module openframe_project_wrapper (por_l,
    porb_h,
    porb_l,
    resetb_h,
    resetb_l,
    analog_io,
    analog_noesd_io,
    gpio_analog_en,
    gpio_analog_pol,
    gpio_analog_sel,
    gpio_dm0,
    gpio_dm1,
    gpio_dm2,
    gpio_holdover,
    gpio_ib_mode_sel,
    gpio_in,
    gpio_in_h,
    gpio_inp_dis,
    gpio_loopback_one,
    gpio_loopback_zero,
    gpio_oeb,
    gpio_out,
    gpio_slow_sel,
    gpio_vtrip_sel,
    mask_rev);
 input por_l;
 input porb_h;
 input porb_l;
 input resetb_h;
 input resetb_l;
 inout [43:0] analog_io;
 inout [43:0] analog_noesd_io;
 output [43:0] gpio_analog_en;
 output [43:0] gpio_analog_pol;
 output [43:0] gpio_analog_sel;
 output [43:0] gpio_dm0;
 output [43:0] gpio_dm1;
 output [43:0] gpio_dm2;
 output [43:0] gpio_holdover;
 output [43:0] gpio_ib_mode_sel;
 input [43:0] gpio_in;
 input [43:0] gpio_in_h;
 output [43:0] gpio_inp_dis;
 input [43:0] gpio_loopback_one;
 input [43:0] gpio_loopback_zero;
 output [43:0] gpio_oeb;
 output [43:0] gpio_out;
 output [43:0] gpio_slow_sel;
 output [43:0] gpio_vtrip_sel;
 input [31:0] mask_rev;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire net2525;
 wire net2559;
 wire _00165_;
 wire _00166_;
 wire net2558;
 wire net2441;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire net2539;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire net2556;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire net2598;
 wire net2600;
 wire _02918_;
 wire net2443;
 wire net2315;
 wire _02921_;
 wire _02922_;
 wire net2617;
 wire net2625;
 wire _02925_;
 wire net2312;
 wire net2612;
 wire _02928_;
 wire net2609;
 wire _02930_;
 wire net2336;
 wire net2608;
 wire _02933_;
 wire net2606;
 wire _02935_;
 wire net2335;
 wire net2604;
 wire _02938_;
 wire net2602;
 wire _02940_;
 wire net2445;
 wire _02942_;
 wire _02943_;
 wire net2446;
 wire net2307;
 wire _02946_;
 wire _02947_;
 wire net2596;
 wire net2448;
 wire net2314;
 wire _02951_;
 wire _02952_;
 wire net2594;
 wire net2450;
 wire net2343;
 wire _02956_;
 wire _02957_;
 wire net2592;
 wire net2368;
 wire net2350;
 wire _02961_;
 wire net2589;
 wire _02963_;
 wire net2367;
 wire net2358;
 wire _02966_;
 wire net2586;
 wire _02968_;
 wire net2453;
 wire net2364;
 wire _02971_;
 wire _02972_;
 wire net2585;
 wire net2390;
 wire net2371;
 wire _02976_;
 wire net2584;
 wire _02978_;
 wire net2389;
 wire net2379;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire net2582;
 wire net2384;
 wire _02987_;
 wire _02988_;
 wire net2581;
 wire net2459;
 wire net2387;
 wire _02992_;
 wire _02993_;
 wire net2580;
 wire net2462;
 wire net2392;
 wire _02997_;
 wire _02998_;
 wire net2579;
 wire _03000_;
 wire net2467;
 wire net2398;
 wire _03003_;
 wire _03004_;
 wire net2578;
 wire _03006_;
 wire net2414;
 wire net2400;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire net2412;
 wire net2403;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire net2472;
 wire net2385;
 wire _03021_;
 wire _03022_;
 wire net2576;
 wire net2474;
 wire net2388;
 wire _03026_;
 wire _03027_;
 wire net2575;
 wire _03029_;
 wire net2574;
 wire net2404;
 wire _03032_;
 wire _03033_;
 wire net2573;
 wire _03035_;
 wire net2572;
 wire net2410;
 wire _03038_;
 wire _03039_;
 wire net2571;
 wire net2483;
 wire net2396;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire net2491;
 wire net2405;
 wire _03048_;
 wire _03049_;
 wire net2570;
 wire net2494;
 wire net2411;
 wire _03053_;
 wire _03054_;
 wire net2569;
 wire _03056_;
 wire net2496;
 wire net2407;
 wire _03059_;
 wire _03060_;
 wire net2567;
 wire net2499;
 wire net2426;
 wire _03064_;
 wire _03065_;
 wire net2565;
 wire net2505;
 wire net2428;
 wire _03069_;
 wire _03070_;
 wire net2562;
 wire _03072_;
 wire net2517;
 wire net2432;
 wire _03075_;
 wire _03076_;
 wire net2560;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire net1378;
 wire net1377;
 wire net1376;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire net1373;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire net1108;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire net2463;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire net2461;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire net2460;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire net2458;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire net2457;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire net2456;
 wire net2455;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire net2454;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire net2452;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire net2451;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire net2449;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire net2447;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire net2444;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire net2442;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire net2440;
 wire _05896_;
 wire _05897_;
 wire net2439;
 wire net2438;
 wire _05900_;
 wire _05901_;
 wire net2437;
 wire _05903_;
 wire net2436;
 wire net2435;
 wire net2434;
 wire _05907_;
 wire _05908_;
 wire net2433;
 wire _05910_;
 wire net2431;
 wire _05912_;
 wire net2430;
 wire net2429;
 wire net2427;
 wire _05916_;
 wire net2425;
 wire net2424;
 wire net2423;
 wire _05920_;
 wire net2422;
 wire net2421;
 wire net2420;
 wire net2419;
 wire net2418;
 wire net2417;
 wire net2416;
 wire _05928_;
 wire net2415;
 wire net2413;
 wire _05931_;
 wire net2409;
 wire net2408;
 wire net2406;
 wire _05935_;
 wire net2402;
 wire net2401;
 wire _05938_;
 wire net2399;
 wire _05940_;
 wire net2397;
 wire net2395;
 wire net2394;
 wire net2393;
 wire _05945_;
 wire net2391;
 wire _05947_;
 wire _05948_;
 wire net2386;
 wire _05950_;
 wire net2383;
 wire net2382;
 wire net2381;
 wire net2380;
 wire net2378;
 wire net2377;
 wire net2376;
 wire net2375;
 wire net2374;
 wire net2373;
 wire net2372;
 wire _05962_;
 wire net2370;
 wire net2369;
 wire net2366;
 wire net2365;
 wire net2363;
 wire _05968_;
 wire net2362;
 wire net2361;
 wire net2360;
 wire _05972_;
 wire net2359;
 wire net2357;
 wire net2356;
 wire net2355;
 wire net2354;
 wire net2353;
 wire net2352;
 wire net2351;
 wire net2349;
 wire net2348;
 wire net2347;
 wire net2346;
 wire net2345;
 wire net2344;
 wire _05987_;
 wire net2342;
 wire net2341;
 wire net2340;
 wire net2339;
 wire net2338;
 wire net2337;
 wire net2334;
 wire net2333;
 wire net2332;
 wire _05997_;
 wire net2331;
 wire net2330;
 wire net2329;
 wire net2328;
 wire _06002_;
 wire net2327;
 wire net2326;
 wire _06005_;
 wire net2325;
 wire net2324;
 wire net2323;
 wire net2322;
 wire net2321;
 wire _06011_;
 wire net2320;
 wire net2319;
 wire _06014_;
 wire net2318;
 wire net2317;
 wire net2316;
 wire _06018_;
 wire net2313;
 wire net2311;
 wire net2310;
 wire net2309;
 wire _06023_;
 wire net2308;
 wire net2306;
 wire net2305;
 wire net2304;
 wire net2303;
 wire net2302;
 wire net2301;
 wire net2300;
 wire net2299;
 wire _06033_;
 wire net2298;
 wire net2297;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire net2294;
 wire net2293;
 wire _06055_;
 wire net2292;
 wire net2291;
 wire net2290;
 wire net2289;
 wire net2288;
 wire _06061_;
 wire net2287;
 wire net2286;
 wire _06064_;
 wire net2285;
 wire net2284;
 wire net2283;
 wire net2282;
 wire _06069_;
 wire _06070_;
 wire net2281;
 wire net2280;
 wire _06073_;
 wire net2279;
 wire net2278;
 wire net2277;
 wire net2276;
 wire _06078_;
 wire net2275;
 wire net2274;
 wire net2273;
 wire net2272;
 wire net2271;
 wire _06084_;
 wire _06085_;
 wire net2270;
 wire net2269;
 wire _06088_;
 wire net2268;
 wire _06090_;
 wire net2267;
 wire net2266;
 wire _06093_;
 wire net2265;
 wire net2264;
 wire net2263;
 wire net2262;
 wire net2261;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire net2260;
 wire net2259;
 wire _06104_;
 wire net2258;
 wire net2257;
 wire _06107_;
 wire net2256;
 wire net2255;
 wire _06110_;
 wire net2254;
 wire net2253;
 wire _06113_;
 wire _06114_;
 wire net2252;
 wire net2251;
 wire net2250;
 wire _06118_;
 wire net2249;
 wire net2248;
 wire _06121_;
 wire net2247;
 wire net2246;
 wire _06124_;
 wire net2245;
 wire net2244;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire net2243;
 wire net2242;
 wire net2241;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire net2240;
 wire net2239;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire net2238;
 wire _06170_;
 wire net2237;
 wire net2236;
 wire _06173_;
 wire net2235;
 wire net2234;
 wire _06176_;
 wire _06177_;
 wire net2233;
 wire _06179_;
 wire net2232;
 wire net2231;
 wire _06182_;
 wire net2230;
 wire net2229;
 wire _06185_;
 wire _06186_;
 wire net2228;
 wire net2227;
 wire _06189_;
 wire net2226;
 wire _06191_;
 wire net2225;
 wire net2224;
 wire _06194_;
 wire net2223;
 wire net2222;
 wire net2221;
 wire _06198_;
 wire _06199_;
 wire net2220;
 wire _06201_;
 wire net2219;
 wire net2218;
 wire _06204_;
 wire net2217;
 wire net2216;
 wire net2215;
 wire _06208_;
 wire _06209_;
 wire net2214;
 wire _06211_;
 wire _06212_;
 wire net2213;
 wire net2212;
 wire _06215_;
 wire net2211;
 wire net2210;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire net2209;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire net2208;
 wire _06227_;
 wire _06228_;
 wire net2207;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire net2206;
 wire net2205;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire net2204;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire net2203;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire net2202;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire net2201;
 wire net2200;
 wire net2199;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire net2198;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire net2197;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire net2196;
 wire net2195;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire net2194;
 wire net2193;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire net2192;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire net2191;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire net2190;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire net2189;
 wire net2188;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire net2187;
 wire net2186;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire net2185;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire net2184;
 wire net2183;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire net2182;
 wire net2181;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire net2180;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire net2179;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire net2178;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire net2177;
 wire _06521_;
 wire _06522_;
 wire net2176;
 wire _06524_;
 wire net2175;
 wire _06526_;
 wire net2174;
 wire net2173;
 wire _06529_;
 wire net2172;
 wire net2171;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire net2170;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire net2169;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire net2168;
 wire net2167;
 wire _06586_;
 wire net2166;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire net2165;
 wire _06593_;
 wire _06594_;
 wire net2164;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire net2163;
 wire net2162;
 wire _06609_;
 wire net2161;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire net2160;
 wire net2159;
 wire _06640_;
 wire net2158;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire net2157;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire net2156;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire net2155;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire net2154;
 wire _06672_;
 wire _06673_;
 wire net2153;
 wire net2152;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire net2151;
 wire net2150;
 wire _06681_;
 wire net2149;
 wire net2148;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire net2147;
 wire _06697_;
 wire _06698_;
 wire net2146;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire net2145;
 wire net2144;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire net2143;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire net2142;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire net2141;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire net2140;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire net2139;
 wire net2138;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire net2137;
 wire net2136;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire net2135;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire net2134;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire net2133;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire net2132;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire net2131;
 wire net2130;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire net2129;
 wire net2128;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire net2127;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire net2126;
 wire net2125;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire net2124;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire net2123;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire net2122;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire net2121;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire net2120;
 wire net2119;
 wire _07043_;
 wire net2118;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire net2117;
 wire _07050_;
 wire _07051_;
 wire net2116;
 wire _07053_;
 wire _07054_;
 wire net2115;
 wire net2114;
 wire _07057_;
 wire net2113;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire net2112;
 wire _07430_;
 wire net2111;
 wire _07432_;
 wire net2110;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire net2109;
 wire _07485_;
 wire net2108;
 wire net2107;
 wire net2106;
 wire _07489_;
 wire net2105;
 wire net2104;
 wire net2103;
 wire net2102;
 wire _07494_;
 wire net2101;
 wire net2100;
 wire net2099;
 wire _07498_;
 wire net2098;
 wire net2097;
 wire net2096;
 wire net2095;
 wire _07503_;
 wire net2094;
 wire net2093;
 wire _07506_;
 wire net2092;
 wire net2091;
 wire _07509_;
 wire net2090;
 wire net2089;
 wire net2088;
 wire _07513_;
 wire net2087;
 wire _07515_;
 wire net2086;
 wire net2085;
 wire _07518_;
 wire net2084;
 wire net2083;
 wire _07521_;
 wire net2082;
 wire _07523_;
 wire net2081;
 wire _07525_;
 wire net2080;
 wire net2079;
 wire net2078;
 wire _07529_;
 wire net2077;
 wire net2076;
 wire _07532_;
 wire net2075;
 wire net2074;
 wire net2073;
 wire _07536_;
 wire net2072;
 wire _07538_;
 wire net2071;
 wire _07540_;
 wire net2070;
 wire net2069;
 wire net2068;
 wire _07544_;
 wire net2067;
 wire _07546_;
 wire net2066;
 wire net2065;
 wire net2064;
 wire _07550_;
 wire net2063;
 wire _07552_;
 wire net2062;
 wire _07554_;
 wire net2061;
 wire net2060;
 wire _07557_;
 wire net2059;
 wire net2058;
 wire _07560_;
 wire net2057;
 wire net2056;
 wire _07563_;
 wire net2055;
 wire net2054;
 wire _07566_;
 wire net2053;
 wire _07568_;
 wire net2052;
 wire _07570_;
 wire net2051;
 wire net2050;
 wire _07573_;
 wire net2049;
 wire net2048;
 wire _07576_;
 wire net2047;
 wire net2046;
 wire _07579_;
 wire net2045;
 wire _07581_;
 wire net2044;
 wire net2043;
 wire _07584_;
 wire net2042;
 wire net2041;
 wire _07587_;
 wire net2040;
 wire net2039;
 wire _07590_;
 wire net2038;
 wire net2037;
 wire _07593_;
 wire net2036;
 wire net2035;
 wire net2034;
 wire net2033;
 wire _07598_;
 wire net2032;
 wire _07600_;
 wire net2031;
 wire _07602_;
 wire net2030;
 wire net2029;
 wire net2028;
 wire _07606_;
 wire net2027;
 wire net2026;
 wire _07609_;
 wire net2025;
 wire net2024;
 wire _07612_;
 wire net2023;
 wire _07614_;
 wire net2022;
 wire _07616_;
 wire net2021;
 wire net2020;
 wire _07619_;
 wire net2019;
 wire _07621_;
 wire _07622_;
 wire net2018;
 wire net2017;
 wire _07625_;
 wire net2016;
 wire _07627_;
 wire _07628_;
 wire net2015;
 wire _07630_;
 wire net2014;
 wire _07632_;
 wire net2013;
 wire net2012;
 wire _07635_;
 wire net2011;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire net2010;
 wire net2009;
 wire _07642_;
 wire _07643_;
 wire net2008;
 wire _07645_;
 wire net2007;
 wire _07647_;
 wire _07648_;
 wire net2006;
 wire _07650_;
 wire net2005;
 wire _07652_;
 wire net2004;
 wire net2003;
 wire _07655_;
 wire _07656_;
 wire net2002;
 wire _07658_;
 wire net2001;
 wire _07660_;
 wire net2000;
 wire net1999;
 wire _07663_;
 wire _07664_;
 wire net1998;
 wire net1997;
 wire _07667_;
 wire net1996;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire net1995;
 wire net1994;
 wire _07675_;
 wire net1993;
 wire _07677_;
 wire net1992;
 wire net1991;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire net1990;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire net1989;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire net1988;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire net1987;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire net1986;
 wire _07718_;
 wire _07719_;
 wire net1985;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire net1984;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire net1983;
 wire _07734_;
 wire net1982;
 wire net1981;
 wire _07737_;
 wire _07738_;
 wire net1980;
 wire net1979;
 wire _07741_;
 wire _07742_;
 wire net1978;
 wire net1977;
 wire _07745_;
 wire net1976;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire net1975;
 wire net1974;
 wire _07756_;
 wire net1973;
 wire net1972;
 wire _07759_;
 wire _07760_;
 wire net1971;
 wire net1970;
 wire _07763_;
 wire _07764_;
 wire net1969;
 wire net1968;
 wire net1967;
 wire _07768_;
 wire net1966;
 wire _07770_;
 wire net1965;
 wire _07772_;
 wire net1964;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire net1963;
 wire net1962;
 wire _07782_;
 wire net1961;
 wire _07784_;
 wire net1960;
 wire net1959;
 wire _07787_;
 wire net1958;
 wire _07789_;
 wire _07790_;
 wire net1957;
 wire net1956;
 wire _07793_;
 wire net1955;
 wire _07795_;
 wire net1954;
 wire net1953;
 wire _07798_;
 wire _07799_;
 wire net1952;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire net1951;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire net1950;
 wire net1949;
 wire _07851_;
 wire net1948;
 wire _07853_;
 wire _07854_;
 wire net1947;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire net1946;
 wire _07860_;
 wire net1945;
 wire _07862_;
 wire net1944;
 wire _07864_;
 wire net1943;
 wire _07866_;
 wire _07867_;
 wire net1942;
 wire _07869_;
 wire _07870_;
 wire net1941;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire net1940;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire net1939;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire net1938;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire net1937;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire net1936;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire net1935;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire net1934;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire net1933;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire net1932;
 wire _07965_;
 wire net1931;
 wire _07967_;
 wire net1930;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire net1929;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire net1928;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire net1927;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire net1926;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire net1925;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire net1924;
 wire _08057_;
 wire net1923;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire net1922;
 wire _08073_;
 wire net1921;
 wire _08075_;
 wire net1920;
 wire _08077_;
 wire _08078_;
 wire net1919;
 wire _08080_;
 wire _08081_;
 wire net1918;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire net1917;
 wire _08089_;
 wire _08090_;
 wire net1916;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire net1915;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire net1914;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire net1913;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire net1912;
 wire _08124_;
 wire net1911;
 wire _08126_;
 wire _08127_;
 wire net1910;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire net1909;
 wire _08142_;
 wire _08143_;
 wire net1908;
 wire net1907;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire net1906;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire net1905;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire net1904;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire net1903;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire net1902;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire net1901;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire net1900;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire net1899;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire net1898;
 wire _08553_;
 wire net1897;
 wire _08555_;
 wire net1896;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire net1895;
 wire _08568_;
 wire net1894;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire net1893;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire net1892;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire net1891;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire net1890;
 wire _09190_;
 wire net1889;
 wire _09192_;
 wire net1888;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire net1887;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire net1886;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire net1884;
 wire _09369_;
 wire _09370_;
 wire net1883;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire net1882;
 wire net1881;
 wire net1880;
 wire net1879;
 wire _09394_;
 wire net1878;
 wire net1877;
 wire net1876;
 wire net1875;
 wire net1874;
 wire net1873;
 wire _09401_;
 wire net1872;
 wire net1871;
 wire _09404_;
 wire _09405_;
 wire net1870;
 wire net1869;
 wire _09408_;
 wire net1868;
 wire net1867;
 wire _09411_;
 wire net1866;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire net1865;
 wire net1864;
 wire _09418_;
 wire net1863;
 wire net1862;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire net1861;
 wire net1860;
 wire net1859;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire net1858;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire net1857;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire net1856;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire net1855;
 wire net1854;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire net1853;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire net1852;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire net1851;
 wire _09843_;
 wire _09844_;
 wire net1850;
 wire net1849;
 wire net1848;
 wire _09848_;
 wire net1847;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire net1846;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire net1845;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire net1844;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire net1843;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire net1842;
 wire net1841;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire net1840;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire net1839;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire net1838;
 wire _09909_;
 wire net1837;
 wire net1836;
 wire _09912_;
 wire net1835;
 wire net1834;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire net1833;
 wire _09922_;
 wire _09923_;
 wire net1832;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire net1831;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire net1830;
 wire net1829;
 wire _10000_;
 wire _10001_;
 wire net1828;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire net1827;
 wire net1826;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire net1825;
 wire net1824;
 wire net1823;
 wire net1822;
 wire _10029_;
 wire _10030_;
 wire net1821;
 wire net1820;
 wire net1819;
 wire net1818;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire net1817;
 wire _10079_;
 wire _10080_;
 wire net1816;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire net1815;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire net1814;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire net1813;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire net1812;
 wire net1811;
 wire _10125_;
 wire _10126_;
 wire net1810;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire net1809;
 wire _10141_;
 wire _10142_;
 wire net1808;
 wire net1807;
 wire _10145_;
 wire _10146_;
 wire net1806;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire net1805;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire net1804;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire net1803;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire net1802;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire net1801;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire net1800;
 wire net1799;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire net1798;
 wire net1797;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire net1796;
 wire _10336_;
 wire _10337_;
 wire net1795;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire net1794;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire net1793;
 wire _10382_;
 wire _10383_;
 wire net1792;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire net1791;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire net1790;
 wire _10503_;
 wire net1789;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire net1788;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire net1787;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire net1786;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire net1785;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire net1784;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire net1783;
 wire net1782;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire net1781;
 wire _10917_;
 wire _10918_;
 wire net1780;
 wire _10920_;
 wire _10921_;
 wire net1779;
 wire net1778;
 wire _10924_;
 wire net1777;
 wire net1776;
 wire _10927_;
 wire net1775;
 wire _10929_;
 wire net1774;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire net1773;
 wire _10953_;
 wire net1772;
 wire _10955_;
 wire net1771;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire net1770;
 wire net1769;
 wire _10980_;
 wire _10981_;
 wire net1768;
 wire net1767;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire net1766;
 wire net1765;
 wire _11005_;
 wire net1764;
 wire net1763;
 wire _11008_;
 wire _11009_;
 wire net1762;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire net1761;
 wire net1760;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire net1759;
 wire _11032_;
 wire _11033_;
 wire net1758;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire net1757;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire net1756;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire net1755;
 wire _11067_;
 wire net1754;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire net1753;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire net1752;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire net1751;
 wire _11101_;
 wire net1750;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire net1749;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire net1748;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire net1747;
 wire _11135_;
 wire net1746;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire net1745;
 wire _11147_;
 wire net1744;
 wire net1743;
 wire _11150_;
 wire _11151_;
 wire net1742;
 wire _11153_;
 wire net1741;
 wire _11155_;
 wire net1740;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire net1739;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire net1738;
 wire net1737;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire net1736;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire net1735;
 wire _11190_;
 wire net1734;
 wire net1733;
 wire _11193_;
 wire _11194_;
 wire net1732;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire net1731;
 wire net1730;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire net1729;
 wire _11242_;
 wire _11243_;
 wire net1728;
 wire net1727;
 wire _11246_;
 wire _11247_;
 wire net1726;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire net1725;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire net1724;
 wire _11263_;
 wire net1723;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire net1722;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire net1721;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire net1720;
 wire net1719;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire net1718;
 wire _11297_;
 wire _11298_;
 wire net1717;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire net1716;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire net1715;
 wire _11317_;
 wire _11318_;
 wire net1714;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire net1713;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire net1712;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire net1711;
 wire _11342_;
 wire _11343_;
 wire net1710;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire net1709;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire net1708;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire net1707;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire net1706;
 wire _11401_;
 wire _11402_;
 wire net1705;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire net1704;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire net1703;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire net1702;
 wire _11436_;
 wire net1701;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire net1700;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire net1699;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire net1698;
 wire _11470_;
 wire net1697;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire net1696;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire net1695;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire net1694;
 wire net1693;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire net1692;
 wire net1691;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire net1690;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire net1689;
 wire net1688;
 wire _11549_;
 wire _11550_;
 wire net1687;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire net1686;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire net1685;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire net1684;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire net1683;
 wire net1682;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire net1681;
 wire _11592_;
 wire net1680;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire net1679;
 wire _11601_;
 wire _11602_;
 wire net1678;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire net1677;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire net1676;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire net1675;
 wire _11629_;
 wire net1674;
 wire _11631_;
 wire net1673;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire net1672;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire net1671;
 wire net1670;
 wire net1669;
 wire net1668;
 wire _11647_;
 wire net1667;
 wire _11649_;
 wire net1666;
 wire net1665;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire net1664;
 wire _11681_;
 wire _11682_;
 wire net1663;
 wire _11684_;
 wire net1662;
 wire net1661;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire net1660;
 wire _11713_;
 wire _11714_;
 wire net1659;
 wire _11716_;
 wire _11717_;
 wire net1658;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire net1657;
 wire _11724_;
 wire net1656;
 wire net1655;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire net1654;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire net1653;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire net1652;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire net1651;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire net1650;
 wire _11779_;
 wire _11780_;
 wire net1649;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire net1648;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire net1647;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire net1646;
 wire net1645;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire net1644;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire net1643;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire net1642;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire net1641;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire net1640;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire net1639;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire net1638;
 wire net1637;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire net1636;
 wire net1635;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire net1634;
 wire net1633;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire net1632;
 wire net1631;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire net1630;
 wire net1629;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire net1628;
 wire net1627;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire net1626;
 wire net1625;
 wire net1624;
 wire net1623;
 wire net1622;
 wire net1621;
 wire _11942_;
 wire _11943_;
 wire net1620;
 wire _11945_;
 wire _11946_;
 wire net1619;
 wire _11948_;
 wire _11949_;
 wire net1618;
 wire net1617;
 wire _11952_;
 wire _11953_;
 wire net1616;
 wire net1615;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire net1614;
 wire _11966_;
 wire net1613;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire net1612;
 wire net1611;
 wire net1610;
 wire _11993_;
 wire _11994_;
 wire net1609;
 wire _11996_;
 wire net1608;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire net1607;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire net1606;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire net1605;
 wire _12117_;
 wire net1604;
 wire net1603;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire net1602;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire net1601;
 wire _12158_;
 wire net1600;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire net1599;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire net1598;
 wire net1597;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire net1596;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire net1595;
 wire _12201_;
 wire net1594;
 wire net1593;
 wire net1592;
 wire _12205_;
 wire _12206_;
 wire net1591;
 wire _12208_;
 wire _12209_;
 wire net1590;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire net1589;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire net1588;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire net1587;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire net1586;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire net1585;
 wire _12698_;
 wire net1584;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire net1583;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire net1582;
 wire net1581;
 wire _12710_;
 wire net1580;
 wire _12712_;
 wire _12713_;
 wire net1579;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire net1578;
 wire _12720_;
 wire _12721_;
 wire net1577;
 wire net1576;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire net1575;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire net1574;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire net1573;
 wire _12788_;
 wire net1572;
 wire _12790_;
 wire net1571;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire net1570;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire net1569;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire net1568;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire net1567;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire net1566;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire net1565;
 wire _12963_;
 wire net1564;
 wire net1563;
 wire _12966_;
 wire _12967_;
 wire net1562;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire net1561;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire net1560;
 wire net1559;
 wire _12987_;
 wire net1558;
 wire net1557;
 wire _12990_;
 wire net1556;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire net1555;
 wire _12996_;
 wire _12997_;
 wire net1554;
 wire net1553;
 wire net1552;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire net1551;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire net1550;
 wire _13013_;
 wire net1549;
 wire _13015_;
 wire _13016_;
 wire net1548;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire net1547;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire net1546;
 wire _13026_;
 wire _13027_;
 wire net1545;
 wire net1544;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire net1543;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire net1542;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire net1541;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire net1540;
 wire net1539;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire net1538;
 wire _13122_;
 wire net1537;
 wire net1536;
 wire _13125_;
 wire net1535;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire net1534;
 wire _13131_;
 wire net1533;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire net1532;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire net1531;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire net1530;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire net1529;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire net1528;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire net1527;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire net1526;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire net1525;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire net1524;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire net1523;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire net1522;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire net1521;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire net1520;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire net1519;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire net1518;
 wire _13373_;
 wire net1517;
 wire net1516;
 wire _13376_;
 wire net1515;
 wire _13378_;
 wire _13379_;
 wire net1514;
 wire net1513;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire net1512;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire net1511;
 wire net1510;
 wire _13593_;
 wire _13594_;
 wire net1509;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire net1508;
 wire _13600_;
 wire net1507;
 wire _13602_;
 wire _13603_;
 wire net1506;
 wire _13605_;
 wire _13606_;
 wire net1505;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire net1504;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire net1503;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire net1502;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire net1501;
 wire _13799_;
 wire net1500;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire net1499;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire net1498;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire net1497;
 wire net1496;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire net1495;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire net1494;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire net1493;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire net1492;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire net1491;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire net1490;
 wire net1489;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire net1488;
 wire _14604_;
 wire net1487;
 wire net1486;
 wire _14607_;
 wire net1485;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire net1484;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire net1483;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire net1482;
 wire _14665_;
 wire net1481;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire net1480;
 wire net1479;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire net1478;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire net1477;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire net1476;
 wire _14816_;
 wire net1475;
 wire net1474;
 wire _14819_;
 wire net1473;
 wire net1472;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire net1471;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire net1470;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire net1469;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire net1468;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire net1467;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire net1466;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire net1465;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire net1464;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire net1463;
 wire net1462;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire net1461;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire net1460;
 wire net1459;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire net1458;
 wire net1457;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire net1456;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire net1455;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire net1454;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire net1453;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire net1452;
 wire net1451;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire net1450;
 wire _15008_;
 wire _15009_;
 wire net1449;
 wire net1448;
 wire net1447;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire net1446;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire net1445;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire net1444;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire net1443;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire net1442;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire net1441;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire net1440;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire net1439;
 wire net1438;
 wire _15120_;
 wire _15121_;
 wire net1437;
 wire net1436;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire net1435;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire net1434;
 wire _15207_;
 wire net1433;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire net1432;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire net1431;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire net1430;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire net1429;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire net1428;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire net1427;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire net1426;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire net1425;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire net1424;
 wire net1423;
 wire _15633_;
 wire net1422;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire net1421;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire net1420;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire net1419;
 wire _15905_;
 wire net1418;
 wire _15907_;
 wire net1417;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire net1416;
 wire net1415;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire net1414;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire net1413;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire net1412;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire net1411;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire net1410;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire net1409;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire net1408;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire net1407;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire net1406;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire net1405;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire net1404;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire net1403;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire net1402;
 wire net1401;
 wire net1400;
 wire _16059_;
 wire net1399;
 wire net1398;
 wire net1397;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire net1396;
 wire net1395;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire net1394;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire net1393;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire net1392;
 wire _16129_;
 wire _16130_;
 wire net1391;
 wire _16132_;
 wire _16133_;
 wire net1390;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire net1389;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire net1388;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire net1387;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire net1386;
 wire net1385;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire net1384;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire net1383;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire net1382;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire net1381;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire net1380;
 wire net1379;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire net1375;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire net1374;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire net1372;
 wire _16433_;
 wire _16434_;
 wire net1371;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire net1370;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire net1369;
 wire _16469_;
 wire _16470_;
 wire net1368;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire net1367;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire net1366;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire net1365;
 wire _16503_;
 wire _16504_;
 wire net1364;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire net1363;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire net1362;
 wire _16526_;
 wire _16527_;
 wire net1361;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire net1360;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire net1359;
 wire net1358;
 wire _16550_;
 wire _16551_;
 wire net1357;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire net1356;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire net1355;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire net1354;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire net1353;
 wire _16624_;
 wire net1352;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire net1351;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire net1350;
 wire _16663_;
 wire net1349;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire net1348;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire net1347;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire net1346;
 wire _16699_;
 wire _16700_;
 wire net1345;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire net1344;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire net1343;
 wire net1342;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire net1341;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire net1340;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire net1339;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire net1338;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire net1337;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire net1336;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire net1335;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire net1334;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire net1333;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire net1332;
 wire net1331;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire net1330;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire net1329;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire net1328;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire net1327;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire net1326;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire net1325;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire net1324;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire net1323;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire net1322;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire net1321;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire net1320;
 wire _16923_;
 wire net1319;
 wire _16925_;
 wire _16926_;
 wire net1318;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire net1317;
 wire _16937_;
 wire net1316;
 wire _16939_;
 wire _16940_;
 wire net1315;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire net1314;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire net1313;
 wire _16954_;
 wire _16955_;
 wire net1312;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire net1311;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire net1310;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire net1309;
 wire _17033_;
 wire _17034_;
 wire net1308;
 wire _17036_;
 wire _17037_;
 wire net1307;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire net1306;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire net1305;
 wire _17062_;
 wire net1304;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire net1303;
 wire net1302;
 wire _17069_;
 wire _17070_;
 wire net1301;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire net1300;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire net1299;
 wire net1298;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire net1297;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire net1296;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire net1295;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire net1294;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire net1293;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire net1292;
 wire _17170_;
 wire net1291;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire net1290;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire net1289;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire net1288;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire net1287;
 wire _17207_;
 wire _17208_;
 wire net1286;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire net1285;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire net1284;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire net1283;
 wire net1282;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire net1281;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire net1280;
 wire _17268_;
 wire net1279;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire net1278;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire net1277;
 wire _17281_;
 wire net1276;
 wire net1275;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire net1274;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire net1273;
 wire net1272;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire net1271;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire net1270;
 wire _17318_;
 wire net1269;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire net1268;
 wire _17326_;
 wire net1267;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire net1266;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire net1265;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire net1264;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire net1263;
 wire _17363_;
 wire net1262;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire net1261;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire net1260;
 wire _17386_;
 wire net1259;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire net1258;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire net1257;
 wire _17409_;
 wire net1256;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire net1255;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire net1254;
 wire _17433_;
 wire net1253;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire net1252;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire net1251;
 wire _17456_;
 wire net1250;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire net1249;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire net1248;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire net1247;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire net1246;
 wire _17491_;
 wire _17492_;
 wire net1245;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire net1244;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire net1243;
 wire _17506_;
 wire _17507_;
 wire net1242;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire net1241;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire net1240;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire net1239;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire net1238;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire net1237;
 wire _17554_;
 wire _17555_;
 wire net1236;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire net1235;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire net1234;
 wire net1233;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire net1232;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire net1231;
 wire _17589_;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire net1230;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire net1229;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire net1228;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire net1227;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire net1226;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire net1225;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire net1224;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire net1223;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire net1222;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire net1221;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire net1220;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire net1219;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire net1218;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire net1217;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire net1216;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire net1215;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire net1214;
 wire _17725_;
 wire net1213;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire net1212;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire net1211;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire net1210;
 wire net1209;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire net1208;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire net1207;
 wire net1206;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire net1205;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire net1204;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire net1203;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire net1202;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire net1201;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire net1200;
 wire net1199;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire net1198;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire net1197;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire net1196;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire net1195;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire net1194;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire net1193;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire net1192;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire net1191;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire net1190;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire _18109_;
 wire net1189;
 wire _18111_;
 wire _18112_;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire _18117_;
 wire net1188;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire _18124_;
 wire _18125_;
 wire _18126_;
 wire net1187;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire net1186;
 wire _18132_;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire _18145_;
 wire _18146_;
 wire _18147_;
 wire net1185;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire _18176_;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire net1184;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire net1183;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire _18244_;
 wire _18245_;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire _18322_;
 wire _18323_;
 wire _18324_;
 wire _18325_;
 wire _18326_;
 wire _18327_;
 wire net1182;
 wire _18329_;
 wire _18330_;
 wire _18331_;
 wire _18332_;
 wire _18333_;
 wire _18334_;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire _18338_;
 wire _18339_;
 wire _18340_;
 wire _18341_;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire _18354_;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire _18358_;
 wire _18359_;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire _18364_;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire _18368_;
 wire _18369_;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire _18378_;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire _18389_;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire _18396_;
 wire _18397_;
 wire _18398_;
 wire _18399_;
 wire _18400_;
 wire _18401_;
 wire _18402_;
 wire _18403_;
 wire net1181;
 wire _18405_;
 wire _18406_;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire _18411_;
 wire _18412_;
 wire net1180;
 wire net1179;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire _18420_;
 wire _18421_;
 wire _18422_;
 wire _18423_;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire _18428_;
 wire _18429_;
 wire _18430_;
 wire _18431_;
 wire _18432_;
 wire _18433_;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire _18438_;
 wire _18439_;
 wire _18440_;
 wire _18441_;
 wire _18442_;
 wire _18443_;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire _18448_;
 wire _18449_;
 wire _18450_;
 wire _18451_;
 wire _18452_;
 wire _18453_;
 wire _18454_;
 wire _18455_;
 wire _18456_;
 wire _18457_;
 wire _18458_;
 wire _18459_;
 wire _18460_;
 wire net1178;
 wire _18462_;
 wire _18463_;
 wire _18464_;
 wire _18465_;
 wire _18466_;
 wire _18467_;
 wire _18468_;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire _18472_;
 wire _18473_;
 wire _18474_;
 wire _18475_;
 wire net1177;
 wire net1176;
 wire _18478_;
 wire _18479_;
 wire _18480_;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire net1175;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire _18491_;
 wire _18492_;
 wire _18493_;
 wire _18494_;
 wire _18495_;
 wire net1174;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire net1173;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire _18508_;
 wire _18509_;
 wire _18510_;
 wire _18511_;
 wire _18512_;
 wire _18513_;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire _18519_;
 wire _18520_;
 wire net1172;
 wire _18522_;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire net1171;
 wire _18528_;
 wire _18529_;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire _18534_;
 wire _18535_;
 wire net1170;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire _18541_;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire _18546_;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire net1169;
 wire _18557_;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire _18566_;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire _18580_;
 wire _18581_;
 wire _18582_;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire _18606_;
 wire _18607_;
 wire _18608_;
 wire _18609_;
 wire _18610_;
 wire _18611_;
 wire _18612_;
 wire _18613_;
 wire _18614_;
 wire _18615_;
 wire _18616_;
 wire _18617_;
 wire _18618_;
 wire _18619_;
 wire _18620_;
 wire _18621_;
 wire _18622_;
 wire _18623_;
 wire _18624_;
 wire _18625_;
 wire _18626_;
 wire _18627_;
 wire _18628_;
 wire net1168;
 wire _18630_;
 wire _18631_;
 wire _18632_;
 wire _18633_;
 wire _18634_;
 wire _18635_;
 wire _18636_;
 wire _18637_;
 wire _18638_;
 wire _18639_;
 wire _18640_;
 wire _18641_;
 wire _18642_;
 wire _18643_;
 wire _18644_;
 wire _18645_;
 wire _18646_;
 wire _18647_;
 wire _18648_;
 wire _18649_;
 wire _18650_;
 wire _18651_;
 wire _18652_;
 wire _18653_;
 wire _18654_;
 wire _18655_;
 wire _18656_;
 wire _18657_;
 wire _18658_;
 wire _18659_;
 wire _18660_;
 wire _18661_;
 wire _18662_;
 wire _18663_;
 wire _18664_;
 wire _18665_;
 wire _18666_;
 wire _18667_;
 wire _18668_;
 wire _18669_;
 wire _18670_;
 wire _18671_;
 wire _18672_;
 wire _18673_;
 wire _18674_;
 wire _18675_;
 wire _18676_;
 wire _18677_;
 wire _18678_;
 wire _18679_;
 wire _18680_;
 wire _18681_;
 wire _18682_;
 wire _18683_;
 wire _18684_;
 wire _18685_;
 wire _18686_;
 wire _18687_;
 wire _18688_;
 wire _18689_;
 wire _18690_;
 wire _18691_;
 wire _18692_;
 wire _18693_;
 wire _18694_;
 wire _18695_;
 wire _18696_;
 wire _18697_;
 wire _18698_;
 wire _18699_;
 wire _18700_;
 wire _18701_;
 wire _18702_;
 wire _18703_;
 wire _18704_;
 wire _18705_;
 wire _18706_;
 wire _18707_;
 wire _18708_;
 wire _18709_;
 wire _18710_;
 wire _18711_;
 wire _18712_;
 wire _18713_;
 wire _18714_;
 wire _18715_;
 wire _18716_;
 wire _18717_;
 wire _18718_;
 wire _18719_;
 wire _18720_;
 wire _18721_;
 wire _18722_;
 wire _18723_;
 wire _18724_;
 wire _18725_;
 wire _18726_;
 wire _18727_;
 wire _18728_;
 wire _18729_;
 wire _18730_;
 wire _18731_;
 wire _18732_;
 wire _18733_;
 wire net1167;
 wire _18735_;
 wire _18736_;
 wire _18737_;
 wire _18738_;
 wire _18739_;
 wire _18740_;
 wire _18741_;
 wire net1166;
 wire net1165;
 wire _18744_;
 wire _18745_;
 wire _18746_;
 wire _18747_;
 wire _18748_;
 wire _18749_;
 wire _18750_;
 wire _18751_;
 wire _18752_;
 wire net1164;
 wire _18754_;
 wire _18755_;
 wire _18756_;
 wire _18757_;
 wire _18758_;
 wire _18759_;
 wire _18760_;
 wire net1163;
 wire _18762_;
 wire _18763_;
 wire _18764_;
 wire net1162;
 wire _18766_;
 wire _18767_;
 wire _18768_;
 wire net1161;
 wire _18770_;
 wire _18771_;
 wire net1160;
 wire _18773_;
 wire _18774_;
 wire _18775_;
 wire _18776_;
 wire _18777_;
 wire _18778_;
 wire _18779_;
 wire net1159;
 wire _18781_;
 wire net1158;
 wire net1157;
 wire _18784_;
 wire _18785_;
 wire _18786_;
 wire _18787_;
 wire _18788_;
 wire _18789_;
 wire _18790_;
 wire _18791_;
 wire _18792_;
 wire _18793_;
 wire _18794_;
 wire _18795_;
 wire _18796_;
 wire _18797_;
 wire _18798_;
 wire _18799_;
 wire _18800_;
 wire _18801_;
 wire _18802_;
 wire _18803_;
 wire _18804_;
 wire _18805_;
 wire _18806_;
 wire _18807_;
 wire net1156;
 wire _18809_;
 wire net1155;
 wire _18811_;
 wire _18812_;
 wire _18813_;
 wire _18814_;
 wire _18815_;
 wire _18816_;
 wire _18817_;
 wire _18818_;
 wire _18819_;
 wire _18820_;
 wire _18821_;
 wire _18822_;
 wire _18823_;
 wire _18824_;
 wire _18825_;
 wire net1154;
 wire _18827_;
 wire _18828_;
 wire _18829_;
 wire _18830_;
 wire _18831_;
 wire _18832_;
 wire _18833_;
 wire _18834_;
 wire _18835_;
 wire _18836_;
 wire _18837_;
 wire _18838_;
 wire _18839_;
 wire _18840_;
 wire _18841_;
 wire _18842_;
 wire _18843_;
 wire _18844_;
 wire _18845_;
 wire _18846_;
 wire _18847_;
 wire _18848_;
 wire _18849_;
 wire _18850_;
 wire _18851_;
 wire _18852_;
 wire _18853_;
 wire _18854_;
 wire _18855_;
 wire _18856_;
 wire _18857_;
 wire _18858_;
 wire net1153;
 wire _18860_;
 wire _18861_;
 wire _18862_;
 wire _18863_;
 wire _18864_;
 wire _18865_;
 wire _18866_;
 wire _18867_;
 wire _18868_;
 wire _18869_;
 wire _18870_;
 wire _18871_;
 wire _18872_;
 wire _18873_;
 wire _18874_;
 wire net1152;
 wire _18876_;
 wire _18877_;
 wire _18878_;
 wire _18879_;
 wire _18880_;
 wire _18881_;
 wire _18882_;
 wire _18883_;
 wire _18884_;
 wire _18885_;
 wire _18886_;
 wire _18887_;
 wire _18888_;
 wire _18889_;
 wire _18890_;
 wire _18891_;
 wire _18892_;
 wire _18893_;
 wire _18894_;
 wire _18895_;
 wire _18896_;
 wire _18897_;
 wire _18898_;
 wire _18899_;
 wire _18900_;
 wire _18901_;
 wire _18902_;
 wire _18903_;
 wire _18904_;
 wire _18905_;
 wire _18906_;
 wire _18907_;
 wire _18908_;
 wire _18909_;
 wire _18910_;
 wire _18911_;
 wire _18912_;
 wire _18913_;
 wire _18914_;
 wire _18915_;
 wire _18916_;
 wire _18917_;
 wire _18918_;
 wire _18919_;
 wire _18920_;
 wire _18921_;
 wire _18922_;
 wire _18923_;
 wire _18924_;
 wire _18925_;
 wire _18926_;
 wire _18927_;
 wire _18928_;
 wire _18929_;
 wire _18930_;
 wire _18931_;
 wire _18932_;
 wire _18933_;
 wire _18934_;
 wire _18935_;
 wire _18936_;
 wire _18937_;
 wire _18938_;
 wire _18939_;
 wire _18940_;
 wire _18941_;
 wire _18942_;
 wire _18943_;
 wire _18944_;
 wire _18945_;
 wire _18946_;
 wire _18947_;
 wire _18948_;
 wire _18949_;
 wire _18950_;
 wire _18951_;
 wire _18952_;
 wire _18953_;
 wire _18954_;
 wire _18955_;
 wire _18956_;
 wire _18957_;
 wire _18958_;
 wire _18959_;
 wire _18960_;
 wire _18961_;
 wire _18962_;
 wire _18963_;
 wire _18964_;
 wire _18965_;
 wire _18966_;
 wire _18967_;
 wire _18968_;
 wire _18969_;
 wire _18970_;
 wire _18971_;
 wire _18972_;
 wire _18973_;
 wire _18974_;
 wire _18975_;
 wire _18976_;
 wire _18977_;
 wire _18978_;
 wire _18979_;
 wire _18980_;
 wire _18981_;
 wire _18982_;
 wire _18983_;
 wire _18984_;
 wire _18985_;
 wire _18986_;
 wire _18987_;
 wire _18988_;
 wire _18989_;
 wire _18990_;
 wire _18991_;
 wire _18992_;
 wire _18993_;
 wire _18994_;
 wire _18995_;
 wire _18996_;
 wire _18997_;
 wire _18998_;
 wire _18999_;
 wire _19000_;
 wire _19001_;
 wire _19002_;
 wire _19003_;
 wire _19004_;
 wire _19005_;
 wire _19006_;
 wire _19007_;
 wire _19008_;
 wire _19009_;
 wire _19010_;
 wire _19011_;
 wire _19012_;
 wire _19013_;
 wire _19014_;
 wire _19015_;
 wire _19016_;
 wire _19017_;
 wire _19018_;
 wire _19019_;
 wire _19020_;
 wire _19021_;
 wire _19022_;
 wire _19023_;
 wire _19024_;
 wire _19025_;
 wire _19026_;
 wire _19027_;
 wire _19028_;
 wire _19029_;
 wire _19030_;
 wire _19031_;
 wire _19032_;
 wire _19033_;
 wire _19034_;
 wire _19035_;
 wire _19036_;
 wire _19037_;
 wire _19038_;
 wire _19039_;
 wire _19040_;
 wire _19041_;
 wire _19042_;
 wire _19043_;
 wire _19044_;
 wire _19045_;
 wire _19046_;
 wire _19047_;
 wire _19048_;
 wire _19049_;
 wire net1151;
 wire _19051_;
 wire _19052_;
 wire _19053_;
 wire _19054_;
 wire _19055_;
 wire _19056_;
 wire _19057_;
 wire _19058_;
 wire _19059_;
 wire _19060_;
 wire net1150;
 wire _19062_;
 wire _19063_;
 wire _19064_;
 wire _19065_;
 wire _19066_;
 wire _19067_;
 wire _19068_;
 wire _19069_;
 wire _19070_;
 wire _19071_;
 wire _19072_;
 wire _19073_;
 wire _19074_;
 wire _19075_;
 wire _19076_;
 wire _19077_;
 wire _19078_;
 wire _19079_;
 wire _19080_;
 wire _19081_;
 wire _19082_;
 wire _19083_;
 wire _19084_;
 wire _19085_;
 wire _19086_;
 wire _19087_;
 wire _19088_;
 wire _19089_;
 wire _19090_;
 wire _19091_;
 wire _19092_;
 wire _19093_;
 wire _19094_;
 wire _19095_;
 wire _19096_;
 wire _19097_;
 wire _19098_;
 wire net1149;
 wire _19100_;
 wire _19101_;
 wire _19102_;
 wire _19103_;
 wire _19104_;
 wire _19105_;
 wire net1148;
 wire net1147;
 wire _19108_;
 wire _19109_;
 wire _19110_;
 wire _19111_;
 wire net1146;
 wire _19113_;
 wire _19114_;
 wire _19115_;
 wire _19116_;
 wire _19117_;
 wire _19118_;
 wire _19119_;
 wire _19120_;
 wire _19121_;
 wire _19122_;
 wire _19123_;
 wire _19124_;
 wire _19125_;
 wire _19126_;
 wire _19127_;
 wire _19128_;
 wire _19129_;
 wire _19130_;
 wire _19131_;
 wire _19132_;
 wire _19133_;
 wire _19134_;
 wire net1145;
 wire _19136_;
 wire net1144;
 wire _19138_;
 wire _19139_;
 wire _19140_;
 wire net1143;
 wire _19142_;
 wire _19143_;
 wire _19144_;
 wire _19145_;
 wire _19146_;
 wire _19147_;
 wire _19148_;
 wire _19149_;
 wire _19150_;
 wire _19151_;
 wire _19152_;
 wire _19153_;
 wire _19154_;
 wire _19155_;
 wire _19156_;
 wire _19157_;
 wire _19158_;
 wire _19159_;
 wire _19160_;
 wire _19161_;
 wire _19162_;
 wire _19163_;
 wire _19164_;
 wire _19165_;
 wire _19166_;
 wire _19167_;
 wire net1142;
 wire _19169_;
 wire _19170_;
 wire net1141;
 wire _19172_;
 wire _19173_;
 wire _19174_;
 wire _19175_;
 wire _19176_;
 wire _19177_;
 wire _19178_;
 wire net1140;
 wire _19180_;
 wire _19181_;
 wire _19182_;
 wire _19183_;
 wire _19184_;
 wire _19185_;
 wire _19186_;
 wire _19187_;
 wire _19188_;
 wire _19189_;
 wire _19190_;
 wire _19191_;
 wire _19192_;
 wire _19193_;
 wire _19194_;
 wire _19195_;
 wire net1139;
 wire _19197_;
 wire _19198_;
 wire net1138;
 wire _19200_;
 wire _19201_;
 wire _19202_;
 wire _19203_;
 wire _19204_;
 wire _19205_;
 wire _19206_;
 wire _19207_;
 wire _19208_;
 wire _19209_;
 wire _19210_;
 wire _19211_;
 wire _19212_;
 wire _19213_;
 wire _19214_;
 wire _19215_;
 wire _19216_;
 wire _19217_;
 wire _19218_;
 wire _19219_;
 wire _19220_;
 wire _19221_;
 wire _19222_;
 wire _19223_;
 wire _19224_;
 wire _19225_;
 wire _19226_;
 wire _19227_;
 wire _19228_;
 wire _19229_;
 wire _19230_;
 wire _19231_;
 wire _19232_;
 wire _19233_;
 wire _19234_;
 wire _19235_;
 wire _19236_;
 wire _19237_;
 wire _19238_;
 wire _19239_;
 wire _19240_;
 wire _19241_;
 wire _19242_;
 wire _19243_;
 wire _19244_;
 wire _19245_;
 wire _19246_;
 wire _19247_;
 wire _19248_;
 wire _19249_;
 wire _19250_;
 wire _19251_;
 wire _19252_;
 wire _19253_;
 wire _19254_;
 wire _19255_;
 wire _19256_;
 wire _19257_;
 wire _19258_;
 wire _19259_;
 wire _19260_;
 wire _19261_;
 wire _19262_;
 wire _19263_;
 wire _19264_;
 wire _19265_;
 wire _19266_;
 wire _19267_;
 wire _19268_;
 wire _19269_;
 wire _19270_;
 wire _19271_;
 wire _19272_;
 wire _19273_;
 wire _19274_;
 wire _19275_;
 wire _19276_;
 wire _19277_;
 wire _19278_;
 wire _19279_;
 wire _19280_;
 wire _19281_;
 wire _19282_;
 wire _19283_;
 wire _19284_;
 wire _19285_;
 wire _19286_;
 wire _19287_;
 wire _19288_;
 wire _19289_;
 wire _19290_;
 wire _19291_;
 wire _19292_;
 wire _19293_;
 wire _19294_;
 wire _19295_;
 wire _19296_;
 wire _19297_;
 wire _19298_;
 wire _19299_;
 wire _19300_;
 wire _19301_;
 wire _19302_;
 wire _19303_;
 wire _19304_;
 wire _19305_;
 wire _19306_;
 wire _19307_;
 wire _19308_;
 wire _19309_;
 wire _19310_;
 wire _19311_;
 wire _19312_;
 wire _19313_;
 wire _19314_;
 wire _19315_;
 wire _19316_;
 wire _19317_;
 wire _19318_;
 wire _19319_;
 wire _19320_;
 wire _19321_;
 wire _19322_;
 wire _19323_;
 wire _19324_;
 wire _19325_;
 wire _19326_;
 wire _19327_;
 wire _19328_;
 wire _19329_;
 wire _19330_;
 wire _19331_;
 wire _19332_;
 wire _19333_;
 wire _19334_;
 wire _19335_;
 wire _19336_;
 wire _19337_;
 wire _19338_;
 wire _19339_;
 wire _19340_;
 wire _19341_;
 wire _19342_;
 wire _19343_;
 wire _19344_;
 wire _19345_;
 wire _19346_;
 wire _19347_;
 wire _19348_;
 wire _19349_;
 wire _19350_;
 wire _19351_;
 wire _19352_;
 wire _19353_;
 wire _19354_;
 wire _19355_;
 wire _19356_;
 wire _19357_;
 wire _19358_;
 wire _19359_;
 wire _19360_;
 wire _19361_;
 wire _19362_;
 wire _19363_;
 wire _19364_;
 wire _19365_;
 wire _19366_;
 wire _19367_;
 wire _19368_;
 wire _19369_;
 wire _19370_;
 wire _19371_;
 wire _19372_;
 wire _19373_;
 wire _19374_;
 wire _19375_;
 wire _19376_;
 wire _19377_;
 wire _19378_;
 wire _19379_;
 wire _19380_;
 wire _19381_;
 wire _19382_;
 wire _19383_;
 wire _19384_;
 wire _19385_;
 wire _19386_;
 wire _19387_;
 wire _19388_;
 wire _19389_;
 wire _19390_;
 wire _19391_;
 wire _19392_;
 wire _19393_;
 wire _19394_;
 wire net1137;
 wire _19396_;
 wire _19397_;
 wire net1136;
 wire net1135;
 wire _19400_;
 wire _19401_;
 wire _19402_;
 wire _19403_;
 wire _19404_;
 wire _19405_;
 wire _19406_;
 wire net1134;
 wire _19408_;
 wire _19409_;
 wire net1133;
 wire _19411_;
 wire _19412_;
 wire _19413_;
 wire _19414_;
 wire _19415_;
 wire _19416_;
 wire _19417_;
 wire _19418_;
 wire _19419_;
 wire _19420_;
 wire _19421_;
 wire _19422_;
 wire _19423_;
 wire net1132;
 wire _19425_;
 wire _19426_;
 wire _19427_;
 wire _19428_;
 wire _19429_;
 wire _19430_;
 wire _19431_;
 wire _19432_;
 wire _19433_;
 wire _19434_;
 wire _19435_;
 wire _19436_;
 wire _19437_;
 wire _19438_;
 wire _19439_;
 wire _19440_;
 wire _19441_;
 wire _19442_;
 wire _19443_;
 wire _19444_;
 wire _19445_;
 wire _19446_;
 wire _19447_;
 wire _19448_;
 wire _19449_;
 wire _19450_;
 wire _19451_;
 wire _19452_;
 wire _19453_;
 wire _19454_;
 wire _19455_;
 wire _19456_;
 wire _19457_;
 wire _19458_;
 wire _19459_;
 wire _19460_;
 wire net1131;
 wire _19462_;
 wire _19463_;
 wire _19464_;
 wire _19465_;
 wire _19466_;
 wire _19467_;
 wire _19468_;
 wire _19469_;
 wire _19470_;
 wire _19471_;
 wire net1130;
 wire _19473_;
 wire _19474_;
 wire _19475_;
 wire _19476_;
 wire _19477_;
 wire _19478_;
 wire _19479_;
 wire _19480_;
 wire _19481_;
 wire _19482_;
 wire _19483_;
 wire _19484_;
 wire _19485_;
 wire _19486_;
 wire _19487_;
 wire _19488_;
 wire _19489_;
 wire _19490_;
 wire _19491_;
 wire _19492_;
 wire _19493_;
 wire _19494_;
 wire _19495_;
 wire _19496_;
 wire _19497_;
 wire _19498_;
 wire _19499_;
 wire _19500_;
 wire _19501_;
 wire _19502_;
 wire _19503_;
 wire _19504_;
 wire _19505_;
 wire net1129;
 wire net1128;
 wire _19508_;
 wire _19509_;
 wire _19510_;
 wire _19511_;
 wire _19512_;
 wire _19513_;
 wire _19514_;
 wire _19515_;
 wire _19516_;
 wire _19517_;
 wire _19518_;
 wire net1127;
 wire _19520_;
 wire _19521_;
 wire _19522_;
 wire _19523_;
 wire net1126;
 wire _19525_;
 wire _19526_;
 wire _19527_;
 wire _19528_;
 wire _19529_;
 wire net1125;
 wire _19531_;
 wire _19532_;
 wire _19533_;
 wire net1124;
 wire _19535_;
 wire _19536_;
 wire _19537_;
 wire _19538_;
 wire _19539_;
 wire _19540_;
 wire _19541_;
 wire _19542_;
 wire _19543_;
 wire _19544_;
 wire net1123;
 wire net1122;
 wire net1121;
 wire _19548_;
 wire _19549_;
 wire _19550_;
 wire _19551_;
 wire _19552_;
 wire _19553_;
 wire _19554_;
 wire _19555_;
 wire _19556_;
 wire net1120;
 wire net1119;
 wire _19559_;
 wire _19560_;
 wire _19561_;
 wire _19562_;
 wire _19563_;
 wire _19564_;
 wire _19565_;
 wire _19566_;
 wire _19567_;
 wire _19568_;
 wire _19569_;
 wire _19570_;
 wire _19571_;
 wire _19572_;
 wire _19573_;
 wire _19574_;
 wire _19575_;
 wire _19576_;
 wire _19577_;
 wire _19578_;
 wire _19579_;
 wire _19580_;
 wire _19581_;
 wire _19582_;
 wire _19583_;
 wire _19584_;
 wire _19585_;
 wire _19586_;
 wire _19587_;
 wire _19588_;
 wire _19589_;
 wire _19590_;
 wire _19591_;
 wire net1118;
 wire _19593_;
 wire _19594_;
 wire _19595_;
 wire _19596_;
 wire _19597_;
 wire _19598_;
 wire _19599_;
 wire _19600_;
 wire _19601_;
 wire _19602_;
 wire _19603_;
 wire _19604_;
 wire net1117;
 wire _19606_;
 wire net1116;
 wire net1115;
 wire _19609_;
 wire _19610_;
 wire _19611_;
 wire _19612_;
 wire _19613_;
 wire _19614_;
 wire _19615_;
 wire _19616_;
 wire _19617_;
 wire _19618_;
 wire _19619_;
 wire _19620_;
 wire _19621_;
 wire _19622_;
 wire _19623_;
 wire net1114;
 wire _19625_;
 wire _19626_;
 wire _19627_;
 wire _19628_;
 wire _19629_;
 wire _19630_;
 wire net1113;
 wire _19632_;
 wire _19633_;
 wire _19634_;
 wire net1112;
 wire _19636_;
 wire _19637_;
 wire _19638_;
 wire _19639_;
 wire _19640_;
 wire _19641_;
 wire net1111;
 wire _19643_;
 wire _19644_;
 wire _19645_;
 wire _19646_;
 wire _19647_;
 wire net1110;
 wire _19649_;
 wire _19650_;
 wire _19651_;
 wire _19652_;
 wire net1109;
 wire _19654_;
 wire _19655_;
 wire _19656_;
 wire _19657_;
 wire _19658_;
 wire _19659_;
 wire _19660_;
 wire _19661_;
 wire _19662_;
 wire _19663_;
 wire _19664_;
 wire _19665_;
 wire _19666_;
 wire _19667_;
 wire _19668_;
 wire _19669_;
 wire _19670_;
 wire net1107;
 wire _19672_;
 wire net1106;
 wire _19674_;
 wire net1105;
 wire _19676_;
 wire _19677_;
 wire _19678_;
 wire _19679_;
 wire _19680_;
 wire _19681_;
 wire _19682_;
 wire _19683_;
 wire _19684_;
 wire _19685_;
 wire _19686_;
 wire _19687_;
 wire _19688_;
 wire _19689_;
 wire _19690_;
 wire _19691_;
 wire net1104;
 wire _19693_;
 wire _19694_;
 wire net1103;
 wire _19696_;
 wire _19697_;
 wire _19698_;
 wire _19699_;
 wire _19700_;
 wire _19701_;
 wire _19702_;
 wire _19703_;
 wire _19704_;
 wire _19705_;
 wire _19706_;
 wire _19707_;
 wire _19708_;
 wire _19709_;
 wire _19710_;
 wire _19711_;
 wire _19712_;
 wire _19713_;
 wire _19714_;
 wire _19715_;
 wire _19716_;
 wire _19717_;
 wire _19718_;
 wire _19719_;
 wire _19720_;
 wire _19721_;
 wire _19722_;
 wire _19723_;
 wire _19724_;
 wire _19725_;
 wire _19726_;
 wire _19727_;
 wire _19728_;
 wire _19729_;
 wire _19730_;
 wire _19731_;
 wire _19732_;
 wire _19733_;
 wire _19734_;
 wire _19735_;
 wire _19736_;
 wire _19737_;
 wire _19738_;
 wire _19739_;
 wire _19740_;
 wire _19741_;
 wire _19742_;
 wire _19743_;
 wire _19744_;
 wire _19745_;
 wire _19746_;
 wire _19747_;
 wire _19748_;
 wire _19749_;
 wire _19750_;
 wire _19751_;
 wire _19752_;
 wire _19753_;
 wire _19754_;
 wire _19755_;
 wire _19756_;
 wire _19757_;
 wire _19758_;
 wire _19759_;
 wire _19760_;
 wire _19761_;
 wire _19762_;
 wire _19763_;
 wire _19764_;
 wire _19765_;
 wire _19766_;
 wire _19767_;
 wire _19768_;
 wire _19769_;
 wire _19770_;
 wire _19771_;
 wire _19772_;
 wire _19773_;
 wire _19774_;
 wire _19775_;
 wire _19776_;
 wire _19777_;
 wire _19778_;
 wire _19779_;
 wire _19780_;
 wire _19781_;
 wire _19782_;
 wire _19783_;
 wire _19784_;
 wire _19785_;
 wire _19786_;
 wire _19787_;
 wire _19788_;
 wire _19789_;
 wire _19790_;
 wire _19791_;
 wire _19792_;
 wire _19793_;
 wire _19794_;
 wire _19795_;
 wire _19796_;
 wire net1102;
 wire _19798_;
 wire _19799_;
 wire _19800_;
 wire _19801_;
 wire _19802_;
 wire _19803_;
 wire _19804_;
 wire _19805_;
 wire _19806_;
 wire _19807_;
 wire _19808_;
 wire _19809_;
 wire _19810_;
 wire _19811_;
 wire _19812_;
 wire _19813_;
 wire _19814_;
 wire _19815_;
 wire _19816_;
 wire _19817_;
 wire _19818_;
 wire _19819_;
 wire _19820_;
 wire _19821_;
 wire _19822_;
 wire _19823_;
 wire _19824_;
 wire _19825_;
 wire _19826_;
 wire _19827_;
 wire _19828_;
 wire _19829_;
 wire _19830_;
 wire _19831_;
 wire _19832_;
 wire _19833_;
 wire _19834_;
 wire _19835_;
 wire _19836_;
 wire _19837_;
 wire _19838_;
 wire _19839_;
 wire _19840_;
 wire _19841_;
 wire _19842_;
 wire _19843_;
 wire _19844_;
 wire _19845_;
 wire net2635;
 wire _19847_;
 wire net2634;
 wire _19849_;
 wire _19850_;
 wire net2633;
 wire _19852_;
 wire net2632;
 wire _19854_;
 wire _19855_;
 wire _19856_;
 wire _19857_;
 wire _19858_;
 wire _19859_;
 wire _19860_;
 wire _19861_;
 wire net2631;
 wire _19863_;
 wire net2630;
 wire _19865_;
 wire net2629;
 wire _19867_;
 wire _19868_;
 wire _19869_;
 wire _19870_;
 wire _19871_;
 wire _19872_;
 wire net2628;
 wire net2627;
 wire _19875_;
 wire net2626;
 wire _19877_;
 wire _19878_;
 wire _19879_;
 wire _19880_;
 wire _19881_;
 wire _19882_;
 wire _19883_;
 wire _19884_;
 wire _19885_;
 wire _19886_;
 wire net2624;
 wire net2623;
 wire _19889_;
 wire net2622;
 wire net2621;
 wire net2620;
 wire _19893_;
 wire net2619;
 wire net2618;
 wire _19896_;
 wire _19897_;
 wire _19898_;
 wire _19899_;
 wire _19900_;
 wire net2616;
 wire _19902_;
 wire net2615;
 wire net2614;
 wire _19905_;
 wire _19906_;
 wire _19907_;
 wire net2613;
 wire _19909_;
 wire _19910_;
 wire _19911_;
 wire net2611;
 wire net2610;
 wire _19914_;
 wire _19915_;
 wire _19916_;
 wire _19917_;
 wire _19918_;
 wire _19919_;
 wire _19920_;
 wire _19921_;
 wire _19922_;
 wire _19923_;
 wire _19924_;
 wire _19925_;
 wire _19926_;
 wire _19927_;
 wire _19928_;
 wire _19929_;
 wire _19930_;
 wire net2607;
 wire _19932_;
 wire net2605;
 wire _19934_;
 wire _19935_;
 wire _19936_;
 wire _19937_;
 wire _19938_;
 wire _19939_;
 wire _19940_;
 wire _19941_;
 wire _19942_;
 wire _19943_;
 wire _19944_;
 wire net2603;
 wire _19946_;
 wire _19947_;
 wire _19948_;
 wire _19949_;
 wire _19950_;
 wire _19951_;
 wire _19952_;
 wire net2601;
 wire _19954_;
 wire _19955_;
 wire _19956_;
 wire _19957_;
 wire net2599;
 wire _19959_;
 wire _19960_;
 wire _19961_;
 wire _19962_;
 wire net2597;
 wire _19964_;
 wire _19965_;
 wire _19966_;
 wire _19967_;
 wire net2595;
 wire _19969_;
 wire _19970_;
 wire _19971_;
 wire _19972_;
 wire _19973_;
 wire _19974_;
 wire net2593;
 wire _19976_;
 wire net2591;
 wire net2590;
 wire _19979_;
 wire _19980_;
 wire _19981_;
 wire _19982_;
 wire _19983_;
 wire _19984_;
 wire net2588;
 wire _19986_;
 wire _19987_;
 wire _19988_;
 wire _19989_;
 wire _19990_;
 wire net2587;
 wire _19992_;
 wire _19993_;
 wire _19994_;
 wire _19995_;
 wire _19996_;
 wire _19997_;
 wire _19998_;
 wire _19999_;
 wire _20000_;
 wire _20001_;
 wire _20002_;
 wire _20003_;
 wire net2583;
 wire _20005_;
 wire _20006_;
 wire _20007_;
 wire _20008_;
 wire _20009_;
 wire _20010_;
 wire _20011_;
 wire _20012_;
 wire _20013_;
 wire _20014_;
 wire _20015_;
 wire _20016_;
 wire _20017_;
 wire _20018_;
 wire _20019_;
 wire _20020_;
 wire _20021_;
 wire _20022_;
 wire _20023_;
 wire _20024_;
 wire _20025_;
 wire _20026_;
 wire _20027_;
 wire _20028_;
 wire _20029_;
 wire _20030_;
 wire _20031_;
 wire _20032_;
 wire _20033_;
 wire _20034_;
 wire _20035_;
 wire _20036_;
 wire _20037_;
 wire _20038_;
 wire _20039_;
 wire _20040_;
 wire _20041_;
 wire _20042_;
 wire _20043_;
 wire _20044_;
 wire _20045_;
 wire _20046_;
 wire _20047_;
 wire _20048_;
 wire net2577;
 wire _20050_;
 wire _20051_;
 wire _20052_;
 wire _20053_;
 wire _20054_;
 wire _20055_;
 wire _20056_;
 wire _20057_;
 wire _20058_;
 wire _20059_;
 wire _20060_;
 wire _20061_;
 wire _20062_;
 wire _20063_;
 wire _20064_;
 wire _20065_;
 wire _20066_;
 wire _20067_;
 wire _20068_;
 wire _20069_;
 wire _20070_;
 wire _20071_;
 wire _20072_;
 wire _20073_;
 wire _20074_;
 wire _20075_;
 wire _20076_;
 wire _20077_;
 wire _20078_;
 wire _20079_;
 wire _20080_;
 wire _20081_;
 wire _20082_;
 wire _20083_;
 wire _20084_;
 wire _20085_;
 wire _20086_;
 wire _20087_;
 wire _20088_;
 wire _20089_;
 wire _20090_;
 wire _20091_;
 wire _20092_;
 wire net2568;
 wire _20094_;
 wire _20095_;
 wire _20096_;
 wire _20097_;
 wire _20098_;
 wire _20099_;
 wire _20100_;
 wire net2566;
 wire _20102_;
 wire _20103_;
 wire _20104_;
 wire _20105_;
 wire _20106_;
 wire _20107_;
 wire net2564;
 wire net2563;
 wire _20110_;
 wire _20111_;
 wire _20112_;
 wire _20113_;
 wire _20114_;
 wire _20115_;
 wire net2561;
 wire _20117_;
 wire _20118_;
 wire _20119_;
 wire _20120_;
 wire _20121_;
 wire _20122_;
 wire _20123_;
 wire _20124_;
 wire _20125_;
 wire _20126_;
 wire _20127_;
 wire _20128_;
 wire _20129_;
 wire _20130_;
 wire net2557;
 wire _20132_;
 wire _20133_;
 wire _20134_;
 wire _20135_;
 wire _20136_;
 wire _20137_;
 wire _20138_;
 wire net2555;
 wire _20140_;
 wire _20141_;
 wire _20142_;
 wire _20143_;
 wire _20144_;
 wire _20145_;
 wire _20146_;
 wire _20147_;
 wire _20148_;
 wire _20149_;
 wire _20150_;
 wire _20151_;
 wire _20152_;
 wire _20153_;
 wire _20154_;
 wire _20155_;
 wire _20156_;
 wire _20157_;
 wire _20158_;
 wire _20159_;
 wire _20160_;
 wire net2554;
 wire _20162_;
 wire _20163_;
 wire _20164_;
 wire _20165_;
 wire _20166_;
 wire _20167_;
 wire _20168_;
 wire _20169_;
 wire _20170_;
 wire _20171_;
 wire _20172_;
 wire _20173_;
 wire _20174_;
 wire _20175_;
 wire _20176_;
 wire _20177_;
 wire _20178_;
 wire _20179_;
 wire _20180_;
 wire _20181_;
 wire _20182_;
 wire _20183_;
 wire _20184_;
 wire _20185_;
 wire net2553;
 wire _20187_;
 wire _20188_;
 wire _20189_;
 wire _20190_;
 wire _20191_;
 wire _20192_;
 wire _20193_;
 wire _20194_;
 wire _20195_;
 wire _20196_;
 wire _20197_;
 wire _20198_;
 wire _20199_;
 wire _20200_;
 wire _20201_;
 wire _20202_;
 wire _20203_;
 wire _20204_;
 wire _20205_;
 wire _20206_;
 wire _20207_;
 wire _20208_;
 wire _20209_;
 wire _20210_;
 wire _20211_;
 wire _20212_;
 wire _20213_;
 wire _20214_;
 wire _20215_;
 wire _20216_;
 wire _20217_;
 wire _20218_;
 wire _20219_;
 wire _20220_;
 wire _20221_;
 wire _20222_;
 wire _20223_;
 wire _20224_;
 wire _20225_;
 wire _20226_;
 wire _20227_;
 wire _20228_;
 wire net2552;
 wire _20230_;
 wire _20231_;
 wire _20232_;
 wire net2551;
 wire net2550;
 wire _20235_;
 wire _20236_;
 wire _20237_;
 wire _20238_;
 wire _20239_;
 wire _20240_;
 wire _20241_;
 wire _20242_;
 wire _20243_;
 wire _20244_;
 wire _20245_;
 wire _20246_;
 wire _20247_;
 wire _20248_;
 wire _20249_;
 wire _20250_;
 wire _20251_;
 wire _20252_;
 wire _20253_;
 wire _20254_;
 wire _20255_;
 wire net2549;
 wire _20257_;
 wire _20258_;
 wire _20259_;
 wire _20260_;
 wire _20261_;
 wire _20262_;
 wire _20263_;
 wire _20264_;
 wire _20265_;
 wire _20266_;
 wire _20267_;
 wire _20268_;
 wire _20269_;
 wire _20270_;
 wire _20271_;
 wire _20272_;
 wire _20273_;
 wire _20274_;
 wire _20275_;
 wire _20276_;
 wire _20277_;
 wire _20278_;
 wire _20279_;
 wire _20280_;
 wire _20281_;
 wire _20282_;
 wire _20283_;
 wire _20284_;
 wire _20285_;
 wire net2548;
 wire _20287_;
 wire _20288_;
 wire _20289_;
 wire _20290_;
 wire _20291_;
 wire _20292_;
 wire _20293_;
 wire _20294_;
 wire _20295_;
 wire _20296_;
 wire _20297_;
 wire _20298_;
 wire _20299_;
 wire _20300_;
 wire _20301_;
 wire _20302_;
 wire _20303_;
 wire _20304_;
 wire _20305_;
 wire _20306_;
 wire _20307_;
 wire _20308_;
 wire _20309_;
 wire _20310_;
 wire _20311_;
 wire _20312_;
 wire _20313_;
 wire _20314_;
 wire net2547;
 wire _20316_;
 wire _20317_;
 wire _20318_;
 wire _20319_;
 wire _20320_;
 wire _20321_;
 wire _20322_;
 wire _20323_;
 wire _20324_;
 wire _20325_;
 wire _20326_;
 wire _20327_;
 wire _20328_;
 wire _20329_;
 wire _20330_;
 wire _20331_;
 wire _20332_;
 wire _20333_;
 wire _20334_;
 wire _20335_;
 wire _20336_;
 wire _20337_;
 wire _20338_;
 wire net2546;
 wire _20340_;
 wire _20341_;
 wire _20342_;
 wire _20343_;
 wire _20344_;
 wire _20345_;
 wire _20346_;
 wire _20347_;
 wire _20348_;
 wire _20349_;
 wire net2545;
 wire _20351_;
 wire _20352_;
 wire _20353_;
 wire _20354_;
 wire _20355_;
 wire _20356_;
 wire _20357_;
 wire _20358_;
 wire _20359_;
 wire _20360_;
 wire _20361_;
 wire _20362_;
 wire _20363_;
 wire _20364_;
 wire _20365_;
 wire _20366_;
 wire _20367_;
 wire _20368_;
 wire _20369_;
 wire _20370_;
 wire net2544;
 wire net2542;
 wire _20373_;
 wire _20374_;
 wire _20375_;
 wire _20376_;
 wire _20377_;
 wire _20378_;
 wire net2541;
 wire net2540;
 wire _20381_;
 wire net2538;
 wire _20383_;
 wire net2537;
 wire _20385_;
 wire _20386_;
 wire net2536;
 wire _20388_;
 wire net2535;
 wire _20390_;
 wire _20391_;
 wire _20392_;
 wire _20393_;
 wire _20394_;
 wire _20395_;
 wire _20396_;
 wire _20397_;
 wire _20398_;
 wire _20399_;
 wire net2534;
 wire net2533;
 wire _20402_;
 wire _20403_;
 wire net2532;
 wire net2531;
 wire _20406_;
 wire _20407_;
 wire _20408_;
 wire _20409_;
 wire _20410_;
 wire _20411_;
 wire _20412_;
 wire _20413_;
 wire _20414_;
 wire net2530;
 wire _20416_;
 wire _20417_;
 wire _20418_;
 wire _20419_;
 wire _20420_;
 wire _20421_;
 wire _20422_;
 wire net2529;
 wire net2528;
 wire _20425_;
 wire _20426_;
 wire _20427_;
 wire net2527;
 wire net2526;
 wire net2524;
 wire net2523;
 wire _20432_;
 wire _20433_;
 wire _20434_;
 wire _20435_;
 wire _20436_;
 wire net2522;
 wire _20438_;
 wire _20439_;
 wire _20440_;
 wire _20441_;
 wire _20442_;
 wire _20443_;
 wire _20444_;
 wire _20445_;
 wire net2521;
 wire _20447_;
 wire _20448_;
 wire _20449_;
 wire _20450_;
 wire net2520;
 wire _20452_;
 wire _20453_;
 wire _20454_;
 wire _20455_;
 wire _20456_;
 wire _20457_;
 wire _20458_;
 wire _20459_;
 wire _20460_;
 wire _20461_;
 wire _20462_;
 wire _20463_;
 wire _20464_;
 wire _20465_;
 wire net2519;
 wire net2518;
 wire net2516;
 wire net2515;
 wire net2514;
 wire _20471_;
 wire _20472_;
 wire _20473_;
 wire _20474_;
 wire net2513;
 wire _20476_;
 wire net2512;
 wire _20478_;
 wire _20479_;
 wire _20480_;
 wire _20481_;
 wire net2511;
 wire _20483_;
 wire _20484_;
 wire _20485_;
 wire net2510;
 wire _20487_;
 wire _20488_;
 wire _20489_;
 wire _20490_;
 wire _20491_;
 wire _20492_;
 wire net2509;
 wire _20494_;
 wire _20495_;
 wire _20496_;
 wire _20497_;
 wire _20498_;
 wire net2508;
 wire _20500_;
 wire _20501_;
 wire _20502_;
 wire _20503_;
 wire _20504_;
 wire _20505_;
 wire _20506_;
 wire net2507;
 wire net2506;
 wire _20509_;
 wire _20510_;
 wire _20511_;
 wire _20512_;
 wire net2504;
 wire _20514_;
 wire net2503;
 wire _20516_;
 wire _20517_;
 wire _20518_;
 wire _20519_;
 wire _20520_;
 wire _20521_;
 wire _20522_;
 wire _20523_;
 wire _20524_;
 wire _20525_;
 wire _20526_;
 wire _20527_;
 wire _20528_;
 wire _20529_;
 wire _20530_;
 wire _20531_;
 wire _20532_;
 wire _20533_;
 wire _20534_;
 wire _20535_;
 wire net2502;
 wire _20537_;
 wire _20538_;
 wire _20539_;
 wire _20540_;
 wire _20541_;
 wire _20542_;
 wire _20543_;
 wire net2501;
 wire net2500;
 wire net2498;
 wire _20547_;
 wire _20548_;
 wire _20549_;
 wire _20550_;
 wire _20551_;
 wire _20552_;
 wire _20553_;
 wire _20554_;
 wire _20555_;
 wire _20556_;
 wire _20557_;
 wire _20558_;
 wire _20559_;
 wire _20560_;
 wire _20561_;
 wire _20562_;
 wire _20563_;
 wire _20564_;
 wire _20565_;
 wire _20566_;
 wire _20567_;
 wire _20568_;
 wire _20569_;
 wire _20570_;
 wire _20571_;
 wire _20572_;
 wire net2497;
 wire _20574_;
 wire _20575_;
 wire _20576_;
 wire _20577_;
 wire _20578_;
 wire _20579_;
 wire _20580_;
 wire _20581_;
 wire _20582_;
 wire _20583_;
 wire _20584_;
 wire _20585_;
 wire _20586_;
 wire _20587_;
 wire _20588_;
 wire _20589_;
 wire _20590_;
 wire _20591_;
 wire _20592_;
 wire _20593_;
 wire _20594_;
 wire _20595_;
 wire _20596_;
 wire _20597_;
 wire _20598_;
 wire _20599_;
 wire net2495;
 wire _20601_;
 wire _20602_;
 wire _20603_;
 wire _20604_;
 wire _20605_;
 wire _20606_;
 wire net2493;
 wire _20608_;
 wire _20609_;
 wire _20610_;
 wire _20611_;
 wire _20612_;
 wire _20613_;
 wire _20614_;
 wire _20615_;
 wire _20616_;
 wire _20617_;
 wire _20618_;
 wire _20619_;
 wire _20620_;
 wire _20621_;
 wire _20622_;
 wire _20623_;
 wire _20624_;
 wire _20625_;
 wire _20626_;
 wire _20627_;
 wire _20628_;
 wire net2492;
 wire _20630_;
 wire _20631_;
 wire net2490;
 wire net2489;
 wire _20634_;
 wire _20635_;
 wire _20636_;
 wire _20637_;
 wire _20638_;
 wire _20639_;
 wire _20640_;
 wire _20641_;
 wire _20642_;
 wire _20643_;
 wire _20644_;
 wire net2488;
 wire _20646_;
 wire net2487;
 wire _20648_;
 wire net2486;
 wire _20650_;
 wire _20651_;
 wire _20652_;
 wire _20653_;
 wire _20654_;
 wire _20655_;
 wire _20656_;
 wire _20657_;
 wire _20658_;
 wire _20659_;
 wire _20660_;
 wire _20661_;
 wire _20662_;
 wire _20663_;
 wire _20664_;
 wire net2485;
 wire _20666_;
 wire _20667_;
 wire _20668_;
 wire _20669_;
 wire _20670_;
 wire net2484;
 wire _20672_;
 wire _20673_;
 wire _20674_;
 wire _20675_;
 wire _20676_;
 wire _20677_;
 wire _20678_;
 wire _20679_;
 wire _20680_;
 wire net2482;
 wire _20682_;
 wire _20683_;
 wire _20684_;
 wire _20685_;
 wire _20686_;
 wire _20687_;
 wire _20688_;
 wire _20689_;
 wire _20690_;
 wire net2481;
 wire _20692_;
 wire _20693_;
 wire _20694_;
 wire _20695_;
 wire _20696_;
 wire _20697_;
 wire _20698_;
 wire _20699_;
 wire _20700_;
 wire net2480;
 wire _20702_;
 wire net2479;
 wire _20704_;
 wire _20705_;
 wire _20706_;
 wire _20707_;
 wire _20708_;
 wire _20709_;
 wire _20710_;
 wire net2478;
 wire net2477;
 wire _20713_;
 wire _20714_;
 wire _20715_;
 wire _20716_;
 wire _20717_;
 wire _20718_;
 wire _20719_;
 wire _20720_;
 wire _20721_;
 wire _20722_;
 wire _20723_;
 wire net2476;
 wire _20725_;
 wire _20726_;
 wire _20727_;
 wire _20728_;
 wire _20729_;
 wire _20730_;
 wire _20731_;
 wire net2475;
 wire _20733_;
 wire _20734_;
 wire _20735_;
 wire _20736_;
 wire _20737_;
 wire _20738_;
 wire _20739_;
 wire _20740_;
 wire _20741_;
 wire _20742_;
 wire _20743_;
 wire _20744_;
 wire _20745_;
 wire _20746_;
 wire _20747_;
 wire _20748_;
 wire _20749_;
 wire _20750_;
 wire _20751_;
 wire _20752_;
 wire _20753_;
 wire _20754_;
 wire _20755_;
 wire _20756_;
 wire net2473;
 wire _20758_;
 wire _20759_;
 wire _20760_;
 wire _20761_;
 wire _20762_;
 wire _20763_;
 wire _20764_;
 wire _20765_;
 wire _20766_;
 wire _20767_;
 wire _20768_;
 wire _20769_;
 wire net2471;
 wire _20771_;
 wire _20772_;
 wire _20773_;
 wire _20774_;
 wire _20775_;
 wire _20776_;
 wire net2470;
 wire _20778_;
 wire _20779_;
 wire _20780_;
 wire _20781_;
 wire _20782_;
 wire _20783_;
 wire _20784_;
 wire _20785_;
 wire _20786_;
 wire _20787_;
 wire _20788_;
 wire _20789_;
 wire _20790_;
 wire _20791_;
 wire _20792_;
 wire _20793_;
 wire _20794_;
 wire net2469;
 wire _20796_;
 wire _20797_;
 wire _20798_;
 wire _20799_;
 wire _20800_;
 wire _20801_;
 wire _20802_;
 wire _20803_;
 wire _20804_;
 wire _20805_;
 wire _20806_;
 wire _20807_;
 wire _20808_;
 wire _20809_;
 wire _20810_;
 wire _20811_;
 wire _20812_;
 wire net2468;
 wire net2466;
 wire net2465;
 wire _20816_;
 wire _20817_;
 wire _20818_;
 wire _20819_;
 wire _20820_;
 wire net2464;
 wire _20822_;
 wire _20823_;
 wire _20824_;
 wire _20825_;
 wire _20826_;
 wire _20827_;
 wire _20828_;
 wire _20829_;
 wire _20830_;
 wire _20831_;
 wire _20832_;
 wire _20833_;
 wire _20834_;
 wire _20835_;
 wire _20836_;
 wire _20837_;
 wire _20838_;
 wire _20839_;
 wire _20840_;
 wire _20841_;
 wire _20842_;
 wire _20843_;
 wire _20844_;
 wire _20845_;
 wire _20846_;
 wire _20847_;
 wire _20848_;
 wire _20849_;
 wire _20850_;
 wire _20851_;
 wire _20852_;
 wire _20853_;
 wire _20854_;
 wire _20855_;
 wire _20856_;
 wire _20857_;
 wire _20858_;
 wire _20859_;
 wire _20860_;
 wire _20861_;
 wire _20862_;
 wire _20863_;
 wire _20864_;
 wire _20865_;
 wire _20866_;
 wire _20867_;
 wire _20868_;
 wire _20869_;
 wire _20870_;
 wire _20871_;
 wire _20872_;
 wire _20873_;
 wire _20874_;
 wire _20875_;
 wire _20876_;
 wire _20877_;
 wire _20878_;
 wire _20879_;
 wire _20880_;
 wire _20881_;
 wire _20882_;
 wire _20883_;
 wire _20884_;
 wire _20885_;
 wire _20886_;
 wire _20887_;
 wire _20888_;
 wire _20889_;
 wire _20890_;
 wire _20891_;
 wire _20892_;
 wire _20893_;
 wire _20894_;
 wire _20895_;
 wire _20896_;
 wire _20897_;
 wire _20898_;
 wire _20899_;
 wire _20900_;
 wire _20901_;
 wire _20902_;
 wire _20903_;
 wire _20904_;
 wire _20905_;
 wire _20906_;
 wire _20907_;
 wire _20908_;
 wire _20909_;
 wire _20910_;
 wire _20911_;
 wire _20912_;
 wire _20913_;
 wire _20914_;
 wire _20915_;
 wire _20916_;
 wire _20917_;
 wire _20918_;
 wire _20919_;
 wire _20920_;
 wire _20921_;
 wire _20922_;
 wire _20923_;
 wire _20924_;
 wire _20925_;
 wire _20926_;
 wire _20927_;
 wire _20928_;
 wire _20929_;
 wire _20930_;
 wire _20931_;
 wire _20932_;
 wire _20933_;
 wire _20934_;
 wire _20935_;
 wire _20936_;
 wire _20937_;
 wire _20938_;
 wire _20939_;
 wire _20940_;
 wire _20941_;
 wire _20942_;
 wire _20943_;
 wire _20944_;
 wire _20945_;
 wire _20946_;
 wire _20947_;
 wire _20948_;
 wire _20949_;
 wire _20950_;
 wire _20951_;
 wire _20952_;
 wire _20953_;
 wire _20954_;
 wire _20955_;
 wire _20956_;
 wire _20957_;
 wire _20958_;
 wire _20959_;
 wire _20960_;
 wire _20961_;
 wire _20962_;
 wire _20963_;
 wire _20964_;
 wire _20965_;
 wire _20966_;
 wire _20967_;
 wire _20968_;
 wire _20969_;
 wire _20970_;
 wire _20971_;
 wire _20972_;
 wire _20973_;
 wire _20974_;
 wire _20975_;
 wire _20976_;
 wire _20977_;
 wire _20978_;
 wire _20979_;
 wire _20980_;
 wire _20981_;
 wire _20982_;
 wire _20983_;
 wire _20984_;
 wire _20985_;
 wire _20986_;
 wire _20987_;
 wire _20988_;
 wire _20989_;
 wire _20990_;
 wire _20991_;
 wire _20992_;
 wire _20993_;
 wire _20994_;
 wire _20995_;
 wire _20996_;
 wire _20997_;
 wire _20998_;
 wire _20999_;
 wire _21000_;
 wire _21001_;
 wire _21002_;
 wire _21003_;
 wire _21004_;
 wire _21005_;
 wire _21006_;
 wire _21007_;
 wire _21008_;
 wire _21009_;
 wire _21010_;
 wire _21011_;
 wire _21012_;
 wire _21013_;
 wire _21014_;
 wire _21015_;
 wire _21016_;
 wire _21017_;
 wire _21018_;
 wire _21019_;
 wire _21020_;
 wire _21021_;
 wire _21022_;
 wire _21023_;
 wire _21024_;
 wire _21025_;
 wire _21026_;
 wire _21027_;
 wire _21028_;
 wire _21029_;
 wire _21030_;
 wire _21031_;
 wire _21032_;
 wire _21033_;
 wire _21034_;
 wire _21035_;
 wire _21036_;
 wire _21037_;
 wire _21038_;
 wire _21039_;
 wire _21040_;
 wire _21041_;
 wire _21042_;
 wire _21043_;
 wire _21044_;
 wire _21045_;
 wire _21046_;
 wire _21047_;
 wire _21048_;
 wire _21049_;
 wire _21050_;
 wire _21051_;
 wire _21052_;
 wire _21053_;
 wire _21054_;
 wire _21055_;
 wire _21056_;
 wire _21057_;
 wire _21058_;
 wire _21059_;
 wire _21060_;
 wire _21061_;
 wire _21062_;
 wire _21063_;
 wire _21064_;
 wire _21065_;
 wire _21066_;
 wire _21067_;
 wire _21068_;
 wire _21069_;
 wire _21070_;
 wire _21071_;
 wire _21072_;
 wire _21073_;
 wire _21074_;
 wire _21075_;
 wire _21076_;
 wire _21077_;
 wire _21078_;
 wire _21079_;
 wire _21080_;
 wire _21081_;
 wire _21082_;
 wire _21083_;
 wire _21084_;
 wire _21085_;
 wire _21086_;
 wire _21087_;
 wire _21088_;
 wire _21089_;
 wire _21090_;
 wire _21091_;
 wire _21092_;
 wire _21093_;
 wire _21094_;
 wire _21095_;
 wire _21096_;
 wire _21097_;
 wire _21098_;
 wire _21099_;
 wire _21100_;
 wire _21101_;
 wire _21102_;
 wire _21103_;
 wire _21104_;
 wire _21105_;
 wire _21106_;
 wire _21107_;
 wire _21108_;
 wire _21109_;
 wire _21110_;
 wire _21111_;
 wire _21112_;
 wire _21113_;
 wire _21114_;
 wire _21115_;
 wire _21116_;
 wire _21117_;
 wire _21118_;
 wire _21119_;
 wire _21120_;
 wire _21121_;
 wire _21122_;
 wire _21123_;
 wire _21124_;
 wire _21125_;
 wire _21126_;
 wire _21127_;
 wire _21128_;
 wire _21129_;
 wire _21130_;
 wire _21131_;
 wire _21132_;
 wire _21133_;
 wire _21134_;
 wire _21135_;
 wire _21136_;
 wire _21137_;
 wire _21138_;
 wire _21139_;
 wire _21140_;
 wire _21141_;
 wire _21142_;
 wire _21143_;
 wire _21144_;
 wire _21145_;
 wire _21146_;
 wire _21147_;
 wire _21148_;
 wire _21149_;
 wire _21150_;
 wire _21151_;
 wire _21152_;
 wire _21153_;
 wire _21154_;
 wire _21155_;
 wire _21156_;
 wire _21157_;
 wire _21158_;
 wire _21159_;
 wire _21160_;
 wire _21161_;
 wire _21162_;
 wire _21163_;
 wire _21164_;
 wire _21165_;
 wire _21166_;
 wire _21167_;
 wire _21168_;
 wire _21169_;
 wire _21170_;
 wire _21171_;
 wire _21172_;
 wire _21173_;
 wire _21174_;
 wire _21175_;
 wire _21176_;
 wire _21177_;
 wire _21178_;
 wire _21179_;
 wire _21180_;
 wire _21181_;
 wire _21182_;
 wire _21183_;
 wire _21184_;
 wire _21185_;
 wire _21186_;
 wire _21187_;
 wire _21188_;
 wire _21189_;
 wire _21190_;
 wire _21191_;
 wire _21192_;
 wire _21193_;
 wire _21194_;
 wire _21195_;
 wire _21196_;
 wire _21197_;
 wire _21198_;
 wire _21199_;
 wire _21200_;
 wire _21201_;
 wire _21202_;
 wire _21203_;
 wire _21204_;
 wire _21205_;
 wire _21206_;
 wire _21207_;
 wire _21208_;
 wire _21209_;
 wire _21210_;
 wire _21211_;
 wire _21212_;
 wire _21213_;
 wire _21214_;
 wire _21215_;
 wire _21216_;
 wire _21217_;
 wire _21218_;
 wire _21219_;
 wire _21220_;
 wire _21221_;
 wire _21222_;
 wire _21223_;
 wire _21224_;
 wire _21225_;
 wire _21226_;
 wire _21227_;
 wire _21228_;
 wire _21229_;
 wire _21230_;
 wire _21231_;
 wire _21232_;
 wire _21233_;
 wire _21234_;
 wire _21235_;
 wire _21236_;
 wire _21237_;
 wire _21238_;
 wire _21239_;
 wire _21240_;
 wire _21241_;
 wire _21242_;
 wire _21243_;
 wire _21244_;
 wire _21245_;
 wire _21246_;
 wire _21247_;
 wire _21248_;
 wire _21249_;
 wire _21250_;
 wire _21251_;
 wire _21252_;
 wire _21253_;
 wire _21254_;
 wire _21255_;
 wire _21256_;
 wire _21257_;
 wire _21258_;
 wire _21259_;
 wire _21260_;
 wire _21261_;
 wire _21262_;
 wire _21263_;
 wire _21264_;
 wire _21265_;
 wire _21266_;
 wire _21267_;
 wire _21268_;
 wire _21269_;
 wire _21270_;
 wire _21271_;
 wire _21272_;
 wire _21273_;
 wire _21274_;
 wire _21275_;
 wire _21276_;
 wire _21277_;
 wire _21278_;
 wire _21279_;
 wire _21280_;
 wire _21281_;
 wire _21282_;
 wire _21283_;
 wire _21284_;
 wire _21285_;
 wire _21286_;
 wire _21287_;
 wire _21288_;
 wire _21289_;
 wire _21290_;
 wire _21291_;
 wire _21292_;
 wire _21293_;
 wire _21294_;
 wire _21295_;
 wire _21296_;
 wire _21297_;
 wire _21298_;
 wire _21299_;
 wire _21300_;
 wire _21301_;
 wire _21302_;
 wire _21303_;
 wire _21304_;
 wire _21305_;
 wire _21306_;
 wire _21307_;
 wire _21308_;
 wire _21309_;
 wire _21310_;
 wire _21311_;
 wire _21312_;
 wire _21313_;
 wire _21314_;
 wire _21315_;
 wire _21316_;
 wire _21317_;
 wire _21318_;
 wire _21319_;
 wire _21320_;
 wire _21321_;
 wire _21322_;
 wire _21323_;
 wire _21324_;
 wire _21325_;
 wire _21326_;
 wire _21327_;
 wire _21328_;
 wire _21329_;
 wire _21330_;
 wire _21331_;
 wire _21332_;
 wire _21333_;
 wire _21334_;
 wire _21335_;
 wire _21336_;
 wire _21337_;
 wire _21338_;
 wire _21339_;
 wire _21340_;
 wire _21341_;
 wire _21342_;
 wire _21343_;
 wire _21344_;
 wire _21345_;
 wire _21346_;
 wire _21347_;
 wire _21348_;
 wire _21349_;
 wire _21350_;
 wire _21351_;
 wire _21352_;
 wire _21353_;
 wire _21354_;
 wire _21355_;
 wire _21356_;
 wire _21357_;
 wire _21358_;
 wire _21359_;
 wire _21360_;
 wire _21361_;
 wire _21362_;
 wire _21363_;
 wire _21364_;
 wire _21365_;
 wire _21366_;
 wire _21367_;
 wire _21368_;
 wire _21369_;
 wire _21370_;
 wire _21371_;
 wire _21372_;
 wire _21373_;
 wire _21374_;
 wire _21375_;
 wire _21376_;
 wire _21377_;
 wire _21378_;
 wire _21379_;
 wire _21380_;
 wire _21381_;
 wire _21382_;
 wire _21383_;
 wire _21384_;
 wire _21385_;
 wire _21386_;
 wire _21387_;
 wire _21388_;
 wire _21389_;
 wire _21390_;
 wire _21391_;
 wire _21392_;
 wire _21393_;
 wire _21394_;
 wire _21395_;
 wire _21396_;
 wire _21397_;
 wire _21398_;
 wire _21399_;
 wire _21400_;
 wire _21401_;
 wire _21402_;
 wire _21403_;
 wire _21404_;
 wire _21405_;
 wire _21406_;
 wire _21407_;
 wire _21408_;
 wire _21409_;
 wire _21410_;
 wire _21411_;
 wire _21412_;
 wire _21413_;
 wire _21414_;
 wire _21415_;
 wire _21416_;
 wire _21417_;
 wire _21418_;
 wire _21419_;
 wire _21420_;
 wire _21421_;
 wire _21422_;
 wire _21423_;
 wire _21424_;
 wire _21425_;
 wire _21426_;
 wire _21427_;
 wire _21428_;
 wire _21429_;
 wire _21430_;
 wire _21431_;
 wire _21432_;
 wire _21433_;
 wire _21434_;
 wire _21435_;
 wire _21436_;
 wire _21437_;
 wire _21438_;
 wire _21439_;
 wire _21440_;
 wire _21441_;
 wire _21442_;
 wire _21443_;
 wire _21444_;
 wire _21445_;
 wire _21446_;
 wire _21447_;
 wire _21448_;
 wire _21449_;
 wire _21450_;
 wire _21451_;
 wire _21452_;
 wire _21453_;
 wire _21454_;
 wire _21455_;
 wire _21456_;
 wire _21457_;
 wire _21458_;
 wire _21459_;
 wire _21460_;
 wire _21461_;
 wire _21462_;
 wire _21463_;
 wire _21464_;
 wire _21465_;
 wire _21466_;
 wire _21467_;
 wire _21468_;
 wire _21469_;
 wire _21470_;
 wire _21471_;
 wire _21472_;
 wire _21473_;
 wire _21474_;
 wire _21475_;
 wire _21476_;
 wire _21477_;
 wire _21478_;
 wire _21479_;
 wire _21480_;
 wire _21481_;
 wire _21482_;
 wire _21483_;
 wire _21484_;
 wire _21485_;
 wire _21486_;
 wire _21487_;
 wire _21488_;
 wire _21489_;
 wire _21490_;
 wire _21491_;
 wire _21492_;
 wire _21493_;
 wire _21494_;
 wire _21495_;
 wire _21496_;
 wire _21497_;
 wire _21498_;
 wire _21499_;
 wire _21500_;
 wire _21501_;
 wire _21502_;
 wire _21503_;
 wire _21504_;
 wire _21505_;
 wire _21506_;
 wire _21507_;
 wire _21508_;
 wire _21509_;
 wire _21510_;
 wire _21511_;
 wire _21512_;
 wire _21513_;
 wire _21514_;
 wire _21515_;
 wire _21516_;
 wire _21517_;
 wire _21518_;
 wire _21519_;
 wire _21520_;
 wire _21521_;
 wire _21522_;
 wire _21523_;
 wire _21524_;
 wire _21525_;
 wire _21526_;
 wire _21527_;
 wire _21528_;
 wire _21529_;
 wire _21530_;
 wire _21531_;
 wire _21532_;
 wire _21533_;
 wire _21534_;
 wire _21535_;
 wire _21536_;
 wire _21537_;
 wire _21538_;
 wire _21539_;
 wire _21540_;
 wire _21541_;
 wire _21542_;
 wire _21543_;
 wire _21544_;
 wire _21545_;
 wire _21546_;
 wire _21547_;
 wire _21548_;
 wire _21549_;
 wire _21550_;
 wire _21551_;
 wire _21552_;
 wire _21553_;
 wire _21554_;
 wire _21555_;
 wire _21556_;
 wire _21557_;
 wire _21558_;
 wire _21559_;
 wire _21560_;
 wire _21561_;
 wire _21562_;
 wire _21563_;
 wire _21564_;
 wire _21565_;
 wire _21566_;
 wire _21567_;
 wire _21568_;
 wire _21569_;
 wire _21570_;
 wire _21571_;
 wire _21572_;
 wire _21573_;
 wire _21574_;
 wire _21575_;
 wire _21576_;
 wire _21577_;
 wire _21578_;
 wire _21579_;
 wire _21580_;
 wire _21581_;
 wire _21582_;
 wire _21583_;
 wire _21584_;
 wire _21585_;
 wire _21586_;
 wire _21587_;
 wire _21588_;
 wire _21589_;
 wire _21590_;
 wire _21591_;
 wire _21592_;
 wire _21593_;
 wire _21594_;
 wire _21595_;
 wire _21596_;
 wire _21597_;
 wire _21598_;
 wire _21599_;
 wire _21600_;
 wire _21601_;
 wire _21602_;
 wire _21603_;
 wire _21604_;
 wire _21605_;
 wire _21606_;
 wire _21607_;
 wire _21608_;
 wire _21609_;
 wire _21610_;
 wire _21611_;
 wire _21612_;
 wire _21613_;
 wire _21614_;
 wire _21615_;
 wire _21616_;
 wire _21617_;
 wire _21618_;
 wire _21619_;
 wire _21620_;
 wire _21621_;
 wire _21622_;
 wire _21623_;
 wire _21624_;
 wire _21625_;
 wire _21626_;
 wire _21627_;
 wire _21628_;
 wire _21629_;
 wire _21630_;
 wire _21631_;
 wire _21632_;
 wire _21633_;
 wire _21634_;
 wire _21635_;
 wire _21636_;
 wire _21637_;
 wire _21638_;
 wire _21639_;
 wire _21640_;
 wire _21641_;
 wire _21642_;
 wire _21643_;
 wire _21644_;
 wire _21645_;
 wire _21646_;
 wire _21647_;
 wire _21648_;
 wire _21649_;
 wire _21650_;
 wire _21651_;
 wire _21652_;
 wire _21653_;
 wire _21654_;
 wire _21655_;
 wire _21656_;
 wire _21657_;
 wire _21658_;
 wire _21659_;
 wire _21660_;
 wire _21661_;
 wire _21662_;
 wire _21663_;
 wire _21664_;
 wire _21665_;
 wire _21666_;
 wire _21667_;
 wire _21668_;
 wire _21669_;
 wire _21670_;
 wire _21671_;
 wire _21672_;
 wire _21673_;
 wire _21674_;
 wire _21675_;
 wire _21676_;
 wire _21677_;
 wire _21678_;
 wire _21679_;
 wire _21680_;
 wire _21681_;
 wire _21682_;
 wire _21683_;
 wire _21684_;
 wire _21685_;
 wire _21686_;
 wire _21687_;
 wire _21688_;
 wire _21689_;
 wire _21690_;
 wire _21691_;
 wire _21692_;
 wire _21693_;
 wire _21694_;
 wire _21695_;
 wire _21696_;
 wire _21697_;
 wire _21698_;
 wire _21699_;
 wire _21700_;
 wire _21701_;
 wire _21702_;
 wire _21703_;
 wire _21704_;
 wire _21705_;
 wire _21706_;
 wire _21707_;
 wire _21708_;
 wire _21709_;
 wire _21710_;
 wire _21711_;
 wire _21712_;
 wire _21713_;
 wire _21714_;
 wire _21715_;
 wire _21716_;
 wire _21717_;
 wire _21718_;
 wire _21719_;
 wire _21720_;
 wire _21721_;
 wire _21722_;
 wire _21723_;
 wire _21724_;
 wire _21725_;
 wire _21726_;
 wire _21727_;
 wire _21728_;
 wire _21729_;
 wire _21730_;
 wire _21731_;
 wire _21732_;
 wire _21733_;
 wire _21734_;
 wire _21735_;
 wire _21736_;
 wire _21737_;
 wire _21738_;
 wire _21739_;
 wire _21740_;
 wire _21741_;
 wire _21742_;
 wire _21743_;
 wire _21744_;
 wire _21745_;
 wire _21746_;
 wire _21747_;
 wire _21748_;
 wire _21749_;
 wire _21750_;
 wire _21751_;
 wire _21752_;
 wire _21753_;
 wire _21754_;
 wire _21755_;
 wire _21756_;
 wire _21757_;
 wire _21758_;
 wire _21759_;
 wire _21760_;
 wire _21761_;
 wire _21762_;
 wire _21763_;
 wire _21764_;
 wire _21765_;
 wire _21766_;
 wire _21767_;
 wire _21768_;
 wire _21769_;
 wire _21770_;
 wire _21771_;
 wire _21772_;
 wire _21773_;
 wire _21774_;
 wire _21775_;
 wire _21776_;
 wire _21777_;
 wire _21778_;
 wire _21779_;
 wire _21780_;
 wire _21781_;
 wire _21782_;
 wire _21783_;
 wire _21784_;
 wire _21785_;
 wire _21786_;
 wire _21787_;
 wire _21788_;
 wire _21789_;
 wire _21790_;
 wire _21791_;
 wire _21792_;
 wire _21793_;
 wire _21794_;
 wire _21795_;
 wire _21796_;
 wire _21797_;
 wire _21798_;
 wire _21799_;
 wire _21800_;
 wire _21801_;
 wire _21802_;
 wire _21803_;
 wire _21804_;
 wire _21805_;
 wire _21806_;
 wire _21807_;
 wire _21808_;
 wire _21809_;
 wire _21810_;
 wire _21811_;
 wire _21812_;
 wire _21813_;
 wire _21814_;
 wire _21815_;
 wire _21816_;
 wire _21817_;
 wire _21818_;
 wire _21819_;
 wire _21820_;
 wire _21821_;
 wire _21822_;
 wire _21823_;
 wire _21824_;
 wire _21825_;
 wire _21826_;
 wire _21827_;
 wire _21828_;
 wire _21829_;
 wire _21830_;
 wire _21831_;
 wire _21832_;
 wire _21833_;
 wire _21834_;
 wire _21835_;
 wire _21836_;
 wire _21837_;
 wire _21838_;
 wire _21839_;
 wire _21840_;
 wire _21841_;
 wire _21842_;
 wire _21843_;
 wire _21844_;
 wire _21845_;
 wire _21846_;
 wire _21847_;
 wire _21848_;
 wire _21849_;
 wire _21850_;
 wire _21851_;
 wire _21852_;
 wire _21853_;
 wire _21854_;
 wire _21855_;
 wire _21856_;
 wire _21857_;
 wire _21858_;
 wire _21859_;
 wire _21860_;
 wire _21861_;
 wire _21862_;
 wire _21863_;
 wire _21864_;
 wire _21865_;
 wire _21866_;
 wire _21867_;
 wire _21868_;
 wire _21869_;
 wire _21870_;
 wire _21871_;
 wire _21872_;
 wire _21873_;
 wire _21874_;
 wire _21875_;
 wire _21876_;
 wire _21877_;
 wire _21878_;
 wire _21879_;
 wire _21880_;
 wire _21881_;
 wire _21882_;
 wire _21883_;
 wire _21884_;
 wire _21885_;
 wire _21886_;
 wire _21887_;
 wire _21888_;
 wire _21889_;
 wire _21890_;
 wire _21891_;
 wire _21892_;
 wire _21893_;
 wire _21894_;
 wire _21895_;
 wire _21896_;
 wire _21897_;
 wire _21898_;
 wire _21899_;
 wire _21900_;
 wire _21901_;
 wire _21902_;
 wire _21903_;
 wire _21904_;
 wire _21905_;
 wire _21906_;
 wire _21907_;
 wire _21908_;
 wire _21909_;
 wire _21910_;
 wire _21911_;
 wire _21912_;
 wire _21913_;
 wire _21914_;
 wire _21915_;
 wire _21916_;
 wire _21917_;
 wire _21918_;
 wire _21919_;
 wire _21920_;
 wire _21921_;
 wire _21922_;
 wire _21923_;
 wire _21924_;
 wire _21925_;
 wire _21926_;
 wire _21927_;
 wire _21928_;
 wire _21929_;
 wire _21930_;
 wire _21931_;
 wire _21932_;
 wire _21933_;
 wire _21934_;
 wire _21935_;
 wire _21936_;
 wire _21937_;
 wire _21938_;
 wire _21939_;
 wire _21940_;
 wire _21941_;
 wire _21942_;
 wire _21943_;
 wire _21944_;
 wire _21945_;
 wire _21946_;
 wire _21947_;
 wire _21948_;
 wire _21949_;
 wire _21950_;
 wire _21951_;
 wire _21952_;
 wire _21953_;
 wire _21954_;
 wire _21955_;
 wire _21956_;
 wire _21957_;
 wire _21958_;
 wire _21959_;
 wire _21960_;
 wire _21961_;
 wire _21962_;
 wire _21963_;
 wire _21964_;
 wire _21965_;
 wire _21966_;
 wire _21967_;
 wire _21968_;
 wire _21969_;
 wire _21970_;
 wire _21971_;
 wire _21972_;
 wire _21973_;
 wire _21974_;
 wire _21975_;
 wire _21976_;
 wire _21977_;
 wire _21978_;
 wire _21979_;
 wire _21980_;
 wire _21981_;
 wire _21982_;
 wire _21983_;
 wire _21984_;
 wire _21985_;
 wire _21986_;
 wire _21987_;
 wire _21988_;
 wire _21989_;
 wire _21990_;
 wire _21991_;
 wire _21992_;
 wire _21993_;
 wire _21994_;
 wire _21995_;
 wire _21996_;
 wire _21997_;
 wire _21998_;
 wire _21999_;
 wire _22000_;
 wire _22001_;
 wire _22002_;
 wire _22003_;
 wire _22004_;
 wire _22005_;
 wire _22006_;
 wire _22007_;
 wire _22008_;
 wire _22009_;
 wire _22010_;
 wire _22011_;
 wire _22012_;
 wire _22013_;
 wire _22014_;
 wire _22015_;
 wire _22016_;
 wire _22017_;
 wire _22018_;
 wire _22019_;
 wire _22020_;
 wire _22021_;
 wire _22022_;
 wire _22023_;
 wire _22024_;
 wire _22025_;
 wire _22026_;
 wire _22027_;
 wire _22028_;
 wire _22029_;
 wire _22030_;
 wire _22031_;
 wire _22032_;
 wire _22033_;
 wire _22034_;
 wire _22035_;
 wire _22036_;
 wire _22037_;
 wire _22038_;
 wire _22039_;
 wire _22040_;
 wire _22041_;
 wire _22042_;
 wire _22043_;
 wire _22044_;
 wire _22045_;
 wire _22046_;
 wire _22047_;
 wire _22048_;
 wire _22049_;
 wire _22050_;
 wire _22051_;
 wire _22052_;
 wire _22053_;
 wire _22054_;
 wire _22055_;
 wire _22056_;
 wire _22057_;
 wire _22058_;
 wire _22059_;
 wire _22060_;
 wire _22061_;
 wire _22062_;
 wire _22063_;
 wire _22064_;
 wire _22065_;
 wire _22066_;
 wire _22067_;
 wire _22068_;
 wire _22069_;
 wire _22070_;
 wire _22071_;
 wire _22072_;
 wire _22073_;
 wire _22074_;
 wire _22075_;
 wire _22076_;
 wire _22077_;
 wire _22078_;
 wire _22079_;
 wire _22080_;
 wire _22081_;
 wire _22082_;
 wire _22083_;
 wire _22084_;
 wire _22085_;
 wire _22086_;
 wire _22087_;
 wire _22088_;
 wire _22089_;
 wire _22090_;
 wire _22091_;
 wire _22092_;
 wire _22093_;
 wire _22094_;
 wire _22095_;
 wire _22096_;
 wire _22097_;
 wire _22098_;
 wire _22099_;
 wire _22100_;
 wire _22101_;
 wire _22102_;
 wire _22103_;
 wire _22104_;
 wire _22105_;
 wire _22106_;
 wire _22107_;
 wire _22108_;
 wire _22109_;
 wire _22110_;
 wire _22111_;
 wire _22112_;
 wire _22113_;
 wire _22114_;
 wire _22115_;
 wire _22116_;
 wire _22117_;
 wire _22118_;
 wire _22119_;
 wire _22120_;
 wire _22121_;
 wire _22122_;
 wire _22123_;
 wire _22124_;
 wire _22125_;
 wire _22126_;
 wire _22127_;
 wire _22128_;
 wire _22129_;
 wire _22130_;
 wire _22131_;
 wire _22132_;
 wire _22133_;
 wire _22134_;
 wire _22135_;
 wire _22136_;
 wire _22137_;
 wire _22138_;
 wire _22139_;
 wire _22140_;
 wire _22141_;
 wire _22142_;
 wire _22143_;
 wire _22144_;
 wire _22145_;
 wire _22146_;
 wire _22147_;
 wire _22148_;
 wire _22149_;
 wire _22150_;
 wire _22151_;
 wire _22152_;
 wire _22153_;
 wire _22154_;
 wire _22155_;
 wire _22156_;
 wire _22157_;
 wire _22158_;
 wire _22159_;
 wire _22160_;
 wire _22161_;
 wire _22162_;
 wire _22163_;
 wire _22164_;
 wire _22165_;
 wire _22166_;
 wire _22167_;
 wire _22168_;
 wire _22169_;
 wire _22170_;
 wire _22171_;
 wire _22172_;
 wire _22173_;
 wire _22174_;
 wire _22175_;
 wire _22176_;
 wire _22177_;
 wire _22178_;
 wire _22179_;
 wire _22180_;
 wire _22181_;
 wire _22182_;
 wire _22183_;
 wire _22184_;
 wire _22185_;
 wire _22186_;
 wire _22187_;
 wire _22188_;
 wire _22189_;
 wire _22190_;
 wire _22191_;
 wire _22192_;
 wire _22193_;
 wire _22194_;
 wire _22195_;
 wire _22196_;
 wire _22197_;
 wire _22198_;
 wire _22199_;
 wire _22200_;
 wire _22201_;
 wire _22202_;
 wire _22203_;
 wire _22204_;
 wire _22205_;
 wire _22206_;
 wire _22207_;
 wire _22208_;
 wire _22209_;
 wire _22210_;
 wire _22211_;
 wire _22212_;
 wire _22213_;
 wire _22214_;
 wire _22215_;
 wire _22216_;
 wire _22217_;
 wire _22218_;
 wire _22219_;
 wire _22220_;
 wire _22221_;
 wire _22222_;
 wire _22223_;
 wire _22224_;
 wire _22225_;
 wire _22226_;
 wire _22227_;
 wire _22228_;
 wire _22229_;
 wire _22230_;
 wire _22231_;
 wire _22232_;
 wire _22233_;
 wire _22234_;
 wire _22235_;
 wire _22236_;
 wire _22237_;
 wire _22238_;
 wire _22239_;
 wire _22240_;
 wire _22241_;
 wire _22242_;
 wire _22243_;
 wire _22244_;
 wire _22245_;
 wire _22246_;
 wire _22247_;
 wire _22248_;
 wire _22249_;
 wire _22250_;
 wire _22251_;
 wire _22252_;
 wire _22253_;
 wire _22254_;
 wire _22255_;
 wire _22256_;
 wire _22257_;
 wire _22258_;
 wire _22259_;
 wire _22260_;
 wire _22261_;
 wire _22262_;
 wire _22263_;
 wire _22264_;
 wire _22265_;
 wire _22266_;
 wire _22267_;
 wire _22268_;
 wire _22269_;
 wire _22270_;
 wire _22271_;
 wire _22272_;
 wire _22273_;
 wire _22274_;
 wire _22275_;
 wire _22276_;
 wire _22277_;
 wire _22278_;
 wire _22279_;
 wire _22280_;
 wire _22281_;
 wire _22282_;
 wire _22283_;
 wire _22284_;
 wire _22285_;
 wire _22286_;
 wire _22287_;
 wire _22288_;
 wire _22289_;
 wire _22290_;
 wire _22291_;
 wire _22292_;
 wire _22293_;
 wire _22294_;
 wire _22295_;
 wire _22296_;
 wire _22297_;
 wire _22298_;
 wire _22299_;
 wire _22300_;
 wire _22301_;
 wire _22302_;
 wire _22303_;
 wire _22304_;
 wire _22305_;
 wire _22306_;
 wire _22307_;
 wire _22308_;
 wire _22309_;
 wire _22310_;
 wire _22311_;
 wire _22312_;
 wire _22313_;
 wire _22314_;
 wire _22315_;
 wire _22316_;
 wire _22317_;
 wire _22318_;
 wire _22319_;
 wire _22320_;
 wire _22321_;
 wire _22322_;
 wire _22323_;
 wire _22324_;
 wire _22325_;
 wire _22326_;
 wire _22327_;
 wire _22328_;
 wire _22329_;
 wire _22330_;
 wire _22331_;
 wire _22332_;
 wire _22333_;
 wire _22334_;
 wire _22335_;
 wire _22336_;
 wire _22337_;
 wire _22338_;
 wire _22339_;
 wire _22340_;
 wire _22341_;
 wire _22342_;
 wire _22343_;
 wire _22344_;
 wire _22345_;
 wire _22346_;
 wire _22347_;
 wire _22348_;
 wire _22349_;
 wire _22350_;
 wire _22351_;
 wire _22352_;
 wire _22353_;
 wire _22354_;
 wire _22355_;
 wire _22356_;
 wire _22357_;
 wire _22358_;
 wire _22359_;
 wire _22360_;
 wire _22361_;
 wire _22362_;
 wire _22363_;
 wire _22364_;
 wire _22365_;
 wire _22366_;
 wire _22367_;
 wire _22368_;
 wire _22369_;
 wire _22370_;
 wire _22371_;
 wire _22372_;
 wire _22373_;
 wire _22374_;
 wire _22375_;
 wire _22376_;
 wire _22377_;
 wire _22378_;
 wire _22379_;
 wire _22380_;
 wire _22381_;
 wire _22382_;
 wire _22383_;
 wire _22384_;
 wire _22385_;
 wire _22386_;
 wire _22387_;
 wire _22388_;
 wire _22389_;
 wire _22390_;
 wire _22391_;
 wire _22392_;
 wire _22393_;
 wire _22394_;
 wire _22395_;
 wire _22396_;
 wire _22397_;
 wire _22398_;
 wire _22399_;
 wire _22400_;
 wire _22401_;
 wire _22402_;
 wire _22403_;
 wire _22404_;
 wire _22405_;
 wire _22406_;
 wire _22407_;
 wire _22408_;
 wire _22409_;
 wire _22410_;
 wire _22411_;
 wire _22412_;
 wire _22413_;
 wire _22414_;
 wire _22415_;
 wire _22416_;
 wire _22417_;
 wire _22418_;
 wire _22419_;
 wire _22420_;
 wire _22421_;
 wire _22422_;
 wire _22423_;
 wire _22424_;
 wire _22425_;
 wire _22426_;
 wire _22427_;
 wire _22428_;
 wire _22429_;
 wire _22430_;
 wire _22431_;
 wire _22432_;
 wire _22433_;
 wire _22434_;
 wire _22435_;
 wire _22436_;
 wire _22437_;
 wire _22438_;
 wire _22439_;
 wire _22440_;
 wire _22441_;
 wire _22442_;
 wire _22443_;
 wire _22444_;
 wire _22445_;
 wire _22446_;
 wire _22447_;
 wire _22448_;
 wire _22449_;
 wire _22450_;
 wire _22451_;
 wire _22452_;
 wire _22453_;
 wire _22454_;
 wire _22455_;
 wire _22456_;
 wire _22457_;
 wire _22458_;
 wire _22459_;
 wire _22460_;
 wire _22461_;
 wire _22462_;
 wire _22463_;
 wire _22464_;
 wire _22465_;
 wire _22466_;
 wire _22467_;
 wire _22468_;
 wire _22469_;
 wire _22470_;
 wire _22471_;
 wire _22472_;
 wire _22473_;
 wire _22474_;
 wire _22475_;
 wire _22476_;
 wire _22477_;
 wire _22478_;
 wire _22479_;
 wire _22480_;
 wire _22481_;
 wire _22482_;
 wire _22483_;
 wire _22484_;
 wire _22485_;
 wire _22486_;
 wire _22487_;
 wire _22488_;
 wire _22489_;
 wire _22490_;
 wire _22491_;
 wire _22492_;
 wire _22493_;
 wire _22494_;
 wire _22495_;
 wire _22496_;
 wire _22497_;
 wire _22498_;
 wire _22499_;
 wire _22500_;
 wire _22501_;
 wire _22502_;
 wire _22503_;
 wire _22504_;
 wire _22505_;
 wire _22506_;
 wire _22507_;
 wire _22508_;
 wire _22509_;
 wire _22510_;
 wire _22511_;
 wire _22512_;
 wire _22513_;
 wire _22514_;
 wire _22515_;
 wire _22516_;
 wire _22517_;
 wire _22518_;
 wire _22519_;
 wire _22520_;
 wire _22521_;
 wire _22522_;
 wire _22523_;
 wire _22524_;
 wire _22525_;
 wire _22526_;
 wire _22527_;
 wire _22528_;
 wire _22529_;
 wire _22530_;
 wire _22531_;
 wire _22532_;
 wire _22533_;
 wire _22534_;
 wire _22535_;
 wire _22536_;
 wire _22537_;
 wire _22538_;
 wire _22539_;
 wire _22540_;
 wire _22541_;
 wire _22542_;
 wire _22543_;
 wire _22544_;
 wire _22545_;
 wire _22546_;
 wire _22547_;
 wire _22548_;
 wire _22549_;
 wire _22550_;
 wire _22551_;
 wire _22552_;
 wire _22553_;
 wire _22554_;
 wire _22555_;
 wire _22556_;
 wire _22557_;
 wire _22558_;
 wire _22559_;
 wire _22560_;
 wire _22561_;
 wire _22562_;
 wire _22563_;
 wire _22564_;
 wire _22565_;
 wire _22566_;
 wire _22567_;
 wire _22568_;
 wire _22569_;
 wire _22570_;
 wire _22571_;
 wire _22572_;
 wire _22573_;
 wire _22574_;
 wire _22575_;
 wire _22576_;
 wire _22577_;
 wire _22578_;
 wire _22579_;
 wire _22580_;
 wire _22581_;
 wire _22582_;
 wire _22583_;
 wire _22584_;
 wire _22585_;
 wire _22586_;
 wire _22587_;
 wire _22588_;
 wire _22589_;
 wire _22590_;
 wire _22591_;
 wire _22592_;
 wire _22593_;
 wire _22594_;
 wire _22595_;
 wire _22596_;
 wire _22597_;
 wire _22598_;
 wire _22599_;
 wire _22600_;
 wire _22601_;
 wire _22602_;
 wire _22603_;
 wire _22604_;
 wire _22605_;
 wire _22606_;
 wire _22607_;
 wire _22608_;
 wire _22609_;
 wire _22610_;
 wire _22611_;
 wire _22612_;
 wire _22613_;
 wire _22614_;
 wire _22615_;
 wire _22616_;
 wire _22617_;
 wire _22618_;
 wire _22619_;
 wire _22620_;
 wire _22621_;
 wire _22622_;
 wire _22623_;
 wire _22624_;
 wire _22625_;
 wire _22626_;
 wire _22627_;
 wire _22628_;
 wire _22629_;
 wire _22630_;
 wire _22631_;
 wire _22632_;
 wire _22633_;
 wire _22634_;
 wire _22635_;
 wire _22636_;
 wire _22637_;
 wire _22638_;
 wire _22639_;
 wire _22640_;
 wire _22641_;
 wire _22642_;
 wire net2636;
 wire net969;
 wire clk_in;
 assign clk_in = gpio_in[38];
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net680;
 wire net703;
 wire net702;
 wire net701;
 wire net700;
 wire net679;
 wire net697;
 wire net696;
 wire net695;
 wire net694;
 wire net693;
 wire net692;
 wire net678;
 wire net691;
 wire net690;
 wire net677;
 wire net724;
 wire net723;
 wire net741;
 wire net740;
 wire net739;
 wire net738;
 wire net737;
 wire net736;
 wire net722;
 wire net735;
 wire net734;
 wire net721;
 wire net660;
 wire \inst$top.i$88 ;
 wire \inst$top.rst_n_sync.rst ;
 wire \inst$top.rst_n_sync.stage0 ;
 wire \inst$top.soc.bus__addr[2] ;
 wire \inst$top.soc.bus__addr[3] ;
 wire \inst$top.soc.bus__adr[2] ;
 wire \inst$top.soc.bus__adr[3] ;
 wire \inst$top.soc.bus__adr[4] ;
 wire \inst$top.soc.bus__adr[5] ;
 wire \inst$top.soc.bus__adr[6] ;
 wire \inst$top.soc.bus__adr[7] ;
 wire \inst$top.soc.bus__dat_w[0] ;
 wire \inst$top.soc.bus__dat_w[10] ;
 wire \inst$top.soc.bus__dat_w[11] ;
 wire \inst$top.soc.bus__dat_w[12] ;
 wire \inst$top.soc.bus__dat_w[13] ;
 wire \inst$top.soc.bus__dat_w[14] ;
 wire \inst$top.soc.bus__dat_w[15] ;
 wire \inst$top.soc.bus__dat_w[16] ;
 wire \inst$top.soc.bus__dat_w[17] ;
 wire \inst$top.soc.bus__dat_w[18] ;
 wire \inst$top.soc.bus__dat_w[19] ;
 wire \inst$top.soc.bus__dat_w[1] ;
 wire \inst$top.soc.bus__dat_w[20] ;
 wire \inst$top.soc.bus__dat_w[21] ;
 wire \inst$top.soc.bus__dat_w[22] ;
 wire \inst$top.soc.bus__dat_w[23] ;
 wire \inst$top.soc.bus__dat_w[24] ;
 wire \inst$top.soc.bus__dat_w[25] ;
 wire \inst$top.soc.bus__dat_w[26] ;
 wire \inst$top.soc.bus__dat_w[27] ;
 wire \inst$top.soc.bus__dat_w[28] ;
 wire \inst$top.soc.bus__dat_w[29] ;
 wire \inst$top.soc.bus__dat_w[2] ;
 wire \inst$top.soc.bus__dat_w[30] ;
 wire \inst$top.soc.bus__dat_w[31] ;
 wire \inst$top.soc.bus__dat_w[3] ;
 wire \inst$top.soc.bus__dat_w[4] ;
 wire \inst$top.soc.bus__dat_w[5] ;
 wire \inst$top.soc.bus__dat_w[6] ;
 wire \inst$top.soc.bus__dat_w[7] ;
 wire \inst$top.soc.bus__dat_w[8] ;
 wire \inst$top.soc.bus__dat_w[9] ;
 wire net2543;
 wire \inst$top.soc.cpu.a.source__valid ;
 wire net1885;
 wire \inst$top.soc.cpu.adder$307.x_sub ;
 wire \inst$top.soc.cpu.csr_fmt_i ;
 wire \inst$top.soc.cpu.csrf.bank_300_m_select ;
 wire \inst$top.soc.cpu.csrf.bank_300_w_select ;
 wire \inst$top.soc.cpu.csrf.bank_300_x_select ;
 wire \inst$top.soc.cpu.csrf.d_addr[10] ;
 wire \inst$top.soc.cpu.csrf.d_addr[11] ;
 wire net2295;
 wire net2296;
 wire \inst$top.soc.cpu.csrf.d_addr[4] ;
 wire \inst$top.soc.cpu.csrf.d_addr[5] ;
 wire \inst$top.soc.cpu.csrf.d_addr[6] ;
 wire \inst$top.soc.cpu.csrf.d_addr[7] ;
 wire \inst$top.soc.cpu.csrf.d_addr[8] ;
 wire \inst$top.soc.cpu.csrf.d_addr[9] ;
 wire \inst$top.soc.cpu.d.sink__payload$16.csr_rdy ;
 wire \inst$top.soc.cpu.d.sink__payload$16.csr_we ;
 wire \inst$top.soc.cpu.d.sink__payload$16.load ;
 wire \inst$top.soc.cpu.d.sink__payload$16.multiply ;
 wire \inst$top.soc.cpu.d.sink__payload$16.rd_we ;
 wire \inst$top.soc.cpu.d.sink__payload$6.branch_predict_taken ;
 wire \inst$top.soc.cpu.d.sink__payload$6.branch_taken ;
 wire \inst$top.soc.cpu.d.sink__payload$6.bypass_m ;
 wire \inst$top.soc.cpu.d.sink__payload$6.compare ;
 wire \inst$top.soc.cpu.d.sink__payload$6.condition_met ;
 wire \inst$top.soc.cpu.d.sink__payload$6.csr_we ;
 wire \inst$top.soc.cpu.d.sink__payload$6.divide ;
 wire \inst$top.soc.cpu.d.sink__payload$6.ebreak ;
 wire \inst$top.soc.cpu.d.sink__payload$6.ecall ;
 wire \inst$top.soc.cpu.d.sink__payload$6.illegal ;
 wire \inst$top.soc.cpu.d.sink__payload$6.load ;
 wire \inst$top.soc.cpu.d.sink__payload$6.loadstore_misaligned ;
 wire \inst$top.soc.cpu.d.sink__payload$6.mret ;
 wire \inst$top.soc.cpu.d.sink__payload$6.multiply ;
 wire \inst$top.soc.cpu.d.sink__payload$6.rd_we ;
 wire \inst$top.soc.cpu.d.sink__payload$6.shift ;
 wire \inst$top.soc.cpu.d.sink__payload$6.store ;
 wire \inst$top.soc.cpu.d.sink__payload.auipc ;
 wire \inst$top.soc.cpu.d.sink__payload.branch ;
 wire \inst$top.soc.cpu.d.sink__payload.branch_predict_taken ;
 wire \inst$top.soc.cpu.d.sink__payload.bypass_m ;
 wire \inst$top.soc.cpu.d.sink__payload.bypass_x ;
 wire \inst$top.soc.cpu.d.sink__payload.compare ;
 wire \inst$top.soc.cpu.d.sink__payload.csr_clear ;
 wire \inst$top.soc.cpu.d.sink__payload.csr_fmt_i ;
 wire \inst$top.soc.cpu.d.sink__payload.csr_re ;
 wire \inst$top.soc.cpu.d.sink__payload.csr_set ;
 wire \inst$top.soc.cpu.d.sink__payload.csr_we ;
 wire \inst$top.soc.cpu.d.sink__payload.direction ;
 wire \inst$top.soc.cpu.d.sink__payload.divide ;
 wire \inst$top.soc.cpu.d.sink__payload.ebreak ;
 wire \inst$top.soc.cpu.d.sink__payload.ecall ;
 wire \inst$top.soc.cpu.d.sink__payload.fence_i ;
 wire \inst$top.soc.cpu.d.sink__payload.illegal ;
 wire \inst$top.soc.cpu.d.sink__payload.jump ;
 wire \inst$top.soc.cpu.d.sink__payload.load ;
 wire \inst$top.soc.cpu.d.sink__payload.logic ;
 wire \inst$top.soc.cpu.d.sink__payload.lui ;
 wire \inst$top.soc.cpu.d.sink__payload.mret ;
 wire \inst$top.soc.cpu.d.sink__payload.multiply ;
 wire \inst$top.soc.cpu.d.sink__payload.rd_we ;
 wire \inst$top.soc.cpu.d.sink__payload.rs1_re ;
 wire \inst$top.soc.cpu.d.sink__payload.rs2_re ;
 wire \inst$top.soc.cpu.d.sink__payload.sext ;
 wire \inst$top.soc.cpu.d.sink__payload.shift ;
 wire \inst$top.soc.cpu.d.sink__payload.store ;
 wire \inst$top.soc.cpu.d.source__valid ;
 wire \inst$top.soc.cpu.d_branch_target[2] ;
 wire \inst$top.soc.cpu.d_branch_target[3] ;
 wire \inst$top.soc.cpu.d_offset[12] ;
 wire \inst$top.soc.cpu.d_offset[13] ;
 wire \inst$top.soc.cpu.d_offset[14] ;
 wire \inst$top.soc.cpu.d_offset[15] ;
 wire \inst$top.soc.cpu.d_offset[16] ;
 wire \inst$top.soc.cpu.d_offset[17] ;
 wire \inst$top.soc.cpu.d_offset[18] ;
 wire \inst$top.soc.cpu.d_offset[19] ;
 wire \inst$top.soc.cpu.d_offset[20] ;
 wire \inst$top.soc.cpu.d_offset[21] ;
 wire \inst$top.soc.cpu.d_offset[22] ;
 wire \inst$top.soc.cpu.d_offset[23] ;
 wire \inst$top.soc.cpu.d_offset[24] ;
 wire \inst$top.soc.cpu.d_offset[25] ;
 wire \inst$top.soc.cpu.d_offset[26] ;
 wire \inst$top.soc.cpu.d_offset[27] ;
 wire \inst$top.soc.cpu.d_offset[28] ;
 wire \inst$top.soc.cpu.d_offset[29] ;
 wire \inst$top.soc.cpu.d_offset[30] ;
 wire \inst$top.soc.cpu.divider.divisor[0] ;
 wire \inst$top.soc.cpu.divider.divisor[10] ;
 wire \inst$top.soc.cpu.divider.divisor[11] ;
 wire \inst$top.soc.cpu.divider.divisor[12] ;
 wire \inst$top.soc.cpu.divider.divisor[13] ;
 wire \inst$top.soc.cpu.divider.divisor[14] ;
 wire \inst$top.soc.cpu.divider.divisor[15] ;
 wire \inst$top.soc.cpu.divider.divisor[16] ;
 wire \inst$top.soc.cpu.divider.divisor[17] ;
 wire \inst$top.soc.cpu.divider.divisor[18] ;
 wire \inst$top.soc.cpu.divider.divisor[19] ;
 wire \inst$top.soc.cpu.divider.divisor[1] ;
 wire \inst$top.soc.cpu.divider.divisor[20] ;
 wire \inst$top.soc.cpu.divider.divisor[21] ;
 wire \inst$top.soc.cpu.divider.divisor[22] ;
 wire \inst$top.soc.cpu.divider.divisor[23] ;
 wire \inst$top.soc.cpu.divider.divisor[24] ;
 wire \inst$top.soc.cpu.divider.divisor[25] ;
 wire \inst$top.soc.cpu.divider.divisor[26] ;
 wire \inst$top.soc.cpu.divider.divisor[27] ;
 wire \inst$top.soc.cpu.divider.divisor[28] ;
 wire \inst$top.soc.cpu.divider.divisor[29] ;
 wire \inst$top.soc.cpu.divider.divisor[2] ;
 wire \inst$top.soc.cpu.divider.divisor[30] ;
 wire \inst$top.soc.cpu.divider.divisor[31] ;
 wire \inst$top.soc.cpu.divider.divisor[3] ;
 wire \inst$top.soc.cpu.divider.divisor[4] ;
 wire \inst$top.soc.cpu.divider.divisor[5] ;
 wire \inst$top.soc.cpu.divider.divisor[6] ;
 wire \inst$top.soc.cpu.divider.divisor[7] ;
 wire \inst$top.soc.cpu.divider.divisor[8] ;
 wire \inst$top.soc.cpu.divider.divisor[9] ;
 wire \inst$top.soc.cpu.divider.fsm_state ;
 wire \inst$top.soc.cpu.divider.m_modulus ;
 wire \inst$top.soc.cpu.divider.m_negative ;
 wire \inst$top.soc.cpu.divider.quotient[0] ;
 wire \inst$top.soc.cpu.divider.quotient[10] ;
 wire \inst$top.soc.cpu.divider.quotient[11] ;
 wire \inst$top.soc.cpu.divider.quotient[12] ;
 wire \inst$top.soc.cpu.divider.quotient[13] ;
 wire \inst$top.soc.cpu.divider.quotient[14] ;
 wire \inst$top.soc.cpu.divider.quotient[15] ;
 wire \inst$top.soc.cpu.divider.quotient[16] ;
 wire \inst$top.soc.cpu.divider.quotient[17] ;
 wire \inst$top.soc.cpu.divider.quotient[18] ;
 wire \inst$top.soc.cpu.divider.quotient[19] ;
 wire \inst$top.soc.cpu.divider.quotient[1] ;
 wire \inst$top.soc.cpu.divider.quotient[20] ;
 wire \inst$top.soc.cpu.divider.quotient[21] ;
 wire \inst$top.soc.cpu.divider.quotient[22] ;
 wire \inst$top.soc.cpu.divider.quotient[23] ;
 wire \inst$top.soc.cpu.divider.quotient[24] ;
 wire \inst$top.soc.cpu.divider.quotient[25] ;
 wire \inst$top.soc.cpu.divider.quotient[26] ;
 wire \inst$top.soc.cpu.divider.quotient[27] ;
 wire \inst$top.soc.cpu.divider.quotient[28] ;
 wire \inst$top.soc.cpu.divider.quotient[29] ;
 wire \inst$top.soc.cpu.divider.quotient[2] ;
 wire \inst$top.soc.cpu.divider.quotient[30] ;
 wire \inst$top.soc.cpu.divider.quotient[31] ;
 wire \inst$top.soc.cpu.divider.quotient[3] ;
 wire \inst$top.soc.cpu.divider.quotient[4] ;
 wire \inst$top.soc.cpu.divider.quotient[5] ;
 wire \inst$top.soc.cpu.divider.quotient[6] ;
 wire \inst$top.soc.cpu.divider.quotient[7] ;
 wire \inst$top.soc.cpu.divider.quotient[8] ;
 wire \inst$top.soc.cpu.divider.quotient[9] ;
 wire \inst$top.soc.cpu.divider.remainder[0] ;
 wire \inst$top.soc.cpu.divider.remainder[10] ;
 wire \inst$top.soc.cpu.divider.remainder[11] ;
 wire \inst$top.soc.cpu.divider.remainder[12] ;
 wire \inst$top.soc.cpu.divider.remainder[13] ;
 wire \inst$top.soc.cpu.divider.remainder[14] ;
 wire \inst$top.soc.cpu.divider.remainder[15] ;
 wire \inst$top.soc.cpu.divider.remainder[16] ;
 wire \inst$top.soc.cpu.divider.remainder[17] ;
 wire \inst$top.soc.cpu.divider.remainder[18] ;
 wire \inst$top.soc.cpu.divider.remainder[19] ;
 wire \inst$top.soc.cpu.divider.remainder[1] ;
 wire \inst$top.soc.cpu.divider.remainder[20] ;
 wire \inst$top.soc.cpu.divider.remainder[21] ;
 wire \inst$top.soc.cpu.divider.remainder[22] ;
 wire \inst$top.soc.cpu.divider.remainder[23] ;
 wire \inst$top.soc.cpu.divider.remainder[24] ;
 wire \inst$top.soc.cpu.divider.remainder[25] ;
 wire \inst$top.soc.cpu.divider.remainder[26] ;
 wire \inst$top.soc.cpu.divider.remainder[27] ;
 wire \inst$top.soc.cpu.divider.remainder[28] ;
 wire \inst$top.soc.cpu.divider.remainder[29] ;
 wire \inst$top.soc.cpu.divider.remainder[2] ;
 wire \inst$top.soc.cpu.divider.remainder[30] ;
 wire \inst$top.soc.cpu.divider.remainder[31] ;
 wire \inst$top.soc.cpu.divider.remainder[3] ;
 wire \inst$top.soc.cpu.divider.remainder[4] ;
 wire \inst$top.soc.cpu.divider.remainder[5] ;
 wire \inst$top.soc.cpu.divider.remainder[6] ;
 wire \inst$top.soc.cpu.divider.remainder[7] ;
 wire \inst$top.soc.cpu.divider.remainder[8] ;
 wire \inst$top.soc.cpu.divider.remainder[9] ;
 wire \inst$top.soc.cpu.divider.timer[0] ;
 wire \inst$top.soc.cpu.divider.timer[1] ;
 wire \inst$top.soc.cpu.divider.timer[2] ;
 wire \inst$top.soc.cpu.divider.timer[3] ;
 wire \inst$top.soc.cpu.divider.timer[4] ;
 wire \inst$top.soc.cpu.divider.timer[5] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[10] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[11] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[12] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[13] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[14] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[15] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[16] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[17] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[18] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[19] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[20] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[21] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[22] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[23] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[24] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[25] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[26] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[27] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[28] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[29] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[2] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[30] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[31] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[3] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[4] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[5] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[6] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[7] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[8] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[9] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[10] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[11] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[12] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[13] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[14] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[15] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[16] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[17] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[18] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[19] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[20] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[21] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[22] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[23] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[24] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[25] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[26] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[27] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[28] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[29] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[2] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[30] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[31] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[3] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[4] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[5] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[6] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[7] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[8] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[9] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[10] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[11] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[12] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[13] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[14] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[15] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[16] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[17] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[18] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[19] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[20] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[21] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[22] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[23] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[24] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[25] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[26] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[27] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[28] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[29] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[2] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[30] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[31] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[3] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[4] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[5] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[6] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[7] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[8] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[9] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause_m_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause_w_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mcause_x_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[10] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[11] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[12] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[13] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[14] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[15] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[16] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[17] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[18] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[19] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[20] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[21] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[22] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[23] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[24] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[25] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[26] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[27] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[28] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[29] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[2] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[3] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[4] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[5] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[6] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[7] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[8] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[9] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc_m_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc_w_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mepc_x_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.meie.x_data ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[10] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[11] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[12] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[13] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[14] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[15] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[2] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[3] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[4] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[5] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[6] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[7] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[8] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[9] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.msie.x_data ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie.mtie.x_data ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie_m_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie_w_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mie_x_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.meip.x_data ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[10] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[11] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[12] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[13] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[14] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[15] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[2] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[3] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[4] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[5] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[6] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[7] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[8] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[9] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.msip.x_data ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip.mtip.x_data ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip_m_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip_w_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mip_x_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[10] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[11] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[12] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[13] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[14] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[15] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[16] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[17] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[18] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[19] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[20] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[21] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[22] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[23] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[24] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[25] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[2] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[3] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[4] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[5] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[6] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[7] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[8] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[9] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.mxl.x_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa.mxl.x_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa_m_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa_w_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.misa_x_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[10] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[11] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[12] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[13] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[14] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[15] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[16] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[17] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[18] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[19] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[20] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[21] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[22] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[23] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[24] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[25] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[26] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[27] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[28] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[29] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[2] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[30] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[31] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[3] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[4] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[5] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[6] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[7] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[8] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[9] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch_m_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch_w_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mscratch_x_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mstatus.mie.x_data ;
 wire \inst$top.soc.cpu.exception.csr_bank.mstatus.mpie.w_data ;
 wire \inst$top.soc.cpu.exception.csr_bank.mstatus.mpie.x_data ;
 wire \inst$top.soc.cpu.exception.csr_bank.mstatus.mpp.x_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mstatus.mpp.x_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mstatus_m_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mstatus_w_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mstatus_x_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[10] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[11] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[12] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[13] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[14] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[15] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[16] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[17] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[18] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[19] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[20] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[21] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[22] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[23] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[24] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[25] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[26] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[27] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[28] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[29] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[2] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[30] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[31] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[3] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[4] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[5] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[6] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[7] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[8] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[9] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval_m_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval_w_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtval_x_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[10] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[11] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[12] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[13] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[14] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[15] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[16] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[17] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[18] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[19] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[20] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[21] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[22] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[23] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[24] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[25] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[26] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[27] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[28] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[29] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[2] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[3] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[4] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[5] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[6] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[7] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[8] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[9] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.mode.x_data[0] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec.mode.x_data[1] ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec_m_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec_w_select ;
 wire \inst$top.soc.cpu.exception.csr_bank.mtvec_x_select ;
 wire \inst$top.soc.cpu.exception.m_mie.meie ;
 wire \inst$top.soc.cpu.exception.m_mie.msie ;
 wire \inst$top.soc.cpu.exception.m_mie.mtie ;
 wire \inst$top.soc.cpu.exception.m_mie[10] ;
 wire \inst$top.soc.cpu.exception.m_mie[11] ;
 wire \inst$top.soc.cpu.exception.m_mie[12] ;
 wire \inst$top.soc.cpu.exception.m_mie[13] ;
 wire \inst$top.soc.cpu.exception.m_mie[14] ;
 wire \inst$top.soc.cpu.exception.m_mie[15] ;
 wire \inst$top.soc.cpu.exception.m_mie[16] ;
 wire \inst$top.soc.cpu.exception.m_mie[17] ;
 wire \inst$top.soc.cpu.exception.m_mie[18] ;
 wire \inst$top.soc.cpu.exception.m_mie[3] ;
 wire \inst$top.soc.cpu.exception.m_mie[4] ;
 wire \inst$top.soc.cpu.exception.m_mie[5] ;
 wire \inst$top.soc.cpu.exception.m_mie[6] ;
 wire \inst$top.soc.cpu.exception.m_mie[7] ;
 wire \inst$top.soc.cpu.exception.m_mie[8] ;
 wire \inst$top.soc.cpu.exception.m_mie[9] ;
 wire \inst$top.soc.cpu.exception.m_mip.meip ;
 wire \inst$top.soc.cpu.exception.m_mip.msip ;
 wire \inst$top.soc.cpu.exception.m_mip.mtip ;
 wire \inst$top.soc.cpu.exception.m_mip[10] ;
 wire \inst$top.soc.cpu.exception.m_mip[11] ;
 wire \inst$top.soc.cpu.exception.m_mip[12] ;
 wire \inst$top.soc.cpu.exception.m_mip[13] ;
 wire \inst$top.soc.cpu.exception.m_mip[14] ;
 wire \inst$top.soc.cpu.exception.m_mip[15] ;
 wire \inst$top.soc.cpu.exception.m_mip[16] ;
 wire \inst$top.soc.cpu.exception.m_mip[17] ;
 wire \inst$top.soc.cpu.exception.m_mip[18] ;
 wire \inst$top.soc.cpu.exception.m_mip[3] ;
 wire \inst$top.soc.cpu.exception.m_mip[4] ;
 wire \inst$top.soc.cpu.exception.m_mip[5] ;
 wire \inst$top.soc.cpu.exception.m_mip[6] ;
 wire \inst$top.soc.cpu.exception.m_mip[7] ;
 wire \inst$top.soc.cpu.exception.m_mip[8] ;
 wire \inst$top.soc.cpu.exception.m_mip[9] ;
 wire \inst$top.soc.cpu.exception.m_mstatus.mie ;
 wire \inst$top.soc.cpu.exception.m_mstatus.mpie ;
 wire \inst$top.soc.cpu.exception.w_data$48[0] ;
 wire \inst$top.soc.cpu.exception.w_data$48[1] ;
 wire \inst$top.soc.cpu.exception.w_data$48[2] ;
 wire \inst$top.soc.cpu.exception.w_data$48[31] ;
 wire \inst$top.soc.cpu.exception.w_data$48[3] ;
 wire \inst$top.soc.cpu.exception.w_data$48[4] ;
 wire \inst$top.soc.cpu.exception.w_data$51[0] ;
 wire \inst$top.soc.cpu.exception.w_data$51[10] ;
 wire \inst$top.soc.cpu.exception.w_data$51[11] ;
 wire \inst$top.soc.cpu.exception.w_data$51[12] ;
 wire \inst$top.soc.cpu.exception.w_data$51[13] ;
 wire \inst$top.soc.cpu.exception.w_data$51[14] ;
 wire \inst$top.soc.cpu.exception.w_data$51[15] ;
 wire \inst$top.soc.cpu.exception.w_data$51[16] ;
 wire \inst$top.soc.cpu.exception.w_data$51[17] ;
 wire \inst$top.soc.cpu.exception.w_data$51[18] ;
 wire \inst$top.soc.cpu.exception.w_data$51[19] ;
 wire \inst$top.soc.cpu.exception.w_data$51[1] ;
 wire \inst$top.soc.cpu.exception.w_data$51[20] ;
 wire \inst$top.soc.cpu.exception.w_data$51[21] ;
 wire \inst$top.soc.cpu.exception.w_data$51[22] ;
 wire \inst$top.soc.cpu.exception.w_data$51[23] ;
 wire \inst$top.soc.cpu.exception.w_data$51[24] ;
 wire \inst$top.soc.cpu.exception.w_data$51[25] ;
 wire \inst$top.soc.cpu.exception.w_data$51[26] ;
 wire \inst$top.soc.cpu.exception.w_data$51[27] ;
 wire \inst$top.soc.cpu.exception.w_data$51[28] ;
 wire \inst$top.soc.cpu.exception.w_data$51[29] ;
 wire \inst$top.soc.cpu.exception.w_data$51[2] ;
 wire \inst$top.soc.cpu.exception.w_data$51[30] ;
 wire \inst$top.soc.cpu.exception.w_data$51[31] ;
 wire \inst$top.soc.cpu.exception.w_data$51[3] ;
 wire \inst$top.soc.cpu.exception.w_data$51[4] ;
 wire \inst$top.soc.cpu.exception.w_data$51[5] ;
 wire \inst$top.soc.cpu.exception.w_data$51[6] ;
 wire \inst$top.soc.cpu.exception.w_data$51[7] ;
 wire \inst$top.soc.cpu.exception.w_data$51[8] ;
 wire \inst$top.soc.cpu.exception.w_data$51[9] ;
 wire \inst$top.soc.cpu.exception.w_mret ;
 wire \inst$top.soc.cpu.exception.w_mstatus.mpie ;
 wire \inst$top.soc.cpu.exception.w_trap ;
 wire \inst$top.soc.cpu.f.source__valid ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[0] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[10] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[11] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[12] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[13] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[14] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[15] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[16] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[17] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[18] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[19] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[1] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[20] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[21] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[22] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[23] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[24] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[25] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[26] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[27] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[28] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[29] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[2] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[3] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[4] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[5] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[6] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[7] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[8] ;
 wire \inst$top.soc.cpu.fetch.ibus__adr[9] ;
 wire \inst$top.soc.cpu.fetch.ibus__cyc ;
 wire \inst$top.soc.cpu.fetch.ibus__stb ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[0] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[10] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[11] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[12] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[13] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[14] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[15] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[16] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[17] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[18] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[19] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[1] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[20] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[21] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[22] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[23] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[24] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[25] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[26] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[27] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[28] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[29] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[2] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[30] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[31] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[3] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[4] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[5] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[6] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[7] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[8] ;
 wire \inst$top.soc.cpu.fetch.ibus_rdata[9] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[0] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[10] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[11] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[12] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[13] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[14] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[15] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[16] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[17] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[18] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[19] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[1] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[20] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[21] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[22] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[23] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[24] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[25] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[26] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[27] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[28] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[29] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[2] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[30] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[31] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[3] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[4] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[5] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[6] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[7] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[8] ;
 wire \inst$top.soc.cpu.gprf.bypass1.w_wp_data[9] ;
 wire \inst$top.soc.cpu.gprf.mem[0][0] ;
 wire \inst$top.soc.cpu.gprf.mem[0][10] ;
 wire \inst$top.soc.cpu.gprf.mem[0][11] ;
 wire \inst$top.soc.cpu.gprf.mem[0][12] ;
 wire \inst$top.soc.cpu.gprf.mem[0][13] ;
 wire \inst$top.soc.cpu.gprf.mem[0][14] ;
 wire \inst$top.soc.cpu.gprf.mem[0][15] ;
 wire \inst$top.soc.cpu.gprf.mem[0][16] ;
 wire \inst$top.soc.cpu.gprf.mem[0][17] ;
 wire \inst$top.soc.cpu.gprf.mem[0][18] ;
 wire \inst$top.soc.cpu.gprf.mem[0][19] ;
 wire \inst$top.soc.cpu.gprf.mem[0][1] ;
 wire \inst$top.soc.cpu.gprf.mem[0][20] ;
 wire \inst$top.soc.cpu.gprf.mem[0][21] ;
 wire \inst$top.soc.cpu.gprf.mem[0][22] ;
 wire \inst$top.soc.cpu.gprf.mem[0][23] ;
 wire \inst$top.soc.cpu.gprf.mem[0][24] ;
 wire \inst$top.soc.cpu.gprf.mem[0][25] ;
 wire \inst$top.soc.cpu.gprf.mem[0][26] ;
 wire \inst$top.soc.cpu.gprf.mem[0][27] ;
 wire \inst$top.soc.cpu.gprf.mem[0][28] ;
 wire \inst$top.soc.cpu.gprf.mem[0][29] ;
 wire \inst$top.soc.cpu.gprf.mem[0][2] ;
 wire \inst$top.soc.cpu.gprf.mem[0][30] ;
 wire \inst$top.soc.cpu.gprf.mem[0][31] ;
 wire \inst$top.soc.cpu.gprf.mem[0][3] ;
 wire \inst$top.soc.cpu.gprf.mem[0][4] ;
 wire \inst$top.soc.cpu.gprf.mem[0][5] ;
 wire \inst$top.soc.cpu.gprf.mem[0][6] ;
 wire \inst$top.soc.cpu.gprf.mem[0][7] ;
 wire \inst$top.soc.cpu.gprf.mem[0][8] ;
 wire \inst$top.soc.cpu.gprf.mem[0][9] ;
 wire \inst$top.soc.cpu.gprf.mem[10][0] ;
 wire \inst$top.soc.cpu.gprf.mem[10][10] ;
 wire \inst$top.soc.cpu.gprf.mem[10][11] ;
 wire \inst$top.soc.cpu.gprf.mem[10][12] ;
 wire \inst$top.soc.cpu.gprf.mem[10][13] ;
 wire \inst$top.soc.cpu.gprf.mem[10][14] ;
 wire \inst$top.soc.cpu.gprf.mem[10][15] ;
 wire \inst$top.soc.cpu.gprf.mem[10][16] ;
 wire \inst$top.soc.cpu.gprf.mem[10][17] ;
 wire \inst$top.soc.cpu.gprf.mem[10][18] ;
 wire \inst$top.soc.cpu.gprf.mem[10][19] ;
 wire \inst$top.soc.cpu.gprf.mem[10][1] ;
 wire \inst$top.soc.cpu.gprf.mem[10][20] ;
 wire \inst$top.soc.cpu.gprf.mem[10][21] ;
 wire \inst$top.soc.cpu.gprf.mem[10][22] ;
 wire \inst$top.soc.cpu.gprf.mem[10][23] ;
 wire \inst$top.soc.cpu.gprf.mem[10][24] ;
 wire \inst$top.soc.cpu.gprf.mem[10][25] ;
 wire \inst$top.soc.cpu.gprf.mem[10][26] ;
 wire \inst$top.soc.cpu.gprf.mem[10][27] ;
 wire \inst$top.soc.cpu.gprf.mem[10][28] ;
 wire \inst$top.soc.cpu.gprf.mem[10][29] ;
 wire \inst$top.soc.cpu.gprf.mem[10][2] ;
 wire \inst$top.soc.cpu.gprf.mem[10][30] ;
 wire \inst$top.soc.cpu.gprf.mem[10][31] ;
 wire \inst$top.soc.cpu.gprf.mem[10][3] ;
 wire \inst$top.soc.cpu.gprf.mem[10][4] ;
 wire \inst$top.soc.cpu.gprf.mem[10][5] ;
 wire \inst$top.soc.cpu.gprf.mem[10][6] ;
 wire \inst$top.soc.cpu.gprf.mem[10][7] ;
 wire \inst$top.soc.cpu.gprf.mem[10][8] ;
 wire \inst$top.soc.cpu.gprf.mem[10][9] ;
 wire \inst$top.soc.cpu.gprf.mem[11][0] ;
 wire \inst$top.soc.cpu.gprf.mem[11][10] ;
 wire \inst$top.soc.cpu.gprf.mem[11][11] ;
 wire \inst$top.soc.cpu.gprf.mem[11][12] ;
 wire \inst$top.soc.cpu.gprf.mem[11][13] ;
 wire \inst$top.soc.cpu.gprf.mem[11][14] ;
 wire \inst$top.soc.cpu.gprf.mem[11][15] ;
 wire \inst$top.soc.cpu.gprf.mem[11][16] ;
 wire \inst$top.soc.cpu.gprf.mem[11][17] ;
 wire \inst$top.soc.cpu.gprf.mem[11][18] ;
 wire \inst$top.soc.cpu.gprf.mem[11][19] ;
 wire \inst$top.soc.cpu.gprf.mem[11][1] ;
 wire \inst$top.soc.cpu.gprf.mem[11][20] ;
 wire \inst$top.soc.cpu.gprf.mem[11][21] ;
 wire \inst$top.soc.cpu.gprf.mem[11][22] ;
 wire \inst$top.soc.cpu.gprf.mem[11][23] ;
 wire \inst$top.soc.cpu.gprf.mem[11][24] ;
 wire \inst$top.soc.cpu.gprf.mem[11][25] ;
 wire \inst$top.soc.cpu.gprf.mem[11][26] ;
 wire \inst$top.soc.cpu.gprf.mem[11][27] ;
 wire \inst$top.soc.cpu.gprf.mem[11][28] ;
 wire \inst$top.soc.cpu.gprf.mem[11][29] ;
 wire \inst$top.soc.cpu.gprf.mem[11][2] ;
 wire \inst$top.soc.cpu.gprf.mem[11][30] ;
 wire \inst$top.soc.cpu.gprf.mem[11][31] ;
 wire \inst$top.soc.cpu.gprf.mem[11][3] ;
 wire \inst$top.soc.cpu.gprf.mem[11][4] ;
 wire \inst$top.soc.cpu.gprf.mem[11][5] ;
 wire \inst$top.soc.cpu.gprf.mem[11][6] ;
 wire \inst$top.soc.cpu.gprf.mem[11][7] ;
 wire \inst$top.soc.cpu.gprf.mem[11][8] ;
 wire \inst$top.soc.cpu.gprf.mem[11][9] ;
 wire \inst$top.soc.cpu.gprf.mem[12][0] ;
 wire \inst$top.soc.cpu.gprf.mem[12][10] ;
 wire \inst$top.soc.cpu.gprf.mem[12][11] ;
 wire \inst$top.soc.cpu.gprf.mem[12][12] ;
 wire \inst$top.soc.cpu.gprf.mem[12][13] ;
 wire \inst$top.soc.cpu.gprf.mem[12][14] ;
 wire \inst$top.soc.cpu.gprf.mem[12][15] ;
 wire \inst$top.soc.cpu.gprf.mem[12][16] ;
 wire \inst$top.soc.cpu.gprf.mem[12][17] ;
 wire \inst$top.soc.cpu.gprf.mem[12][18] ;
 wire \inst$top.soc.cpu.gprf.mem[12][19] ;
 wire \inst$top.soc.cpu.gprf.mem[12][1] ;
 wire \inst$top.soc.cpu.gprf.mem[12][20] ;
 wire \inst$top.soc.cpu.gprf.mem[12][21] ;
 wire \inst$top.soc.cpu.gprf.mem[12][22] ;
 wire \inst$top.soc.cpu.gprf.mem[12][23] ;
 wire \inst$top.soc.cpu.gprf.mem[12][24] ;
 wire \inst$top.soc.cpu.gprf.mem[12][25] ;
 wire \inst$top.soc.cpu.gprf.mem[12][26] ;
 wire \inst$top.soc.cpu.gprf.mem[12][27] ;
 wire \inst$top.soc.cpu.gprf.mem[12][28] ;
 wire \inst$top.soc.cpu.gprf.mem[12][29] ;
 wire \inst$top.soc.cpu.gprf.mem[12][2] ;
 wire \inst$top.soc.cpu.gprf.mem[12][30] ;
 wire \inst$top.soc.cpu.gprf.mem[12][31] ;
 wire \inst$top.soc.cpu.gprf.mem[12][3] ;
 wire \inst$top.soc.cpu.gprf.mem[12][4] ;
 wire \inst$top.soc.cpu.gprf.mem[12][5] ;
 wire \inst$top.soc.cpu.gprf.mem[12][6] ;
 wire \inst$top.soc.cpu.gprf.mem[12][7] ;
 wire \inst$top.soc.cpu.gprf.mem[12][8] ;
 wire \inst$top.soc.cpu.gprf.mem[12][9] ;
 wire \inst$top.soc.cpu.gprf.mem[13][0] ;
 wire \inst$top.soc.cpu.gprf.mem[13][10] ;
 wire \inst$top.soc.cpu.gprf.mem[13][11] ;
 wire \inst$top.soc.cpu.gprf.mem[13][12] ;
 wire \inst$top.soc.cpu.gprf.mem[13][13] ;
 wire \inst$top.soc.cpu.gprf.mem[13][14] ;
 wire \inst$top.soc.cpu.gprf.mem[13][15] ;
 wire \inst$top.soc.cpu.gprf.mem[13][16] ;
 wire \inst$top.soc.cpu.gprf.mem[13][17] ;
 wire \inst$top.soc.cpu.gprf.mem[13][18] ;
 wire \inst$top.soc.cpu.gprf.mem[13][19] ;
 wire \inst$top.soc.cpu.gprf.mem[13][1] ;
 wire \inst$top.soc.cpu.gprf.mem[13][20] ;
 wire \inst$top.soc.cpu.gprf.mem[13][21] ;
 wire \inst$top.soc.cpu.gprf.mem[13][22] ;
 wire \inst$top.soc.cpu.gprf.mem[13][23] ;
 wire \inst$top.soc.cpu.gprf.mem[13][24] ;
 wire \inst$top.soc.cpu.gprf.mem[13][25] ;
 wire \inst$top.soc.cpu.gprf.mem[13][26] ;
 wire \inst$top.soc.cpu.gprf.mem[13][27] ;
 wire \inst$top.soc.cpu.gprf.mem[13][28] ;
 wire \inst$top.soc.cpu.gprf.mem[13][29] ;
 wire \inst$top.soc.cpu.gprf.mem[13][2] ;
 wire \inst$top.soc.cpu.gprf.mem[13][30] ;
 wire \inst$top.soc.cpu.gprf.mem[13][31] ;
 wire \inst$top.soc.cpu.gprf.mem[13][3] ;
 wire \inst$top.soc.cpu.gprf.mem[13][4] ;
 wire \inst$top.soc.cpu.gprf.mem[13][5] ;
 wire \inst$top.soc.cpu.gprf.mem[13][6] ;
 wire \inst$top.soc.cpu.gprf.mem[13][7] ;
 wire \inst$top.soc.cpu.gprf.mem[13][8] ;
 wire \inst$top.soc.cpu.gprf.mem[13][9] ;
 wire \inst$top.soc.cpu.gprf.mem[14][0] ;
 wire \inst$top.soc.cpu.gprf.mem[14][10] ;
 wire \inst$top.soc.cpu.gprf.mem[14][11] ;
 wire \inst$top.soc.cpu.gprf.mem[14][12] ;
 wire \inst$top.soc.cpu.gprf.mem[14][13] ;
 wire \inst$top.soc.cpu.gprf.mem[14][14] ;
 wire \inst$top.soc.cpu.gprf.mem[14][15] ;
 wire \inst$top.soc.cpu.gprf.mem[14][16] ;
 wire \inst$top.soc.cpu.gprf.mem[14][17] ;
 wire \inst$top.soc.cpu.gprf.mem[14][18] ;
 wire \inst$top.soc.cpu.gprf.mem[14][19] ;
 wire \inst$top.soc.cpu.gprf.mem[14][1] ;
 wire \inst$top.soc.cpu.gprf.mem[14][20] ;
 wire \inst$top.soc.cpu.gprf.mem[14][21] ;
 wire \inst$top.soc.cpu.gprf.mem[14][22] ;
 wire \inst$top.soc.cpu.gprf.mem[14][23] ;
 wire \inst$top.soc.cpu.gprf.mem[14][24] ;
 wire \inst$top.soc.cpu.gprf.mem[14][25] ;
 wire \inst$top.soc.cpu.gprf.mem[14][26] ;
 wire \inst$top.soc.cpu.gprf.mem[14][27] ;
 wire \inst$top.soc.cpu.gprf.mem[14][28] ;
 wire \inst$top.soc.cpu.gprf.mem[14][29] ;
 wire \inst$top.soc.cpu.gprf.mem[14][2] ;
 wire \inst$top.soc.cpu.gprf.mem[14][30] ;
 wire \inst$top.soc.cpu.gprf.mem[14][31] ;
 wire \inst$top.soc.cpu.gprf.mem[14][3] ;
 wire \inst$top.soc.cpu.gprf.mem[14][4] ;
 wire \inst$top.soc.cpu.gprf.mem[14][5] ;
 wire \inst$top.soc.cpu.gprf.mem[14][6] ;
 wire \inst$top.soc.cpu.gprf.mem[14][7] ;
 wire \inst$top.soc.cpu.gprf.mem[14][8] ;
 wire \inst$top.soc.cpu.gprf.mem[14][9] ;
 wire \inst$top.soc.cpu.gprf.mem[15][0] ;
 wire \inst$top.soc.cpu.gprf.mem[15][10] ;
 wire \inst$top.soc.cpu.gprf.mem[15][11] ;
 wire \inst$top.soc.cpu.gprf.mem[15][12] ;
 wire \inst$top.soc.cpu.gprf.mem[15][13] ;
 wire \inst$top.soc.cpu.gprf.mem[15][14] ;
 wire \inst$top.soc.cpu.gprf.mem[15][15] ;
 wire \inst$top.soc.cpu.gprf.mem[15][16] ;
 wire \inst$top.soc.cpu.gprf.mem[15][17] ;
 wire \inst$top.soc.cpu.gprf.mem[15][18] ;
 wire \inst$top.soc.cpu.gprf.mem[15][19] ;
 wire \inst$top.soc.cpu.gprf.mem[15][1] ;
 wire \inst$top.soc.cpu.gprf.mem[15][20] ;
 wire \inst$top.soc.cpu.gprf.mem[15][21] ;
 wire \inst$top.soc.cpu.gprf.mem[15][22] ;
 wire \inst$top.soc.cpu.gprf.mem[15][23] ;
 wire \inst$top.soc.cpu.gprf.mem[15][24] ;
 wire \inst$top.soc.cpu.gprf.mem[15][25] ;
 wire \inst$top.soc.cpu.gprf.mem[15][26] ;
 wire \inst$top.soc.cpu.gprf.mem[15][27] ;
 wire \inst$top.soc.cpu.gprf.mem[15][28] ;
 wire \inst$top.soc.cpu.gprf.mem[15][29] ;
 wire \inst$top.soc.cpu.gprf.mem[15][2] ;
 wire \inst$top.soc.cpu.gprf.mem[15][30] ;
 wire \inst$top.soc.cpu.gprf.mem[15][31] ;
 wire \inst$top.soc.cpu.gprf.mem[15][3] ;
 wire \inst$top.soc.cpu.gprf.mem[15][4] ;
 wire \inst$top.soc.cpu.gprf.mem[15][5] ;
 wire \inst$top.soc.cpu.gprf.mem[15][6] ;
 wire \inst$top.soc.cpu.gprf.mem[15][7] ;
 wire \inst$top.soc.cpu.gprf.mem[15][8] ;
 wire \inst$top.soc.cpu.gprf.mem[15][9] ;
 wire \inst$top.soc.cpu.gprf.mem[16][0] ;
 wire \inst$top.soc.cpu.gprf.mem[16][10] ;
 wire \inst$top.soc.cpu.gprf.mem[16][11] ;
 wire \inst$top.soc.cpu.gprf.mem[16][12] ;
 wire \inst$top.soc.cpu.gprf.mem[16][13] ;
 wire \inst$top.soc.cpu.gprf.mem[16][14] ;
 wire \inst$top.soc.cpu.gprf.mem[16][15] ;
 wire \inst$top.soc.cpu.gprf.mem[16][16] ;
 wire \inst$top.soc.cpu.gprf.mem[16][17] ;
 wire \inst$top.soc.cpu.gprf.mem[16][18] ;
 wire \inst$top.soc.cpu.gprf.mem[16][19] ;
 wire \inst$top.soc.cpu.gprf.mem[16][1] ;
 wire \inst$top.soc.cpu.gprf.mem[16][20] ;
 wire \inst$top.soc.cpu.gprf.mem[16][21] ;
 wire \inst$top.soc.cpu.gprf.mem[16][22] ;
 wire \inst$top.soc.cpu.gprf.mem[16][23] ;
 wire \inst$top.soc.cpu.gprf.mem[16][24] ;
 wire \inst$top.soc.cpu.gprf.mem[16][25] ;
 wire \inst$top.soc.cpu.gprf.mem[16][26] ;
 wire \inst$top.soc.cpu.gprf.mem[16][27] ;
 wire \inst$top.soc.cpu.gprf.mem[16][28] ;
 wire \inst$top.soc.cpu.gprf.mem[16][29] ;
 wire \inst$top.soc.cpu.gprf.mem[16][2] ;
 wire \inst$top.soc.cpu.gprf.mem[16][30] ;
 wire \inst$top.soc.cpu.gprf.mem[16][31] ;
 wire \inst$top.soc.cpu.gprf.mem[16][3] ;
 wire \inst$top.soc.cpu.gprf.mem[16][4] ;
 wire \inst$top.soc.cpu.gprf.mem[16][5] ;
 wire \inst$top.soc.cpu.gprf.mem[16][6] ;
 wire \inst$top.soc.cpu.gprf.mem[16][7] ;
 wire \inst$top.soc.cpu.gprf.mem[16][8] ;
 wire \inst$top.soc.cpu.gprf.mem[16][9] ;
 wire \inst$top.soc.cpu.gprf.mem[17][0] ;
 wire \inst$top.soc.cpu.gprf.mem[17][10] ;
 wire \inst$top.soc.cpu.gprf.mem[17][11] ;
 wire \inst$top.soc.cpu.gprf.mem[17][12] ;
 wire \inst$top.soc.cpu.gprf.mem[17][13] ;
 wire \inst$top.soc.cpu.gprf.mem[17][14] ;
 wire \inst$top.soc.cpu.gprf.mem[17][15] ;
 wire \inst$top.soc.cpu.gprf.mem[17][16] ;
 wire \inst$top.soc.cpu.gprf.mem[17][17] ;
 wire \inst$top.soc.cpu.gprf.mem[17][18] ;
 wire \inst$top.soc.cpu.gprf.mem[17][19] ;
 wire \inst$top.soc.cpu.gprf.mem[17][1] ;
 wire \inst$top.soc.cpu.gprf.mem[17][20] ;
 wire \inst$top.soc.cpu.gprf.mem[17][21] ;
 wire \inst$top.soc.cpu.gprf.mem[17][22] ;
 wire \inst$top.soc.cpu.gprf.mem[17][23] ;
 wire \inst$top.soc.cpu.gprf.mem[17][24] ;
 wire \inst$top.soc.cpu.gprf.mem[17][25] ;
 wire \inst$top.soc.cpu.gprf.mem[17][26] ;
 wire \inst$top.soc.cpu.gprf.mem[17][27] ;
 wire \inst$top.soc.cpu.gprf.mem[17][28] ;
 wire \inst$top.soc.cpu.gprf.mem[17][29] ;
 wire \inst$top.soc.cpu.gprf.mem[17][2] ;
 wire \inst$top.soc.cpu.gprf.mem[17][30] ;
 wire \inst$top.soc.cpu.gprf.mem[17][31] ;
 wire \inst$top.soc.cpu.gprf.mem[17][3] ;
 wire \inst$top.soc.cpu.gprf.mem[17][4] ;
 wire \inst$top.soc.cpu.gprf.mem[17][5] ;
 wire \inst$top.soc.cpu.gprf.mem[17][6] ;
 wire \inst$top.soc.cpu.gprf.mem[17][7] ;
 wire \inst$top.soc.cpu.gprf.mem[17][8] ;
 wire \inst$top.soc.cpu.gprf.mem[17][9] ;
 wire \inst$top.soc.cpu.gprf.mem[18][0] ;
 wire \inst$top.soc.cpu.gprf.mem[18][10] ;
 wire \inst$top.soc.cpu.gprf.mem[18][11] ;
 wire \inst$top.soc.cpu.gprf.mem[18][12] ;
 wire \inst$top.soc.cpu.gprf.mem[18][13] ;
 wire \inst$top.soc.cpu.gprf.mem[18][14] ;
 wire \inst$top.soc.cpu.gprf.mem[18][15] ;
 wire \inst$top.soc.cpu.gprf.mem[18][16] ;
 wire \inst$top.soc.cpu.gprf.mem[18][17] ;
 wire \inst$top.soc.cpu.gprf.mem[18][18] ;
 wire \inst$top.soc.cpu.gprf.mem[18][19] ;
 wire \inst$top.soc.cpu.gprf.mem[18][1] ;
 wire \inst$top.soc.cpu.gprf.mem[18][20] ;
 wire \inst$top.soc.cpu.gprf.mem[18][21] ;
 wire \inst$top.soc.cpu.gprf.mem[18][22] ;
 wire \inst$top.soc.cpu.gprf.mem[18][23] ;
 wire \inst$top.soc.cpu.gprf.mem[18][24] ;
 wire \inst$top.soc.cpu.gprf.mem[18][25] ;
 wire \inst$top.soc.cpu.gprf.mem[18][26] ;
 wire \inst$top.soc.cpu.gprf.mem[18][27] ;
 wire \inst$top.soc.cpu.gprf.mem[18][28] ;
 wire \inst$top.soc.cpu.gprf.mem[18][29] ;
 wire \inst$top.soc.cpu.gprf.mem[18][2] ;
 wire \inst$top.soc.cpu.gprf.mem[18][30] ;
 wire \inst$top.soc.cpu.gprf.mem[18][31] ;
 wire \inst$top.soc.cpu.gprf.mem[18][3] ;
 wire \inst$top.soc.cpu.gprf.mem[18][4] ;
 wire \inst$top.soc.cpu.gprf.mem[18][5] ;
 wire \inst$top.soc.cpu.gprf.mem[18][6] ;
 wire \inst$top.soc.cpu.gprf.mem[18][7] ;
 wire \inst$top.soc.cpu.gprf.mem[18][8] ;
 wire \inst$top.soc.cpu.gprf.mem[18][9] ;
 wire \inst$top.soc.cpu.gprf.mem[19][0] ;
 wire \inst$top.soc.cpu.gprf.mem[19][10] ;
 wire \inst$top.soc.cpu.gprf.mem[19][11] ;
 wire \inst$top.soc.cpu.gprf.mem[19][12] ;
 wire \inst$top.soc.cpu.gprf.mem[19][13] ;
 wire \inst$top.soc.cpu.gprf.mem[19][14] ;
 wire \inst$top.soc.cpu.gprf.mem[19][15] ;
 wire \inst$top.soc.cpu.gprf.mem[19][16] ;
 wire \inst$top.soc.cpu.gprf.mem[19][17] ;
 wire \inst$top.soc.cpu.gprf.mem[19][18] ;
 wire \inst$top.soc.cpu.gprf.mem[19][19] ;
 wire \inst$top.soc.cpu.gprf.mem[19][1] ;
 wire \inst$top.soc.cpu.gprf.mem[19][20] ;
 wire \inst$top.soc.cpu.gprf.mem[19][21] ;
 wire \inst$top.soc.cpu.gprf.mem[19][22] ;
 wire \inst$top.soc.cpu.gprf.mem[19][23] ;
 wire \inst$top.soc.cpu.gprf.mem[19][24] ;
 wire \inst$top.soc.cpu.gprf.mem[19][25] ;
 wire \inst$top.soc.cpu.gprf.mem[19][26] ;
 wire \inst$top.soc.cpu.gprf.mem[19][27] ;
 wire \inst$top.soc.cpu.gprf.mem[19][28] ;
 wire \inst$top.soc.cpu.gprf.mem[19][29] ;
 wire \inst$top.soc.cpu.gprf.mem[19][2] ;
 wire \inst$top.soc.cpu.gprf.mem[19][30] ;
 wire \inst$top.soc.cpu.gprf.mem[19][31] ;
 wire \inst$top.soc.cpu.gprf.mem[19][3] ;
 wire \inst$top.soc.cpu.gprf.mem[19][4] ;
 wire \inst$top.soc.cpu.gprf.mem[19][5] ;
 wire \inst$top.soc.cpu.gprf.mem[19][6] ;
 wire \inst$top.soc.cpu.gprf.mem[19][7] ;
 wire \inst$top.soc.cpu.gprf.mem[19][8] ;
 wire \inst$top.soc.cpu.gprf.mem[19][9] ;
 wire \inst$top.soc.cpu.gprf.mem[1][0] ;
 wire \inst$top.soc.cpu.gprf.mem[1][10] ;
 wire \inst$top.soc.cpu.gprf.mem[1][11] ;
 wire \inst$top.soc.cpu.gprf.mem[1][12] ;
 wire \inst$top.soc.cpu.gprf.mem[1][13] ;
 wire \inst$top.soc.cpu.gprf.mem[1][14] ;
 wire \inst$top.soc.cpu.gprf.mem[1][15] ;
 wire \inst$top.soc.cpu.gprf.mem[1][16] ;
 wire \inst$top.soc.cpu.gprf.mem[1][17] ;
 wire \inst$top.soc.cpu.gprf.mem[1][18] ;
 wire \inst$top.soc.cpu.gprf.mem[1][19] ;
 wire \inst$top.soc.cpu.gprf.mem[1][1] ;
 wire \inst$top.soc.cpu.gprf.mem[1][20] ;
 wire \inst$top.soc.cpu.gprf.mem[1][21] ;
 wire \inst$top.soc.cpu.gprf.mem[1][22] ;
 wire \inst$top.soc.cpu.gprf.mem[1][23] ;
 wire \inst$top.soc.cpu.gprf.mem[1][24] ;
 wire \inst$top.soc.cpu.gprf.mem[1][25] ;
 wire \inst$top.soc.cpu.gprf.mem[1][26] ;
 wire \inst$top.soc.cpu.gprf.mem[1][27] ;
 wire \inst$top.soc.cpu.gprf.mem[1][28] ;
 wire \inst$top.soc.cpu.gprf.mem[1][29] ;
 wire \inst$top.soc.cpu.gprf.mem[1][2] ;
 wire \inst$top.soc.cpu.gprf.mem[1][30] ;
 wire \inst$top.soc.cpu.gprf.mem[1][31] ;
 wire \inst$top.soc.cpu.gprf.mem[1][3] ;
 wire \inst$top.soc.cpu.gprf.mem[1][4] ;
 wire \inst$top.soc.cpu.gprf.mem[1][5] ;
 wire \inst$top.soc.cpu.gprf.mem[1][6] ;
 wire \inst$top.soc.cpu.gprf.mem[1][7] ;
 wire \inst$top.soc.cpu.gprf.mem[1][8] ;
 wire \inst$top.soc.cpu.gprf.mem[1][9] ;
 wire \inst$top.soc.cpu.gprf.mem[20][0] ;
 wire \inst$top.soc.cpu.gprf.mem[20][10] ;
 wire \inst$top.soc.cpu.gprf.mem[20][11] ;
 wire \inst$top.soc.cpu.gprf.mem[20][12] ;
 wire \inst$top.soc.cpu.gprf.mem[20][13] ;
 wire \inst$top.soc.cpu.gprf.mem[20][14] ;
 wire \inst$top.soc.cpu.gprf.mem[20][15] ;
 wire \inst$top.soc.cpu.gprf.mem[20][16] ;
 wire \inst$top.soc.cpu.gprf.mem[20][17] ;
 wire \inst$top.soc.cpu.gprf.mem[20][18] ;
 wire \inst$top.soc.cpu.gprf.mem[20][19] ;
 wire \inst$top.soc.cpu.gprf.mem[20][1] ;
 wire \inst$top.soc.cpu.gprf.mem[20][20] ;
 wire \inst$top.soc.cpu.gprf.mem[20][21] ;
 wire \inst$top.soc.cpu.gprf.mem[20][22] ;
 wire \inst$top.soc.cpu.gprf.mem[20][23] ;
 wire \inst$top.soc.cpu.gprf.mem[20][24] ;
 wire \inst$top.soc.cpu.gprf.mem[20][25] ;
 wire \inst$top.soc.cpu.gprf.mem[20][26] ;
 wire \inst$top.soc.cpu.gprf.mem[20][27] ;
 wire \inst$top.soc.cpu.gprf.mem[20][28] ;
 wire \inst$top.soc.cpu.gprf.mem[20][29] ;
 wire \inst$top.soc.cpu.gprf.mem[20][2] ;
 wire \inst$top.soc.cpu.gprf.mem[20][30] ;
 wire \inst$top.soc.cpu.gprf.mem[20][31] ;
 wire \inst$top.soc.cpu.gprf.mem[20][3] ;
 wire \inst$top.soc.cpu.gprf.mem[20][4] ;
 wire \inst$top.soc.cpu.gprf.mem[20][5] ;
 wire \inst$top.soc.cpu.gprf.mem[20][6] ;
 wire \inst$top.soc.cpu.gprf.mem[20][7] ;
 wire \inst$top.soc.cpu.gprf.mem[20][8] ;
 wire \inst$top.soc.cpu.gprf.mem[20][9] ;
 wire \inst$top.soc.cpu.gprf.mem[21][0] ;
 wire \inst$top.soc.cpu.gprf.mem[21][10] ;
 wire \inst$top.soc.cpu.gprf.mem[21][11] ;
 wire \inst$top.soc.cpu.gprf.mem[21][12] ;
 wire \inst$top.soc.cpu.gprf.mem[21][13] ;
 wire \inst$top.soc.cpu.gprf.mem[21][14] ;
 wire \inst$top.soc.cpu.gprf.mem[21][15] ;
 wire \inst$top.soc.cpu.gprf.mem[21][16] ;
 wire \inst$top.soc.cpu.gprf.mem[21][17] ;
 wire \inst$top.soc.cpu.gprf.mem[21][18] ;
 wire \inst$top.soc.cpu.gprf.mem[21][19] ;
 wire \inst$top.soc.cpu.gprf.mem[21][1] ;
 wire \inst$top.soc.cpu.gprf.mem[21][20] ;
 wire \inst$top.soc.cpu.gprf.mem[21][21] ;
 wire \inst$top.soc.cpu.gprf.mem[21][22] ;
 wire \inst$top.soc.cpu.gprf.mem[21][23] ;
 wire \inst$top.soc.cpu.gprf.mem[21][24] ;
 wire \inst$top.soc.cpu.gprf.mem[21][25] ;
 wire \inst$top.soc.cpu.gprf.mem[21][26] ;
 wire \inst$top.soc.cpu.gprf.mem[21][27] ;
 wire \inst$top.soc.cpu.gprf.mem[21][28] ;
 wire \inst$top.soc.cpu.gprf.mem[21][29] ;
 wire \inst$top.soc.cpu.gprf.mem[21][2] ;
 wire \inst$top.soc.cpu.gprf.mem[21][30] ;
 wire \inst$top.soc.cpu.gprf.mem[21][31] ;
 wire \inst$top.soc.cpu.gprf.mem[21][3] ;
 wire \inst$top.soc.cpu.gprf.mem[21][4] ;
 wire \inst$top.soc.cpu.gprf.mem[21][5] ;
 wire \inst$top.soc.cpu.gprf.mem[21][6] ;
 wire \inst$top.soc.cpu.gprf.mem[21][7] ;
 wire \inst$top.soc.cpu.gprf.mem[21][8] ;
 wire \inst$top.soc.cpu.gprf.mem[21][9] ;
 wire \inst$top.soc.cpu.gprf.mem[22][0] ;
 wire \inst$top.soc.cpu.gprf.mem[22][10] ;
 wire \inst$top.soc.cpu.gprf.mem[22][11] ;
 wire \inst$top.soc.cpu.gprf.mem[22][12] ;
 wire \inst$top.soc.cpu.gprf.mem[22][13] ;
 wire \inst$top.soc.cpu.gprf.mem[22][14] ;
 wire \inst$top.soc.cpu.gprf.mem[22][15] ;
 wire \inst$top.soc.cpu.gprf.mem[22][16] ;
 wire \inst$top.soc.cpu.gprf.mem[22][17] ;
 wire \inst$top.soc.cpu.gprf.mem[22][18] ;
 wire \inst$top.soc.cpu.gprf.mem[22][19] ;
 wire \inst$top.soc.cpu.gprf.mem[22][1] ;
 wire \inst$top.soc.cpu.gprf.mem[22][20] ;
 wire \inst$top.soc.cpu.gprf.mem[22][21] ;
 wire \inst$top.soc.cpu.gprf.mem[22][22] ;
 wire \inst$top.soc.cpu.gprf.mem[22][23] ;
 wire \inst$top.soc.cpu.gprf.mem[22][24] ;
 wire \inst$top.soc.cpu.gprf.mem[22][25] ;
 wire \inst$top.soc.cpu.gprf.mem[22][26] ;
 wire \inst$top.soc.cpu.gprf.mem[22][27] ;
 wire \inst$top.soc.cpu.gprf.mem[22][28] ;
 wire \inst$top.soc.cpu.gprf.mem[22][29] ;
 wire \inst$top.soc.cpu.gprf.mem[22][2] ;
 wire \inst$top.soc.cpu.gprf.mem[22][30] ;
 wire \inst$top.soc.cpu.gprf.mem[22][31] ;
 wire \inst$top.soc.cpu.gprf.mem[22][3] ;
 wire \inst$top.soc.cpu.gprf.mem[22][4] ;
 wire \inst$top.soc.cpu.gprf.mem[22][5] ;
 wire \inst$top.soc.cpu.gprf.mem[22][6] ;
 wire \inst$top.soc.cpu.gprf.mem[22][7] ;
 wire \inst$top.soc.cpu.gprf.mem[22][8] ;
 wire \inst$top.soc.cpu.gprf.mem[22][9] ;
 wire \inst$top.soc.cpu.gprf.mem[23][0] ;
 wire \inst$top.soc.cpu.gprf.mem[23][10] ;
 wire \inst$top.soc.cpu.gprf.mem[23][11] ;
 wire \inst$top.soc.cpu.gprf.mem[23][12] ;
 wire \inst$top.soc.cpu.gprf.mem[23][13] ;
 wire \inst$top.soc.cpu.gprf.mem[23][14] ;
 wire \inst$top.soc.cpu.gprf.mem[23][15] ;
 wire \inst$top.soc.cpu.gprf.mem[23][16] ;
 wire \inst$top.soc.cpu.gprf.mem[23][17] ;
 wire \inst$top.soc.cpu.gprf.mem[23][18] ;
 wire \inst$top.soc.cpu.gprf.mem[23][19] ;
 wire \inst$top.soc.cpu.gprf.mem[23][1] ;
 wire \inst$top.soc.cpu.gprf.mem[23][20] ;
 wire \inst$top.soc.cpu.gprf.mem[23][21] ;
 wire \inst$top.soc.cpu.gprf.mem[23][22] ;
 wire \inst$top.soc.cpu.gprf.mem[23][23] ;
 wire \inst$top.soc.cpu.gprf.mem[23][24] ;
 wire \inst$top.soc.cpu.gprf.mem[23][25] ;
 wire \inst$top.soc.cpu.gprf.mem[23][26] ;
 wire \inst$top.soc.cpu.gprf.mem[23][27] ;
 wire \inst$top.soc.cpu.gprf.mem[23][28] ;
 wire \inst$top.soc.cpu.gprf.mem[23][29] ;
 wire \inst$top.soc.cpu.gprf.mem[23][2] ;
 wire \inst$top.soc.cpu.gprf.mem[23][30] ;
 wire \inst$top.soc.cpu.gprf.mem[23][31] ;
 wire \inst$top.soc.cpu.gprf.mem[23][3] ;
 wire \inst$top.soc.cpu.gprf.mem[23][4] ;
 wire \inst$top.soc.cpu.gprf.mem[23][5] ;
 wire \inst$top.soc.cpu.gprf.mem[23][6] ;
 wire \inst$top.soc.cpu.gprf.mem[23][7] ;
 wire \inst$top.soc.cpu.gprf.mem[23][8] ;
 wire \inst$top.soc.cpu.gprf.mem[23][9] ;
 wire \inst$top.soc.cpu.gprf.mem[24][0] ;
 wire \inst$top.soc.cpu.gprf.mem[24][10] ;
 wire \inst$top.soc.cpu.gprf.mem[24][11] ;
 wire \inst$top.soc.cpu.gprf.mem[24][12] ;
 wire \inst$top.soc.cpu.gprf.mem[24][13] ;
 wire \inst$top.soc.cpu.gprf.mem[24][14] ;
 wire \inst$top.soc.cpu.gprf.mem[24][15] ;
 wire \inst$top.soc.cpu.gprf.mem[24][16] ;
 wire \inst$top.soc.cpu.gprf.mem[24][17] ;
 wire \inst$top.soc.cpu.gprf.mem[24][18] ;
 wire \inst$top.soc.cpu.gprf.mem[24][19] ;
 wire \inst$top.soc.cpu.gprf.mem[24][1] ;
 wire \inst$top.soc.cpu.gprf.mem[24][20] ;
 wire \inst$top.soc.cpu.gprf.mem[24][21] ;
 wire \inst$top.soc.cpu.gprf.mem[24][22] ;
 wire \inst$top.soc.cpu.gprf.mem[24][23] ;
 wire \inst$top.soc.cpu.gprf.mem[24][24] ;
 wire \inst$top.soc.cpu.gprf.mem[24][25] ;
 wire \inst$top.soc.cpu.gprf.mem[24][26] ;
 wire \inst$top.soc.cpu.gprf.mem[24][27] ;
 wire \inst$top.soc.cpu.gprf.mem[24][28] ;
 wire \inst$top.soc.cpu.gprf.mem[24][29] ;
 wire \inst$top.soc.cpu.gprf.mem[24][2] ;
 wire \inst$top.soc.cpu.gprf.mem[24][30] ;
 wire \inst$top.soc.cpu.gprf.mem[24][31] ;
 wire \inst$top.soc.cpu.gprf.mem[24][3] ;
 wire \inst$top.soc.cpu.gprf.mem[24][4] ;
 wire \inst$top.soc.cpu.gprf.mem[24][5] ;
 wire \inst$top.soc.cpu.gprf.mem[24][6] ;
 wire \inst$top.soc.cpu.gprf.mem[24][7] ;
 wire \inst$top.soc.cpu.gprf.mem[24][8] ;
 wire \inst$top.soc.cpu.gprf.mem[24][9] ;
 wire \inst$top.soc.cpu.gprf.mem[25][0] ;
 wire \inst$top.soc.cpu.gprf.mem[25][10] ;
 wire \inst$top.soc.cpu.gprf.mem[25][11] ;
 wire \inst$top.soc.cpu.gprf.mem[25][12] ;
 wire \inst$top.soc.cpu.gprf.mem[25][13] ;
 wire \inst$top.soc.cpu.gprf.mem[25][14] ;
 wire \inst$top.soc.cpu.gprf.mem[25][15] ;
 wire \inst$top.soc.cpu.gprf.mem[25][16] ;
 wire \inst$top.soc.cpu.gprf.mem[25][17] ;
 wire \inst$top.soc.cpu.gprf.mem[25][18] ;
 wire \inst$top.soc.cpu.gprf.mem[25][19] ;
 wire \inst$top.soc.cpu.gprf.mem[25][1] ;
 wire \inst$top.soc.cpu.gprf.mem[25][20] ;
 wire \inst$top.soc.cpu.gprf.mem[25][21] ;
 wire \inst$top.soc.cpu.gprf.mem[25][22] ;
 wire \inst$top.soc.cpu.gprf.mem[25][23] ;
 wire \inst$top.soc.cpu.gprf.mem[25][24] ;
 wire \inst$top.soc.cpu.gprf.mem[25][25] ;
 wire \inst$top.soc.cpu.gprf.mem[25][26] ;
 wire \inst$top.soc.cpu.gprf.mem[25][27] ;
 wire \inst$top.soc.cpu.gprf.mem[25][28] ;
 wire \inst$top.soc.cpu.gprf.mem[25][29] ;
 wire \inst$top.soc.cpu.gprf.mem[25][2] ;
 wire \inst$top.soc.cpu.gprf.mem[25][30] ;
 wire \inst$top.soc.cpu.gprf.mem[25][31] ;
 wire \inst$top.soc.cpu.gprf.mem[25][3] ;
 wire \inst$top.soc.cpu.gprf.mem[25][4] ;
 wire \inst$top.soc.cpu.gprf.mem[25][5] ;
 wire \inst$top.soc.cpu.gprf.mem[25][6] ;
 wire \inst$top.soc.cpu.gprf.mem[25][7] ;
 wire \inst$top.soc.cpu.gprf.mem[25][8] ;
 wire \inst$top.soc.cpu.gprf.mem[25][9] ;
 wire \inst$top.soc.cpu.gprf.mem[26][0] ;
 wire \inst$top.soc.cpu.gprf.mem[26][10] ;
 wire \inst$top.soc.cpu.gprf.mem[26][11] ;
 wire \inst$top.soc.cpu.gprf.mem[26][12] ;
 wire \inst$top.soc.cpu.gprf.mem[26][13] ;
 wire \inst$top.soc.cpu.gprf.mem[26][14] ;
 wire \inst$top.soc.cpu.gprf.mem[26][15] ;
 wire \inst$top.soc.cpu.gprf.mem[26][16] ;
 wire \inst$top.soc.cpu.gprf.mem[26][17] ;
 wire \inst$top.soc.cpu.gprf.mem[26][18] ;
 wire \inst$top.soc.cpu.gprf.mem[26][19] ;
 wire \inst$top.soc.cpu.gprf.mem[26][1] ;
 wire \inst$top.soc.cpu.gprf.mem[26][20] ;
 wire \inst$top.soc.cpu.gprf.mem[26][21] ;
 wire \inst$top.soc.cpu.gprf.mem[26][22] ;
 wire \inst$top.soc.cpu.gprf.mem[26][23] ;
 wire \inst$top.soc.cpu.gprf.mem[26][24] ;
 wire \inst$top.soc.cpu.gprf.mem[26][25] ;
 wire \inst$top.soc.cpu.gprf.mem[26][26] ;
 wire \inst$top.soc.cpu.gprf.mem[26][27] ;
 wire \inst$top.soc.cpu.gprf.mem[26][28] ;
 wire \inst$top.soc.cpu.gprf.mem[26][29] ;
 wire \inst$top.soc.cpu.gprf.mem[26][2] ;
 wire \inst$top.soc.cpu.gprf.mem[26][30] ;
 wire \inst$top.soc.cpu.gprf.mem[26][31] ;
 wire \inst$top.soc.cpu.gprf.mem[26][3] ;
 wire \inst$top.soc.cpu.gprf.mem[26][4] ;
 wire \inst$top.soc.cpu.gprf.mem[26][5] ;
 wire \inst$top.soc.cpu.gprf.mem[26][6] ;
 wire \inst$top.soc.cpu.gprf.mem[26][7] ;
 wire \inst$top.soc.cpu.gprf.mem[26][8] ;
 wire \inst$top.soc.cpu.gprf.mem[26][9] ;
 wire \inst$top.soc.cpu.gprf.mem[27][0] ;
 wire \inst$top.soc.cpu.gprf.mem[27][10] ;
 wire \inst$top.soc.cpu.gprf.mem[27][11] ;
 wire \inst$top.soc.cpu.gprf.mem[27][12] ;
 wire \inst$top.soc.cpu.gprf.mem[27][13] ;
 wire \inst$top.soc.cpu.gprf.mem[27][14] ;
 wire \inst$top.soc.cpu.gprf.mem[27][15] ;
 wire \inst$top.soc.cpu.gprf.mem[27][16] ;
 wire \inst$top.soc.cpu.gprf.mem[27][17] ;
 wire \inst$top.soc.cpu.gprf.mem[27][18] ;
 wire \inst$top.soc.cpu.gprf.mem[27][19] ;
 wire \inst$top.soc.cpu.gprf.mem[27][1] ;
 wire \inst$top.soc.cpu.gprf.mem[27][20] ;
 wire \inst$top.soc.cpu.gprf.mem[27][21] ;
 wire \inst$top.soc.cpu.gprf.mem[27][22] ;
 wire \inst$top.soc.cpu.gprf.mem[27][23] ;
 wire \inst$top.soc.cpu.gprf.mem[27][24] ;
 wire \inst$top.soc.cpu.gprf.mem[27][25] ;
 wire \inst$top.soc.cpu.gprf.mem[27][26] ;
 wire \inst$top.soc.cpu.gprf.mem[27][27] ;
 wire \inst$top.soc.cpu.gprf.mem[27][28] ;
 wire \inst$top.soc.cpu.gprf.mem[27][29] ;
 wire \inst$top.soc.cpu.gprf.mem[27][2] ;
 wire \inst$top.soc.cpu.gprf.mem[27][30] ;
 wire \inst$top.soc.cpu.gprf.mem[27][31] ;
 wire \inst$top.soc.cpu.gprf.mem[27][3] ;
 wire \inst$top.soc.cpu.gprf.mem[27][4] ;
 wire \inst$top.soc.cpu.gprf.mem[27][5] ;
 wire \inst$top.soc.cpu.gprf.mem[27][6] ;
 wire \inst$top.soc.cpu.gprf.mem[27][7] ;
 wire \inst$top.soc.cpu.gprf.mem[27][8] ;
 wire \inst$top.soc.cpu.gprf.mem[27][9] ;
 wire \inst$top.soc.cpu.gprf.mem[28][0] ;
 wire \inst$top.soc.cpu.gprf.mem[28][10] ;
 wire \inst$top.soc.cpu.gprf.mem[28][11] ;
 wire \inst$top.soc.cpu.gprf.mem[28][12] ;
 wire \inst$top.soc.cpu.gprf.mem[28][13] ;
 wire \inst$top.soc.cpu.gprf.mem[28][14] ;
 wire \inst$top.soc.cpu.gprf.mem[28][15] ;
 wire \inst$top.soc.cpu.gprf.mem[28][16] ;
 wire \inst$top.soc.cpu.gprf.mem[28][17] ;
 wire \inst$top.soc.cpu.gprf.mem[28][18] ;
 wire \inst$top.soc.cpu.gprf.mem[28][19] ;
 wire \inst$top.soc.cpu.gprf.mem[28][1] ;
 wire \inst$top.soc.cpu.gprf.mem[28][20] ;
 wire \inst$top.soc.cpu.gprf.mem[28][21] ;
 wire \inst$top.soc.cpu.gprf.mem[28][22] ;
 wire \inst$top.soc.cpu.gprf.mem[28][23] ;
 wire \inst$top.soc.cpu.gprf.mem[28][24] ;
 wire \inst$top.soc.cpu.gprf.mem[28][25] ;
 wire \inst$top.soc.cpu.gprf.mem[28][26] ;
 wire \inst$top.soc.cpu.gprf.mem[28][27] ;
 wire \inst$top.soc.cpu.gprf.mem[28][28] ;
 wire \inst$top.soc.cpu.gprf.mem[28][29] ;
 wire \inst$top.soc.cpu.gprf.mem[28][2] ;
 wire \inst$top.soc.cpu.gprf.mem[28][30] ;
 wire \inst$top.soc.cpu.gprf.mem[28][31] ;
 wire \inst$top.soc.cpu.gprf.mem[28][3] ;
 wire \inst$top.soc.cpu.gprf.mem[28][4] ;
 wire \inst$top.soc.cpu.gprf.mem[28][5] ;
 wire \inst$top.soc.cpu.gprf.mem[28][6] ;
 wire \inst$top.soc.cpu.gprf.mem[28][7] ;
 wire \inst$top.soc.cpu.gprf.mem[28][8] ;
 wire \inst$top.soc.cpu.gprf.mem[28][9] ;
 wire \inst$top.soc.cpu.gprf.mem[29][0] ;
 wire \inst$top.soc.cpu.gprf.mem[29][10] ;
 wire \inst$top.soc.cpu.gprf.mem[29][11] ;
 wire \inst$top.soc.cpu.gprf.mem[29][12] ;
 wire \inst$top.soc.cpu.gprf.mem[29][13] ;
 wire \inst$top.soc.cpu.gprf.mem[29][14] ;
 wire \inst$top.soc.cpu.gprf.mem[29][15] ;
 wire \inst$top.soc.cpu.gprf.mem[29][16] ;
 wire \inst$top.soc.cpu.gprf.mem[29][17] ;
 wire \inst$top.soc.cpu.gprf.mem[29][18] ;
 wire \inst$top.soc.cpu.gprf.mem[29][19] ;
 wire \inst$top.soc.cpu.gprf.mem[29][1] ;
 wire \inst$top.soc.cpu.gprf.mem[29][20] ;
 wire \inst$top.soc.cpu.gprf.mem[29][21] ;
 wire \inst$top.soc.cpu.gprf.mem[29][22] ;
 wire \inst$top.soc.cpu.gprf.mem[29][23] ;
 wire \inst$top.soc.cpu.gprf.mem[29][24] ;
 wire \inst$top.soc.cpu.gprf.mem[29][25] ;
 wire \inst$top.soc.cpu.gprf.mem[29][26] ;
 wire \inst$top.soc.cpu.gprf.mem[29][27] ;
 wire \inst$top.soc.cpu.gprf.mem[29][28] ;
 wire \inst$top.soc.cpu.gprf.mem[29][29] ;
 wire \inst$top.soc.cpu.gprf.mem[29][2] ;
 wire \inst$top.soc.cpu.gprf.mem[29][30] ;
 wire \inst$top.soc.cpu.gprf.mem[29][31] ;
 wire \inst$top.soc.cpu.gprf.mem[29][3] ;
 wire \inst$top.soc.cpu.gprf.mem[29][4] ;
 wire \inst$top.soc.cpu.gprf.mem[29][5] ;
 wire \inst$top.soc.cpu.gprf.mem[29][6] ;
 wire \inst$top.soc.cpu.gprf.mem[29][7] ;
 wire \inst$top.soc.cpu.gprf.mem[29][8] ;
 wire \inst$top.soc.cpu.gprf.mem[29][9] ;
 wire \inst$top.soc.cpu.gprf.mem[2][0] ;
 wire \inst$top.soc.cpu.gprf.mem[2][10] ;
 wire \inst$top.soc.cpu.gprf.mem[2][11] ;
 wire \inst$top.soc.cpu.gprf.mem[2][12] ;
 wire \inst$top.soc.cpu.gprf.mem[2][13] ;
 wire \inst$top.soc.cpu.gprf.mem[2][14] ;
 wire \inst$top.soc.cpu.gprf.mem[2][15] ;
 wire \inst$top.soc.cpu.gprf.mem[2][16] ;
 wire \inst$top.soc.cpu.gprf.mem[2][17] ;
 wire \inst$top.soc.cpu.gprf.mem[2][18] ;
 wire \inst$top.soc.cpu.gprf.mem[2][19] ;
 wire \inst$top.soc.cpu.gprf.mem[2][1] ;
 wire \inst$top.soc.cpu.gprf.mem[2][20] ;
 wire \inst$top.soc.cpu.gprf.mem[2][21] ;
 wire \inst$top.soc.cpu.gprf.mem[2][22] ;
 wire \inst$top.soc.cpu.gprf.mem[2][23] ;
 wire \inst$top.soc.cpu.gprf.mem[2][24] ;
 wire \inst$top.soc.cpu.gprf.mem[2][25] ;
 wire \inst$top.soc.cpu.gprf.mem[2][26] ;
 wire \inst$top.soc.cpu.gprf.mem[2][27] ;
 wire \inst$top.soc.cpu.gprf.mem[2][28] ;
 wire \inst$top.soc.cpu.gprf.mem[2][29] ;
 wire \inst$top.soc.cpu.gprf.mem[2][2] ;
 wire \inst$top.soc.cpu.gprf.mem[2][30] ;
 wire \inst$top.soc.cpu.gprf.mem[2][31] ;
 wire \inst$top.soc.cpu.gprf.mem[2][3] ;
 wire \inst$top.soc.cpu.gprf.mem[2][4] ;
 wire \inst$top.soc.cpu.gprf.mem[2][5] ;
 wire \inst$top.soc.cpu.gprf.mem[2][6] ;
 wire \inst$top.soc.cpu.gprf.mem[2][7] ;
 wire \inst$top.soc.cpu.gprf.mem[2][8] ;
 wire \inst$top.soc.cpu.gprf.mem[2][9] ;
 wire \inst$top.soc.cpu.gprf.mem[30][0] ;
 wire \inst$top.soc.cpu.gprf.mem[30][10] ;
 wire \inst$top.soc.cpu.gprf.mem[30][11] ;
 wire \inst$top.soc.cpu.gprf.mem[30][12] ;
 wire \inst$top.soc.cpu.gprf.mem[30][13] ;
 wire \inst$top.soc.cpu.gprf.mem[30][14] ;
 wire \inst$top.soc.cpu.gprf.mem[30][15] ;
 wire \inst$top.soc.cpu.gprf.mem[30][16] ;
 wire \inst$top.soc.cpu.gprf.mem[30][17] ;
 wire \inst$top.soc.cpu.gprf.mem[30][18] ;
 wire \inst$top.soc.cpu.gprf.mem[30][19] ;
 wire \inst$top.soc.cpu.gprf.mem[30][1] ;
 wire \inst$top.soc.cpu.gprf.mem[30][20] ;
 wire \inst$top.soc.cpu.gprf.mem[30][21] ;
 wire \inst$top.soc.cpu.gprf.mem[30][22] ;
 wire \inst$top.soc.cpu.gprf.mem[30][23] ;
 wire \inst$top.soc.cpu.gprf.mem[30][24] ;
 wire \inst$top.soc.cpu.gprf.mem[30][25] ;
 wire \inst$top.soc.cpu.gprf.mem[30][26] ;
 wire \inst$top.soc.cpu.gprf.mem[30][27] ;
 wire \inst$top.soc.cpu.gprf.mem[30][28] ;
 wire \inst$top.soc.cpu.gprf.mem[30][29] ;
 wire \inst$top.soc.cpu.gprf.mem[30][2] ;
 wire \inst$top.soc.cpu.gprf.mem[30][30] ;
 wire \inst$top.soc.cpu.gprf.mem[30][31] ;
 wire \inst$top.soc.cpu.gprf.mem[30][3] ;
 wire \inst$top.soc.cpu.gprf.mem[30][4] ;
 wire \inst$top.soc.cpu.gprf.mem[30][5] ;
 wire \inst$top.soc.cpu.gprf.mem[30][6] ;
 wire \inst$top.soc.cpu.gprf.mem[30][7] ;
 wire \inst$top.soc.cpu.gprf.mem[30][8] ;
 wire \inst$top.soc.cpu.gprf.mem[30][9] ;
 wire \inst$top.soc.cpu.gprf.mem[31][0] ;
 wire \inst$top.soc.cpu.gprf.mem[31][10] ;
 wire \inst$top.soc.cpu.gprf.mem[31][11] ;
 wire \inst$top.soc.cpu.gprf.mem[31][12] ;
 wire \inst$top.soc.cpu.gprf.mem[31][13] ;
 wire \inst$top.soc.cpu.gprf.mem[31][14] ;
 wire \inst$top.soc.cpu.gprf.mem[31][15] ;
 wire \inst$top.soc.cpu.gprf.mem[31][16] ;
 wire \inst$top.soc.cpu.gprf.mem[31][17] ;
 wire \inst$top.soc.cpu.gprf.mem[31][18] ;
 wire \inst$top.soc.cpu.gprf.mem[31][19] ;
 wire \inst$top.soc.cpu.gprf.mem[31][1] ;
 wire \inst$top.soc.cpu.gprf.mem[31][20] ;
 wire \inst$top.soc.cpu.gprf.mem[31][21] ;
 wire \inst$top.soc.cpu.gprf.mem[31][22] ;
 wire \inst$top.soc.cpu.gprf.mem[31][23] ;
 wire \inst$top.soc.cpu.gprf.mem[31][24] ;
 wire \inst$top.soc.cpu.gprf.mem[31][25] ;
 wire \inst$top.soc.cpu.gprf.mem[31][26] ;
 wire \inst$top.soc.cpu.gprf.mem[31][27] ;
 wire \inst$top.soc.cpu.gprf.mem[31][28] ;
 wire \inst$top.soc.cpu.gprf.mem[31][29] ;
 wire \inst$top.soc.cpu.gprf.mem[31][2] ;
 wire \inst$top.soc.cpu.gprf.mem[31][30] ;
 wire \inst$top.soc.cpu.gprf.mem[31][31] ;
 wire \inst$top.soc.cpu.gprf.mem[31][3] ;
 wire \inst$top.soc.cpu.gprf.mem[31][4] ;
 wire \inst$top.soc.cpu.gprf.mem[31][5] ;
 wire \inst$top.soc.cpu.gprf.mem[31][6] ;
 wire \inst$top.soc.cpu.gprf.mem[31][7] ;
 wire \inst$top.soc.cpu.gprf.mem[31][8] ;
 wire \inst$top.soc.cpu.gprf.mem[31][9] ;
 wire \inst$top.soc.cpu.gprf.mem[3][0] ;
 wire \inst$top.soc.cpu.gprf.mem[3][10] ;
 wire \inst$top.soc.cpu.gprf.mem[3][11] ;
 wire \inst$top.soc.cpu.gprf.mem[3][12] ;
 wire \inst$top.soc.cpu.gprf.mem[3][13] ;
 wire \inst$top.soc.cpu.gprf.mem[3][14] ;
 wire \inst$top.soc.cpu.gprf.mem[3][15] ;
 wire \inst$top.soc.cpu.gprf.mem[3][16] ;
 wire \inst$top.soc.cpu.gprf.mem[3][17] ;
 wire \inst$top.soc.cpu.gprf.mem[3][18] ;
 wire \inst$top.soc.cpu.gprf.mem[3][19] ;
 wire \inst$top.soc.cpu.gprf.mem[3][1] ;
 wire \inst$top.soc.cpu.gprf.mem[3][20] ;
 wire \inst$top.soc.cpu.gprf.mem[3][21] ;
 wire \inst$top.soc.cpu.gprf.mem[3][22] ;
 wire \inst$top.soc.cpu.gprf.mem[3][23] ;
 wire \inst$top.soc.cpu.gprf.mem[3][24] ;
 wire \inst$top.soc.cpu.gprf.mem[3][25] ;
 wire \inst$top.soc.cpu.gprf.mem[3][26] ;
 wire \inst$top.soc.cpu.gprf.mem[3][27] ;
 wire \inst$top.soc.cpu.gprf.mem[3][28] ;
 wire \inst$top.soc.cpu.gprf.mem[3][29] ;
 wire \inst$top.soc.cpu.gprf.mem[3][2] ;
 wire \inst$top.soc.cpu.gprf.mem[3][30] ;
 wire \inst$top.soc.cpu.gprf.mem[3][31] ;
 wire \inst$top.soc.cpu.gprf.mem[3][3] ;
 wire \inst$top.soc.cpu.gprf.mem[3][4] ;
 wire \inst$top.soc.cpu.gprf.mem[3][5] ;
 wire \inst$top.soc.cpu.gprf.mem[3][6] ;
 wire \inst$top.soc.cpu.gprf.mem[3][7] ;
 wire \inst$top.soc.cpu.gprf.mem[3][8] ;
 wire \inst$top.soc.cpu.gprf.mem[3][9] ;
 wire \inst$top.soc.cpu.gprf.mem[4][0] ;
 wire \inst$top.soc.cpu.gprf.mem[4][10] ;
 wire \inst$top.soc.cpu.gprf.mem[4][11] ;
 wire \inst$top.soc.cpu.gprf.mem[4][12] ;
 wire \inst$top.soc.cpu.gprf.mem[4][13] ;
 wire \inst$top.soc.cpu.gprf.mem[4][14] ;
 wire \inst$top.soc.cpu.gprf.mem[4][15] ;
 wire \inst$top.soc.cpu.gprf.mem[4][16] ;
 wire \inst$top.soc.cpu.gprf.mem[4][17] ;
 wire \inst$top.soc.cpu.gprf.mem[4][18] ;
 wire \inst$top.soc.cpu.gprf.mem[4][19] ;
 wire \inst$top.soc.cpu.gprf.mem[4][1] ;
 wire \inst$top.soc.cpu.gprf.mem[4][20] ;
 wire \inst$top.soc.cpu.gprf.mem[4][21] ;
 wire \inst$top.soc.cpu.gprf.mem[4][22] ;
 wire \inst$top.soc.cpu.gprf.mem[4][23] ;
 wire \inst$top.soc.cpu.gprf.mem[4][24] ;
 wire \inst$top.soc.cpu.gprf.mem[4][25] ;
 wire \inst$top.soc.cpu.gprf.mem[4][26] ;
 wire \inst$top.soc.cpu.gprf.mem[4][27] ;
 wire \inst$top.soc.cpu.gprf.mem[4][28] ;
 wire \inst$top.soc.cpu.gprf.mem[4][29] ;
 wire \inst$top.soc.cpu.gprf.mem[4][2] ;
 wire \inst$top.soc.cpu.gprf.mem[4][30] ;
 wire \inst$top.soc.cpu.gprf.mem[4][31] ;
 wire \inst$top.soc.cpu.gprf.mem[4][3] ;
 wire \inst$top.soc.cpu.gprf.mem[4][4] ;
 wire \inst$top.soc.cpu.gprf.mem[4][5] ;
 wire \inst$top.soc.cpu.gprf.mem[4][6] ;
 wire \inst$top.soc.cpu.gprf.mem[4][7] ;
 wire \inst$top.soc.cpu.gprf.mem[4][8] ;
 wire \inst$top.soc.cpu.gprf.mem[4][9] ;
 wire \inst$top.soc.cpu.gprf.mem[5][0] ;
 wire \inst$top.soc.cpu.gprf.mem[5][10] ;
 wire \inst$top.soc.cpu.gprf.mem[5][11] ;
 wire \inst$top.soc.cpu.gprf.mem[5][12] ;
 wire \inst$top.soc.cpu.gprf.mem[5][13] ;
 wire \inst$top.soc.cpu.gprf.mem[5][14] ;
 wire \inst$top.soc.cpu.gprf.mem[5][15] ;
 wire \inst$top.soc.cpu.gprf.mem[5][16] ;
 wire \inst$top.soc.cpu.gprf.mem[5][17] ;
 wire \inst$top.soc.cpu.gprf.mem[5][18] ;
 wire \inst$top.soc.cpu.gprf.mem[5][19] ;
 wire \inst$top.soc.cpu.gprf.mem[5][1] ;
 wire \inst$top.soc.cpu.gprf.mem[5][20] ;
 wire \inst$top.soc.cpu.gprf.mem[5][21] ;
 wire \inst$top.soc.cpu.gprf.mem[5][22] ;
 wire \inst$top.soc.cpu.gprf.mem[5][23] ;
 wire \inst$top.soc.cpu.gprf.mem[5][24] ;
 wire \inst$top.soc.cpu.gprf.mem[5][25] ;
 wire \inst$top.soc.cpu.gprf.mem[5][26] ;
 wire \inst$top.soc.cpu.gprf.mem[5][27] ;
 wire \inst$top.soc.cpu.gprf.mem[5][28] ;
 wire \inst$top.soc.cpu.gprf.mem[5][29] ;
 wire \inst$top.soc.cpu.gprf.mem[5][2] ;
 wire \inst$top.soc.cpu.gprf.mem[5][30] ;
 wire \inst$top.soc.cpu.gprf.mem[5][31] ;
 wire \inst$top.soc.cpu.gprf.mem[5][3] ;
 wire \inst$top.soc.cpu.gprf.mem[5][4] ;
 wire \inst$top.soc.cpu.gprf.mem[5][5] ;
 wire \inst$top.soc.cpu.gprf.mem[5][6] ;
 wire \inst$top.soc.cpu.gprf.mem[5][7] ;
 wire \inst$top.soc.cpu.gprf.mem[5][8] ;
 wire \inst$top.soc.cpu.gprf.mem[5][9] ;
 wire \inst$top.soc.cpu.gprf.mem[6][0] ;
 wire \inst$top.soc.cpu.gprf.mem[6][10] ;
 wire \inst$top.soc.cpu.gprf.mem[6][11] ;
 wire \inst$top.soc.cpu.gprf.mem[6][12] ;
 wire \inst$top.soc.cpu.gprf.mem[6][13] ;
 wire \inst$top.soc.cpu.gprf.mem[6][14] ;
 wire \inst$top.soc.cpu.gprf.mem[6][15] ;
 wire \inst$top.soc.cpu.gprf.mem[6][16] ;
 wire \inst$top.soc.cpu.gprf.mem[6][17] ;
 wire \inst$top.soc.cpu.gprf.mem[6][18] ;
 wire \inst$top.soc.cpu.gprf.mem[6][19] ;
 wire \inst$top.soc.cpu.gprf.mem[6][1] ;
 wire \inst$top.soc.cpu.gprf.mem[6][20] ;
 wire \inst$top.soc.cpu.gprf.mem[6][21] ;
 wire \inst$top.soc.cpu.gprf.mem[6][22] ;
 wire \inst$top.soc.cpu.gprf.mem[6][23] ;
 wire \inst$top.soc.cpu.gprf.mem[6][24] ;
 wire \inst$top.soc.cpu.gprf.mem[6][25] ;
 wire \inst$top.soc.cpu.gprf.mem[6][26] ;
 wire \inst$top.soc.cpu.gprf.mem[6][27] ;
 wire \inst$top.soc.cpu.gprf.mem[6][28] ;
 wire \inst$top.soc.cpu.gprf.mem[6][29] ;
 wire \inst$top.soc.cpu.gprf.mem[6][2] ;
 wire \inst$top.soc.cpu.gprf.mem[6][30] ;
 wire \inst$top.soc.cpu.gprf.mem[6][31] ;
 wire \inst$top.soc.cpu.gprf.mem[6][3] ;
 wire \inst$top.soc.cpu.gprf.mem[6][4] ;
 wire \inst$top.soc.cpu.gprf.mem[6][5] ;
 wire \inst$top.soc.cpu.gprf.mem[6][6] ;
 wire \inst$top.soc.cpu.gprf.mem[6][7] ;
 wire \inst$top.soc.cpu.gprf.mem[6][8] ;
 wire \inst$top.soc.cpu.gprf.mem[6][9] ;
 wire \inst$top.soc.cpu.gprf.mem[7][0] ;
 wire \inst$top.soc.cpu.gprf.mem[7][10] ;
 wire \inst$top.soc.cpu.gprf.mem[7][11] ;
 wire \inst$top.soc.cpu.gprf.mem[7][12] ;
 wire \inst$top.soc.cpu.gprf.mem[7][13] ;
 wire \inst$top.soc.cpu.gprf.mem[7][14] ;
 wire \inst$top.soc.cpu.gprf.mem[7][15] ;
 wire \inst$top.soc.cpu.gprf.mem[7][16] ;
 wire \inst$top.soc.cpu.gprf.mem[7][17] ;
 wire \inst$top.soc.cpu.gprf.mem[7][18] ;
 wire \inst$top.soc.cpu.gprf.mem[7][19] ;
 wire \inst$top.soc.cpu.gprf.mem[7][1] ;
 wire \inst$top.soc.cpu.gprf.mem[7][20] ;
 wire \inst$top.soc.cpu.gprf.mem[7][21] ;
 wire \inst$top.soc.cpu.gprf.mem[7][22] ;
 wire \inst$top.soc.cpu.gprf.mem[7][23] ;
 wire \inst$top.soc.cpu.gprf.mem[7][24] ;
 wire \inst$top.soc.cpu.gprf.mem[7][25] ;
 wire \inst$top.soc.cpu.gprf.mem[7][26] ;
 wire \inst$top.soc.cpu.gprf.mem[7][27] ;
 wire \inst$top.soc.cpu.gprf.mem[7][28] ;
 wire \inst$top.soc.cpu.gprf.mem[7][29] ;
 wire \inst$top.soc.cpu.gprf.mem[7][2] ;
 wire \inst$top.soc.cpu.gprf.mem[7][30] ;
 wire \inst$top.soc.cpu.gprf.mem[7][31] ;
 wire \inst$top.soc.cpu.gprf.mem[7][3] ;
 wire \inst$top.soc.cpu.gprf.mem[7][4] ;
 wire \inst$top.soc.cpu.gprf.mem[7][5] ;
 wire \inst$top.soc.cpu.gprf.mem[7][6] ;
 wire \inst$top.soc.cpu.gprf.mem[7][7] ;
 wire \inst$top.soc.cpu.gprf.mem[7][8] ;
 wire \inst$top.soc.cpu.gprf.mem[7][9] ;
 wire \inst$top.soc.cpu.gprf.mem[8][0] ;
 wire \inst$top.soc.cpu.gprf.mem[8][10] ;
 wire \inst$top.soc.cpu.gprf.mem[8][11] ;
 wire \inst$top.soc.cpu.gprf.mem[8][12] ;
 wire \inst$top.soc.cpu.gprf.mem[8][13] ;
 wire \inst$top.soc.cpu.gprf.mem[8][14] ;
 wire \inst$top.soc.cpu.gprf.mem[8][15] ;
 wire \inst$top.soc.cpu.gprf.mem[8][16] ;
 wire \inst$top.soc.cpu.gprf.mem[8][17] ;
 wire \inst$top.soc.cpu.gprf.mem[8][18] ;
 wire \inst$top.soc.cpu.gprf.mem[8][19] ;
 wire \inst$top.soc.cpu.gprf.mem[8][1] ;
 wire \inst$top.soc.cpu.gprf.mem[8][20] ;
 wire \inst$top.soc.cpu.gprf.mem[8][21] ;
 wire \inst$top.soc.cpu.gprf.mem[8][22] ;
 wire \inst$top.soc.cpu.gprf.mem[8][23] ;
 wire \inst$top.soc.cpu.gprf.mem[8][24] ;
 wire \inst$top.soc.cpu.gprf.mem[8][25] ;
 wire \inst$top.soc.cpu.gprf.mem[8][26] ;
 wire \inst$top.soc.cpu.gprf.mem[8][27] ;
 wire \inst$top.soc.cpu.gprf.mem[8][28] ;
 wire \inst$top.soc.cpu.gprf.mem[8][29] ;
 wire \inst$top.soc.cpu.gprf.mem[8][2] ;
 wire \inst$top.soc.cpu.gprf.mem[8][30] ;
 wire \inst$top.soc.cpu.gprf.mem[8][31] ;
 wire \inst$top.soc.cpu.gprf.mem[8][3] ;
 wire \inst$top.soc.cpu.gprf.mem[8][4] ;
 wire \inst$top.soc.cpu.gprf.mem[8][5] ;
 wire \inst$top.soc.cpu.gprf.mem[8][6] ;
 wire \inst$top.soc.cpu.gprf.mem[8][7] ;
 wire \inst$top.soc.cpu.gprf.mem[8][8] ;
 wire \inst$top.soc.cpu.gprf.mem[8][9] ;
 wire \inst$top.soc.cpu.gprf.mem[9][0] ;
 wire \inst$top.soc.cpu.gprf.mem[9][10] ;
 wire \inst$top.soc.cpu.gprf.mem[9][11] ;
 wire \inst$top.soc.cpu.gprf.mem[9][12] ;
 wire \inst$top.soc.cpu.gprf.mem[9][13] ;
 wire \inst$top.soc.cpu.gprf.mem[9][14] ;
 wire \inst$top.soc.cpu.gprf.mem[9][15] ;
 wire \inst$top.soc.cpu.gprf.mem[9][16] ;
 wire \inst$top.soc.cpu.gprf.mem[9][17] ;
 wire \inst$top.soc.cpu.gprf.mem[9][18] ;
 wire \inst$top.soc.cpu.gprf.mem[9][19] ;
 wire \inst$top.soc.cpu.gprf.mem[9][1] ;
 wire \inst$top.soc.cpu.gprf.mem[9][20] ;
 wire \inst$top.soc.cpu.gprf.mem[9][21] ;
 wire \inst$top.soc.cpu.gprf.mem[9][22] ;
 wire \inst$top.soc.cpu.gprf.mem[9][23] ;
 wire \inst$top.soc.cpu.gprf.mem[9][24] ;
 wire \inst$top.soc.cpu.gprf.mem[9][25] ;
 wire \inst$top.soc.cpu.gprf.mem[9][26] ;
 wire \inst$top.soc.cpu.gprf.mem[9][27] ;
 wire \inst$top.soc.cpu.gprf.mem[9][28] ;
 wire \inst$top.soc.cpu.gprf.mem[9][29] ;
 wire \inst$top.soc.cpu.gprf.mem[9][2] ;
 wire \inst$top.soc.cpu.gprf.mem[9][30] ;
 wire \inst$top.soc.cpu.gprf.mem[9][31] ;
 wire \inst$top.soc.cpu.gprf.mem[9][3] ;
 wire \inst$top.soc.cpu.gprf.mem[9][4] ;
 wire \inst$top.soc.cpu.gprf.mem[9][5] ;
 wire \inst$top.soc.cpu.gprf.mem[9][6] ;
 wire \inst$top.soc.cpu.gprf.mem[9][7] ;
 wire \inst$top.soc.cpu.gprf.mem[9][8] ;
 wire \inst$top.soc.cpu.gprf.mem[9][9] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[0] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[10] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[11] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[12] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[13] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[14] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[15] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[16] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[17] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[18] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[19] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[1] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[20] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[21] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[22] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[23] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[24] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[25] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[26] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[27] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[28] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[29] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[2] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[30] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[31] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[3] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[4] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[5] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[6] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[7] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[8] ;
 wire \inst$top.soc.cpu.gprf.mem_rp1__data[9] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[0] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[10] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[11] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[12] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[13] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[14] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[15] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[16] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[17] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[18] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[19] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[1] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[20] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[21] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[22] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[23] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[24] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[25] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[26] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[27] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[28] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[29] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[2] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[30] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[31] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[3] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[4] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[5] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[6] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[7] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[8] ;
 wire \inst$top.soc.cpu.gprf.mem_rp2__data[9] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[0] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[10] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[11] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[12] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[13] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[14] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[15] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[16] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[17] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[18] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[19] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[1] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[20] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[21] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[22] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[23] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[24] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[25] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[26] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[27] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[28] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[29] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[2] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[30] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[31] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[3] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[4] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[5] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[6] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[7] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[8] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_data[9] ;
 wire \inst$top.soc.cpu.gprf.x_bypass1_raw ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[0] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[10] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[11] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[12] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[13] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[14] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[15] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[16] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[17] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[18] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[19] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[1] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[20] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[21] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[22] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[23] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[24] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[25] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[26] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[27] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[28] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[29] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[2] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[30] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[31] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[3] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[4] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[5] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[6] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[7] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[8] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_data[9] ;
 wire \inst$top.soc.cpu.gprf.x_bypass2_raw ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[0] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[10] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[11] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[12] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[13] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[14] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[15] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[16] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[17] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[18] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[19] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[1] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[20] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[21] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[22] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[23] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[24] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[25] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[26] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[27] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[28] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[29] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[2] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[3] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[4] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[5] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[6] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[7] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[8] ;
 wire \inst$top.soc.cpu.loadstore.dbus__adr[9] ;
 wire \inst$top.soc.cpu.loadstore.dbus__cyc ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[0] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[10] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[11] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[12] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[13] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[14] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[15] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[16] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[17] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[18] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[19] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[1] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[20] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[21] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[22] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[23] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[24] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[25] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[26] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[27] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[28] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[29] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[2] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[30] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[31] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[3] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[4] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[5] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[6] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[7] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[8] ;
 wire \inst$top.soc.cpu.loadstore.dbus__dat_w[9] ;
 wire \inst$top.soc.cpu.loadstore.dbus__sel[0] ;
 wire \inst$top.soc.cpu.loadstore.dbus__sel[1] ;
 wire \inst$top.soc.cpu.loadstore.dbus__sel[2] ;
 wire \inst$top.soc.cpu.loadstore.dbus__sel[3] ;
 wire \inst$top.soc.cpu.loadstore.dbus__stb ;
 wire \inst$top.soc.cpu.loadstore.dbus__we ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[0] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[10] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[11] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[12] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[13] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[14] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[15] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[16] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[17] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[18] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[19] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[1] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[20] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[21] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[22] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[23] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[24] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[25] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[26] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[27] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[28] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[29] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[2] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[30] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[31] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[3] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[4] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[5] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[6] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[7] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[8] ;
 wire \inst$top.soc.cpu.loadstore.m_load_data[9] ;
 wire \inst$top.soc.cpu.m.source__valid ;
 wire \inst$top.soc.cpu.multiplier.m_low ;
 wire \inst$top.soc.cpu.multiplier.m_prod[0] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[10] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[11] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[12] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[13] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[14] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[15] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[16] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[17] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[18] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[19] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[1] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[20] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[21] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[22] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[23] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[24] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[25] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[26] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[27] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[28] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[29] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[2] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[30] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[31] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[32] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[33] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[34] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[35] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[36] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[37] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[38] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[39] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[3] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[40] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[41] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[42] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[43] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[44] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[45] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[46] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[47] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[48] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[49] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[4] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[50] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[51] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[52] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[53] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[54] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[55] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[56] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[57] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[58] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[59] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[5] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[60] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[61] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[62] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[63] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[6] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[7] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[8] ;
 wire \inst$top.soc.cpu.multiplier.m_prod[9] ;
 wire \inst$top.soc.cpu.multiplier.w_result[0] ;
 wire \inst$top.soc.cpu.multiplier.w_result[10] ;
 wire \inst$top.soc.cpu.multiplier.w_result[11] ;
 wire \inst$top.soc.cpu.multiplier.w_result[12] ;
 wire \inst$top.soc.cpu.multiplier.w_result[13] ;
 wire \inst$top.soc.cpu.multiplier.w_result[14] ;
 wire \inst$top.soc.cpu.multiplier.w_result[15] ;
 wire \inst$top.soc.cpu.multiplier.w_result[16] ;
 wire \inst$top.soc.cpu.multiplier.w_result[17] ;
 wire \inst$top.soc.cpu.multiplier.w_result[18] ;
 wire \inst$top.soc.cpu.multiplier.w_result[19] ;
 wire \inst$top.soc.cpu.multiplier.w_result[1] ;
 wire \inst$top.soc.cpu.multiplier.w_result[20] ;
 wire \inst$top.soc.cpu.multiplier.w_result[21] ;
 wire \inst$top.soc.cpu.multiplier.w_result[22] ;
 wire \inst$top.soc.cpu.multiplier.w_result[23] ;
 wire \inst$top.soc.cpu.multiplier.w_result[24] ;
 wire \inst$top.soc.cpu.multiplier.w_result[25] ;
 wire \inst$top.soc.cpu.multiplier.w_result[26] ;
 wire \inst$top.soc.cpu.multiplier.w_result[27] ;
 wire \inst$top.soc.cpu.multiplier.w_result[28] ;
 wire \inst$top.soc.cpu.multiplier.w_result[29] ;
 wire \inst$top.soc.cpu.multiplier.w_result[2] ;
 wire \inst$top.soc.cpu.multiplier.w_result[30] ;
 wire \inst$top.soc.cpu.multiplier.w_result[31] ;
 wire \inst$top.soc.cpu.multiplier.w_result[3] ;
 wire \inst$top.soc.cpu.multiplier.w_result[4] ;
 wire \inst$top.soc.cpu.multiplier.w_result[5] ;
 wire \inst$top.soc.cpu.multiplier.w_result[6] ;
 wire \inst$top.soc.cpu.multiplier.w_result[7] ;
 wire \inst$top.soc.cpu.multiplier.w_result[8] ;
 wire \inst$top.soc.cpu.multiplier.w_result[9] ;
 wire \inst$top.soc.cpu.multiplier.x_low ;
 wire \inst$top.soc.cpu.multiplier.x_prod[0] ;
 wire \inst$top.soc.cpu.multiplier.x_prod[1] ;
 wire \inst$top.soc.cpu.multiplier.x_prod[2] ;
 wire \inst$top.soc.cpu.multiplier.x_prod[3] ;
 wire \inst$top.soc.cpu.multiplier.x_prod[4] ;
 wire \inst$top.soc.cpu.multiplier.x_prod[5] ;
 wire \inst$top.soc.cpu.multiplier.x_prod[6] ;
 wire \inst$top.soc.cpu.multiplier.x_src1_signed ;
 wire \inst$top.soc.cpu.multiplier.x_src2_signed ;
 wire \inst$top.soc.cpu.shifter.m_direction ;
 wire \inst$top.soc.cpu.shifter.m_result$7[0] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[10] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[11] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[12] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[13] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[14] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[15] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[16] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[17] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[18] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[19] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[1] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[20] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[21] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[22] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[23] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[24] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[25] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[26] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[27] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[28] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[29] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[2] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[30] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[31] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[3] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[4] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[5] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[6] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[7] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[8] ;
 wire \inst$top.soc.cpu.shifter.m_result$7[9] ;
 wire \inst$top.soc.cpu.sink__payload$12[100] ;
 wire \inst$top.soc.cpu.sink__payload$12[101] ;
 wire \inst$top.soc.cpu.sink__payload$12[102] ;
 wire \inst$top.soc.cpu.sink__payload$12[103] ;
 wire \inst$top.soc.cpu.sink__payload$12[104] ;
 wire \inst$top.soc.cpu.sink__payload$12[105] ;
 wire \inst$top.soc.cpu.sink__payload$12[109] ;
 wire \inst$top.soc.cpu.sink__payload$12[10] ;
 wire \inst$top.soc.cpu.sink__payload$12[110] ;
 wire \inst$top.soc.cpu.sink__payload$12[111] ;
 wire \inst$top.soc.cpu.sink__payload$12[112] ;
 wire \inst$top.soc.cpu.sink__payload$12[113] ;
 wire \inst$top.soc.cpu.sink__payload$12[114] ;
 wire \inst$top.soc.cpu.sink__payload$12[115] ;
 wire \inst$top.soc.cpu.sink__payload$12[116] ;
 wire \inst$top.soc.cpu.sink__payload$12[117] ;
 wire \inst$top.soc.cpu.sink__payload$12[118] ;
 wire \inst$top.soc.cpu.sink__payload$12[119] ;
 wire \inst$top.soc.cpu.sink__payload$12[11] ;
 wire \inst$top.soc.cpu.sink__payload$12[120] ;
 wire \inst$top.soc.cpu.sink__payload$12[121] ;
 wire \inst$top.soc.cpu.sink__payload$12[122] ;
 wire \inst$top.soc.cpu.sink__payload$12[123] ;
 wire \inst$top.soc.cpu.sink__payload$12[124] ;
 wire \inst$top.soc.cpu.sink__payload$12[125] ;
 wire \inst$top.soc.cpu.sink__payload$12[126] ;
 wire \inst$top.soc.cpu.sink__payload$12[127] ;
 wire \inst$top.soc.cpu.sink__payload$12[128] ;
 wire \inst$top.soc.cpu.sink__payload$12[129] ;
 wire \inst$top.soc.cpu.sink__payload$12[12] ;
 wire \inst$top.soc.cpu.sink__payload$12[130] ;
 wire \inst$top.soc.cpu.sink__payload$12[131] ;
 wire \inst$top.soc.cpu.sink__payload$12[132] ;
 wire \inst$top.soc.cpu.sink__payload$12[133] ;
 wire \inst$top.soc.cpu.sink__payload$12[134] ;
 wire \inst$top.soc.cpu.sink__payload$12[135] ;
 wire \inst$top.soc.cpu.sink__payload$12[136] ;
 wire \inst$top.soc.cpu.sink__payload$12[137] ;
 wire \inst$top.soc.cpu.sink__payload$12[138] ;
 wire \inst$top.soc.cpu.sink__payload$12[139] ;
 wire \inst$top.soc.cpu.sink__payload$12[13] ;
 wire \inst$top.soc.cpu.sink__payload$12[140] ;
 wire \inst$top.soc.cpu.sink__payload$12[143] ;
 wire \inst$top.soc.cpu.sink__payload$12[144] ;
 wire \inst$top.soc.cpu.sink__payload$12[14] ;
 wire \inst$top.soc.cpu.sink__payload$12[15] ;
 wire \inst$top.soc.cpu.sink__payload$12[162] ;
 wire \inst$top.soc.cpu.sink__payload$12[163] ;
 wire \inst$top.soc.cpu.sink__payload$12[164] ;
 wire \inst$top.soc.cpu.sink__payload$12[165] ;
 wire \inst$top.soc.cpu.sink__payload$12[166] ;
 wire \inst$top.soc.cpu.sink__payload$12[167] ;
 wire \inst$top.soc.cpu.sink__payload$12[168] ;
 wire \inst$top.soc.cpu.sink__payload$12[169] ;
 wire \inst$top.soc.cpu.sink__payload$12[16] ;
 wire \inst$top.soc.cpu.sink__payload$12[170] ;
 wire \inst$top.soc.cpu.sink__payload$12[171] ;
 wire \inst$top.soc.cpu.sink__payload$12[172] ;
 wire \inst$top.soc.cpu.sink__payload$12[173] ;
 wire \inst$top.soc.cpu.sink__payload$12[174] ;
 wire \inst$top.soc.cpu.sink__payload$12[175] ;
 wire \inst$top.soc.cpu.sink__payload$12[176] ;
 wire \inst$top.soc.cpu.sink__payload$12[177] ;
 wire \inst$top.soc.cpu.sink__payload$12[178] ;
 wire \inst$top.soc.cpu.sink__payload$12[179] ;
 wire \inst$top.soc.cpu.sink__payload$12[17] ;
 wire \inst$top.soc.cpu.sink__payload$12[180] ;
 wire \inst$top.soc.cpu.sink__payload$12[181] ;
 wire \inst$top.soc.cpu.sink__payload$12[182] ;
 wire \inst$top.soc.cpu.sink__payload$12[183] ;
 wire \inst$top.soc.cpu.sink__payload$12[184] ;
 wire \inst$top.soc.cpu.sink__payload$12[185] ;
 wire \inst$top.soc.cpu.sink__payload$12[186] ;
 wire \inst$top.soc.cpu.sink__payload$12[187] ;
 wire \inst$top.soc.cpu.sink__payload$12[188] ;
 wire \inst$top.soc.cpu.sink__payload$12[189] ;
 wire \inst$top.soc.cpu.sink__payload$12[18] ;
 wire \inst$top.soc.cpu.sink__payload$12[190] ;
 wire \inst$top.soc.cpu.sink__payload$12[191] ;
 wire \inst$top.soc.cpu.sink__payload$12[19] ;
 wire \inst$top.soc.cpu.sink__payload$12[20] ;
 wire \inst$top.soc.cpu.sink__payload$12[21] ;
 wire \inst$top.soc.cpu.sink__payload$12[22] ;
 wire \inst$top.soc.cpu.sink__payload$12[23] ;
 wire \inst$top.soc.cpu.sink__payload$12[24] ;
 wire \inst$top.soc.cpu.sink__payload$12[25] ;
 wire \inst$top.soc.cpu.sink__payload$12[26] ;
 wire \inst$top.soc.cpu.sink__payload$12[27] ;
 wire \inst$top.soc.cpu.sink__payload$12[28] ;
 wire \inst$top.soc.cpu.sink__payload$12[29] ;
 wire \inst$top.soc.cpu.sink__payload$12[2] ;
 wire \inst$top.soc.cpu.sink__payload$12[30] ;
 wire \inst$top.soc.cpu.sink__payload$12[31] ;
 wire \inst$top.soc.cpu.sink__payload$12[32] ;
 wire \inst$top.soc.cpu.sink__payload$12[33] ;
 wire \inst$top.soc.cpu.sink__payload$12[34] ;
 wire \inst$top.soc.cpu.sink__payload$12[35] ;
 wire \inst$top.soc.cpu.sink__payload$12[36] ;
 wire \inst$top.soc.cpu.sink__payload$12[37] ;
 wire \inst$top.soc.cpu.sink__payload$12[38] ;
 wire \inst$top.soc.cpu.sink__payload$12[39] ;
 wire \inst$top.soc.cpu.sink__payload$12[3] ;
 wire \inst$top.soc.cpu.sink__payload$12[40] ;
 wire \inst$top.soc.cpu.sink__payload$12[41] ;
 wire \inst$top.soc.cpu.sink__payload$12[42] ;
 wire \inst$top.soc.cpu.sink__payload$12[4] ;
 wire \inst$top.soc.cpu.sink__payload$12[52] ;
 wire \inst$top.soc.cpu.sink__payload$12[53] ;
 wire \inst$top.soc.cpu.sink__payload$12[54] ;
 wire \inst$top.soc.cpu.sink__payload$12[55] ;
 wire \inst$top.soc.cpu.sink__payload$12[56] ;
 wire \inst$top.soc.cpu.sink__payload$12[57] ;
 wire \inst$top.soc.cpu.sink__payload$12[58] ;
 wire \inst$top.soc.cpu.sink__payload$12[59] ;
 wire \inst$top.soc.cpu.sink__payload$12[5] ;
 wire \inst$top.soc.cpu.sink__payload$12[60] ;
 wire \inst$top.soc.cpu.sink__payload$12[61] ;
 wire \inst$top.soc.cpu.sink__payload$12[62] ;
 wire \inst$top.soc.cpu.sink__payload$12[63] ;
 wire \inst$top.soc.cpu.sink__payload$12[6] ;
 wire \inst$top.soc.cpu.sink__payload$12[7] ;
 wire \inst$top.soc.cpu.sink__payload$12[8] ;
 wire \inst$top.soc.cpu.sink__payload$12[9] ;
 wire \inst$top.soc.cpu.sink__payload$18[100] ;
 wire \inst$top.soc.cpu.sink__payload$18[101] ;
 wire \inst$top.soc.cpu.sink__payload$18[102] ;
 wire \inst$top.soc.cpu.sink__payload$18[103] ;
 wire \inst$top.soc.cpu.sink__payload$18[106] ;
 wire \inst$top.soc.cpu.sink__payload$18[107] ;
 wire \inst$top.soc.cpu.sink__payload$18[108] ;
 wire \inst$top.soc.cpu.sink__payload$18[109] ;
 wire \inst$top.soc.cpu.sink__payload$18[10] ;
 wire \inst$top.soc.cpu.sink__payload$18[110] ;
 wire \inst$top.soc.cpu.sink__payload$18[111] ;
 wire \inst$top.soc.cpu.sink__payload$18[112] ;
 wire \inst$top.soc.cpu.sink__payload$18[113] ;
 wire \inst$top.soc.cpu.sink__payload$18[114] ;
 wire \inst$top.soc.cpu.sink__payload$18[115] ;
 wire \inst$top.soc.cpu.sink__payload$18[116] ;
 wire \inst$top.soc.cpu.sink__payload$18[117] ;
 wire \inst$top.soc.cpu.sink__payload$18[118] ;
 wire \inst$top.soc.cpu.sink__payload$18[119] ;
 wire \inst$top.soc.cpu.sink__payload$18[11] ;
 wire \inst$top.soc.cpu.sink__payload$18[120] ;
 wire \inst$top.soc.cpu.sink__payload$18[121] ;
 wire \inst$top.soc.cpu.sink__payload$18[122] ;
 wire \inst$top.soc.cpu.sink__payload$18[123] ;
 wire \inst$top.soc.cpu.sink__payload$18[124] ;
 wire \inst$top.soc.cpu.sink__payload$18[125] ;
 wire \inst$top.soc.cpu.sink__payload$18[126] ;
 wire \inst$top.soc.cpu.sink__payload$18[127] ;
 wire \inst$top.soc.cpu.sink__payload$18[128] ;
 wire \inst$top.soc.cpu.sink__payload$18[129] ;
 wire \inst$top.soc.cpu.sink__payload$18[12] ;
 wire \inst$top.soc.cpu.sink__payload$18[130] ;
 wire \inst$top.soc.cpu.sink__payload$18[131] ;
 wire \inst$top.soc.cpu.sink__payload$18[132] ;
 wire \inst$top.soc.cpu.sink__payload$18[133] ;
 wire \inst$top.soc.cpu.sink__payload$18[134] ;
 wire \inst$top.soc.cpu.sink__payload$18[135] ;
 wire \inst$top.soc.cpu.sink__payload$18[136] ;
 wire \inst$top.soc.cpu.sink__payload$18[137] ;
 wire \inst$top.soc.cpu.sink__payload$18[138] ;
 wire \inst$top.soc.cpu.sink__payload$18[139] ;
 wire \inst$top.soc.cpu.sink__payload$18[13] ;
 wire \inst$top.soc.cpu.sink__payload$18[140] ;
 wire \inst$top.soc.cpu.sink__payload$18[14] ;
 wire \inst$top.soc.cpu.sink__payload$18[15] ;
 wire \inst$top.soc.cpu.sink__payload$18[16] ;
 wire \inst$top.soc.cpu.sink__payload$18[17] ;
 wire \inst$top.soc.cpu.sink__payload$18[180] ;
 wire \inst$top.soc.cpu.sink__payload$18[181] ;
 wire \inst$top.soc.cpu.sink__payload$18[182] ;
 wire \inst$top.soc.cpu.sink__payload$18[183] ;
 wire \inst$top.soc.cpu.sink__payload$18[184] ;
 wire \inst$top.soc.cpu.sink__payload$18[185] ;
 wire \inst$top.soc.cpu.sink__payload$18[186] ;
 wire \inst$top.soc.cpu.sink__payload$18[187] ;
 wire \inst$top.soc.cpu.sink__payload$18[188] ;
 wire \inst$top.soc.cpu.sink__payload$18[189] ;
 wire \inst$top.soc.cpu.sink__payload$18[18] ;
 wire \inst$top.soc.cpu.sink__payload$18[190] ;
 wire \inst$top.soc.cpu.sink__payload$18[191] ;
 wire \inst$top.soc.cpu.sink__payload$18[192] ;
 wire \inst$top.soc.cpu.sink__payload$18[193] ;
 wire \inst$top.soc.cpu.sink__payload$18[194] ;
 wire \inst$top.soc.cpu.sink__payload$18[195] ;
 wire \inst$top.soc.cpu.sink__payload$18[196] ;
 wire \inst$top.soc.cpu.sink__payload$18[197] ;
 wire \inst$top.soc.cpu.sink__payload$18[198] ;
 wire \inst$top.soc.cpu.sink__payload$18[199] ;
 wire \inst$top.soc.cpu.sink__payload$18[19] ;
 wire \inst$top.soc.cpu.sink__payload$18[200] ;
 wire \inst$top.soc.cpu.sink__payload$18[201] ;
 wire \inst$top.soc.cpu.sink__payload$18[202] ;
 wire \inst$top.soc.cpu.sink__payload$18[203] ;
 wire \inst$top.soc.cpu.sink__payload$18[204] ;
 wire \inst$top.soc.cpu.sink__payload$18[205] ;
 wire \inst$top.soc.cpu.sink__payload$18[206] ;
 wire \inst$top.soc.cpu.sink__payload$18[207] ;
 wire \inst$top.soc.cpu.sink__payload$18[208] ;
 wire \inst$top.soc.cpu.sink__payload$18[209] ;
 wire \inst$top.soc.cpu.sink__payload$18[20] ;
 wire \inst$top.soc.cpu.sink__payload$18[210] ;
 wire \inst$top.soc.cpu.sink__payload$18[211] ;
 wire \inst$top.soc.cpu.sink__payload$18[21] ;
 wire \inst$top.soc.cpu.sink__payload$18[22] ;
 wire \inst$top.soc.cpu.sink__payload$18[23] ;
 wire \inst$top.soc.cpu.sink__payload$18[24] ;
 wire \inst$top.soc.cpu.sink__payload$18[25] ;
 wire \inst$top.soc.cpu.sink__payload$18[26] ;
 wire \inst$top.soc.cpu.sink__payload$18[27] ;
 wire \inst$top.soc.cpu.sink__payload$18[28] ;
 wire \inst$top.soc.cpu.sink__payload$18[29] ;
 wire \inst$top.soc.cpu.sink__payload$18[2] ;
 wire \inst$top.soc.cpu.sink__payload$18[30] ;
 wire \inst$top.soc.cpu.sink__payload$18[31] ;
 wire \inst$top.soc.cpu.sink__payload$18[32] ;
 wire \inst$top.soc.cpu.sink__payload$18[33] ;
 wire \inst$top.soc.cpu.sink__payload$18[34] ;
 wire \inst$top.soc.cpu.sink__payload$18[35] ;
 wire \inst$top.soc.cpu.sink__payload$18[36] ;
 wire \inst$top.soc.cpu.sink__payload$18[37] ;
 wire \inst$top.soc.cpu.sink__payload$18[38] ;
 wire \inst$top.soc.cpu.sink__payload$18[39] ;
 wire \inst$top.soc.cpu.sink__payload$18[3] ;
 wire \inst$top.soc.cpu.sink__payload$18[47] ;
 wire \inst$top.soc.cpu.sink__payload$18[48] ;
 wire \inst$top.soc.cpu.sink__payload$18[49] ;
 wire \inst$top.soc.cpu.sink__payload$18[4] ;
 wire \inst$top.soc.cpu.sink__payload$18[50] ;
 wire \inst$top.soc.cpu.sink__payload$18[51] ;
 wire \inst$top.soc.cpu.sink__payload$18[52] ;
 wire \inst$top.soc.cpu.sink__payload$18[53] ;
 wire \inst$top.soc.cpu.sink__payload$18[54] ;
 wire \inst$top.soc.cpu.sink__payload$18[55] ;
 wire \inst$top.soc.cpu.sink__payload$18[56] ;
 wire \inst$top.soc.cpu.sink__payload$18[57] ;
 wire \inst$top.soc.cpu.sink__payload$18[58] ;
 wire \inst$top.soc.cpu.sink__payload$18[59] ;
 wire \inst$top.soc.cpu.sink__payload$18[5] ;
 wire \inst$top.soc.cpu.sink__payload$18[60] ;
 wire \inst$top.soc.cpu.sink__payload$18[61] ;
 wire \inst$top.soc.cpu.sink__payload$18[62] ;
 wire \inst$top.soc.cpu.sink__payload$18[63] ;
 wire \inst$top.soc.cpu.sink__payload$18[6] ;
 wire \inst$top.soc.cpu.sink__payload$18[7] ;
 wire \inst$top.soc.cpu.sink__payload$18[8] ;
 wire \inst$top.soc.cpu.sink__payload$18[9] ;
 wire \inst$top.soc.cpu.sink__payload$24[100] ;
 wire \inst$top.soc.cpu.sink__payload$24[101] ;
 wire \inst$top.soc.cpu.sink__payload$24[102] ;
 wire \inst$top.soc.cpu.sink__payload$24[103] ;
 wire \inst$top.soc.cpu.sink__payload$24[104] ;
 wire \inst$top.soc.cpu.sink__payload$24[105] ;
 wire \inst$top.soc.cpu.sink__payload$24[10] ;
 wire \inst$top.soc.cpu.sink__payload$24[11] ;
 wire \inst$top.soc.cpu.sink__payload$24[12] ;
 wire \inst$top.soc.cpu.sink__payload$24[13] ;
 wire \inst$top.soc.cpu.sink__payload$24[14] ;
 wire \inst$top.soc.cpu.sink__payload$24[15] ;
 wire \inst$top.soc.cpu.sink__payload$24[16] ;
 wire \inst$top.soc.cpu.sink__payload$24[17] ;
 wire \inst$top.soc.cpu.sink__payload$24[18] ;
 wire \inst$top.soc.cpu.sink__payload$24[19] ;
 wire \inst$top.soc.cpu.sink__payload$24[20] ;
 wire \inst$top.soc.cpu.sink__payload$24[21] ;
 wire \inst$top.soc.cpu.sink__payload$24[22] ;
 wire \inst$top.soc.cpu.sink__payload$24[23] ;
 wire \inst$top.soc.cpu.sink__payload$24[24] ;
 wire \inst$top.soc.cpu.sink__payload$24[25] ;
 wire \inst$top.soc.cpu.sink__payload$24[26] ;
 wire \inst$top.soc.cpu.sink__payload$24[27] ;
 wire \inst$top.soc.cpu.sink__payload$24[28] ;
 wire \inst$top.soc.cpu.sink__payload$24[29] ;
 wire \inst$top.soc.cpu.sink__payload$24[2] ;
 wire \inst$top.soc.cpu.sink__payload$24[30] ;
 wire \inst$top.soc.cpu.sink__payload$24[31] ;
 wire \inst$top.soc.cpu.sink__payload$24[32] ;
 wire \inst$top.soc.cpu.sink__payload$24[33] ;
 wire \inst$top.soc.cpu.sink__payload$24[34] ;
 wire \inst$top.soc.cpu.sink__payload$24[35] ;
 wire \inst$top.soc.cpu.sink__payload$24[36] ;
 wire \inst$top.soc.cpu.sink__payload$24[38] ;
 wire \inst$top.soc.cpu.sink__payload$24[39] ;
 wire \inst$top.soc.cpu.sink__payload$24[3] ;
 wire \inst$top.soc.cpu.sink__payload$24[40] ;
 wire \inst$top.soc.cpu.sink__payload$24[41] ;
 wire \inst$top.soc.cpu.sink__payload$24[42] ;
 wire \inst$top.soc.cpu.sink__payload$24[43] ;
 wire \inst$top.soc.cpu.sink__payload$24[44] ;
 wire \inst$top.soc.cpu.sink__payload$24[45] ;
 wire \inst$top.soc.cpu.sink__payload$24[46] ;
 wire \inst$top.soc.cpu.sink__payload$24[47] ;
 wire \inst$top.soc.cpu.sink__payload$24[48] ;
 wire \inst$top.soc.cpu.sink__payload$24[49] ;
 wire \inst$top.soc.cpu.sink__payload$24[4] ;
 wire \inst$top.soc.cpu.sink__payload$24[50] ;
 wire \inst$top.soc.cpu.sink__payload$24[51] ;
 wire \inst$top.soc.cpu.sink__payload$24[52] ;
 wire \inst$top.soc.cpu.sink__payload$24[53] ;
 wire \inst$top.soc.cpu.sink__payload$24[54] ;
 wire \inst$top.soc.cpu.sink__payload$24[55] ;
 wire \inst$top.soc.cpu.sink__payload$24[56] ;
 wire \inst$top.soc.cpu.sink__payload$24[57] ;
 wire \inst$top.soc.cpu.sink__payload$24[58] ;
 wire \inst$top.soc.cpu.sink__payload$24[59] ;
 wire \inst$top.soc.cpu.sink__payload$24[5] ;
 wire \inst$top.soc.cpu.sink__payload$24[60] ;
 wire \inst$top.soc.cpu.sink__payload$24[61] ;
 wire \inst$top.soc.cpu.sink__payload$24[62] ;
 wire \inst$top.soc.cpu.sink__payload$24[63] ;
 wire \inst$top.soc.cpu.sink__payload$24[64] ;
 wire \inst$top.soc.cpu.sink__payload$24[65] ;
 wire \inst$top.soc.cpu.sink__payload$24[66] ;
 wire \inst$top.soc.cpu.sink__payload$24[67] ;
 wire \inst$top.soc.cpu.sink__payload$24[68] ;
 wire \inst$top.soc.cpu.sink__payload$24[69] ;
 wire \inst$top.soc.cpu.sink__payload$24[6] ;
 wire \inst$top.soc.cpu.sink__payload$24[70] ;
 wire \inst$top.soc.cpu.sink__payload$24[71] ;
 wire \inst$top.soc.cpu.sink__payload$24[72] ;
 wire \inst$top.soc.cpu.sink__payload$24[74] ;
 wire \inst$top.soc.cpu.sink__payload$24[75] ;
 wire \inst$top.soc.cpu.sink__payload$24[76] ;
 wire \inst$top.soc.cpu.sink__payload$24[77] ;
 wire \inst$top.soc.cpu.sink__payload$24[78] ;
 wire \inst$top.soc.cpu.sink__payload$24[79] ;
 wire \inst$top.soc.cpu.sink__payload$24[7] ;
 wire \inst$top.soc.cpu.sink__payload$24[80] ;
 wire \inst$top.soc.cpu.sink__payload$24[81] ;
 wire \inst$top.soc.cpu.sink__payload$24[82] ;
 wire \inst$top.soc.cpu.sink__payload$24[83] ;
 wire \inst$top.soc.cpu.sink__payload$24[84] ;
 wire \inst$top.soc.cpu.sink__payload$24[85] ;
 wire \inst$top.soc.cpu.sink__payload$24[86] ;
 wire \inst$top.soc.cpu.sink__payload$24[87] ;
 wire \inst$top.soc.cpu.sink__payload$24[88] ;
 wire \inst$top.soc.cpu.sink__payload$24[89] ;
 wire \inst$top.soc.cpu.sink__payload$24[8] ;
 wire \inst$top.soc.cpu.sink__payload$24[90] ;
 wire \inst$top.soc.cpu.sink__payload$24[91] ;
 wire \inst$top.soc.cpu.sink__payload$24[92] ;
 wire \inst$top.soc.cpu.sink__payload$24[93] ;
 wire \inst$top.soc.cpu.sink__payload$24[94] ;
 wire \inst$top.soc.cpu.sink__payload$24[95] ;
 wire \inst$top.soc.cpu.sink__payload$24[96] ;
 wire \inst$top.soc.cpu.sink__payload$24[97] ;
 wire \inst$top.soc.cpu.sink__payload$24[98] ;
 wire \inst$top.soc.cpu.sink__payload$24[99] ;
 wire \inst$top.soc.cpu.sink__payload$24[9] ;
 wire \inst$top.soc.cpu.sink__payload$6[10] ;
 wire \inst$top.soc.cpu.sink__payload$6[11] ;
 wire \inst$top.soc.cpu.sink__payload$6[12] ;
 wire \inst$top.soc.cpu.sink__payload$6[13] ;
 wire \inst$top.soc.cpu.sink__payload$6[14] ;
 wire \inst$top.soc.cpu.sink__payload$6[15] ;
 wire \inst$top.soc.cpu.sink__payload$6[16] ;
 wire \inst$top.soc.cpu.sink__payload$6[17] ;
 wire \inst$top.soc.cpu.sink__payload$6[18] ;
 wire \inst$top.soc.cpu.sink__payload$6[19] ;
 wire \inst$top.soc.cpu.sink__payload$6[20] ;
 wire \inst$top.soc.cpu.sink__payload$6[21] ;
 wire \inst$top.soc.cpu.sink__payload$6[22] ;
 wire \inst$top.soc.cpu.sink__payload$6[23] ;
 wire \inst$top.soc.cpu.sink__payload$6[24] ;
 wire \inst$top.soc.cpu.sink__payload$6[25] ;
 wire \inst$top.soc.cpu.sink__payload$6[26] ;
 wire \inst$top.soc.cpu.sink__payload$6[27] ;
 wire \inst$top.soc.cpu.sink__payload$6[28] ;
 wire \inst$top.soc.cpu.sink__payload$6[29] ;
 wire \inst$top.soc.cpu.sink__payload$6[2] ;
 wire \inst$top.soc.cpu.sink__payload$6[30] ;
 wire \inst$top.soc.cpu.sink__payload$6[31] ;
 wire \inst$top.soc.cpu.sink__payload$6[32] ;
 wire \inst$top.soc.cpu.sink__payload$6[33] ;
 wire \inst$top.soc.cpu.sink__payload$6[34] ;
 wire \inst$top.soc.cpu.sink__payload$6[35] ;
 wire \inst$top.soc.cpu.sink__payload$6[36] ;
 wire \inst$top.soc.cpu.sink__payload$6[37] ;
 wire \inst$top.soc.cpu.sink__payload$6[38] ;
 wire \inst$top.soc.cpu.sink__payload$6[39] ;
 wire \inst$top.soc.cpu.sink__payload$6[3] ;
 wire \inst$top.soc.cpu.sink__payload$6[40] ;
 wire \inst$top.soc.cpu.sink__payload$6[41] ;
 wire \inst$top.soc.cpu.sink__payload$6[42] ;
 wire \inst$top.soc.cpu.sink__payload$6[43] ;
 wire \inst$top.soc.cpu.sink__payload$6[44] ;
 wire \inst$top.soc.cpu.sink__payload$6[45] ;
 wire \inst$top.soc.cpu.sink__payload$6[47] ;
 wire \inst$top.soc.cpu.sink__payload$6[48] ;
 wire \inst$top.soc.cpu.sink__payload$6[49] ;
 wire \inst$top.soc.cpu.sink__payload$6[4] ;
 wire \inst$top.soc.cpu.sink__payload$6[50] ;
 wire \inst$top.soc.cpu.sink__payload$6[51] ;
 wire \inst$top.soc.cpu.sink__payload$6[52] ;
 wire \inst$top.soc.cpu.sink__payload$6[53] ;
 wire \inst$top.soc.cpu.sink__payload$6[54] ;
 wire \inst$top.soc.cpu.sink__payload$6[55] ;
 wire \inst$top.soc.cpu.sink__payload$6[56] ;
 wire \inst$top.soc.cpu.sink__payload$6[57] ;
 wire \inst$top.soc.cpu.sink__payload$6[58] ;
 wire \inst$top.soc.cpu.sink__payload$6[59] ;
 wire \inst$top.soc.cpu.sink__payload$6[5] ;
 wire \inst$top.soc.cpu.sink__payload$6[60] ;
 wire \inst$top.soc.cpu.sink__payload$6[61] ;
 wire \inst$top.soc.cpu.sink__payload$6[62] ;
 wire \inst$top.soc.cpu.sink__payload$6[63] ;
 wire \inst$top.soc.cpu.sink__payload$6[6] ;
 wire \inst$top.soc.cpu.sink__payload$6[7] ;
 wire \inst$top.soc.cpu.sink__payload$6[8] ;
 wire \inst$top.soc.cpu.sink__payload$6[9] ;
 wire \inst$top.soc.cpu.sink__payload[10] ;
 wire \inst$top.soc.cpu.sink__payload[11] ;
 wire \inst$top.soc.cpu.sink__payload[12] ;
 wire \inst$top.soc.cpu.sink__payload[13] ;
 wire \inst$top.soc.cpu.sink__payload[14] ;
 wire \inst$top.soc.cpu.sink__payload[15] ;
 wire \inst$top.soc.cpu.sink__payload[16] ;
 wire \inst$top.soc.cpu.sink__payload[17] ;
 wire \inst$top.soc.cpu.sink__payload[18] ;
 wire \inst$top.soc.cpu.sink__payload[19] ;
 wire \inst$top.soc.cpu.sink__payload[20] ;
 wire \inst$top.soc.cpu.sink__payload[21] ;
 wire \inst$top.soc.cpu.sink__payload[22] ;
 wire \inst$top.soc.cpu.sink__payload[23] ;
 wire \inst$top.soc.cpu.sink__payload[24] ;
 wire \inst$top.soc.cpu.sink__payload[25] ;
 wire \inst$top.soc.cpu.sink__payload[26] ;
 wire \inst$top.soc.cpu.sink__payload[27] ;
 wire \inst$top.soc.cpu.sink__payload[28] ;
 wire \inst$top.soc.cpu.sink__payload[29] ;
 wire \inst$top.soc.cpu.sink__payload[2] ;
 wire \inst$top.soc.cpu.sink__payload[30] ;
 wire \inst$top.soc.cpu.sink__payload[31] ;
 wire \inst$top.soc.cpu.sink__payload[3] ;
 wire \inst$top.soc.cpu.sink__payload[4] ;
 wire \inst$top.soc.cpu.sink__payload[5] ;
 wire \inst$top.soc.cpu.sink__payload[6] ;
 wire \inst$top.soc.cpu.sink__payload[7] ;
 wire \inst$top.soc.cpu.sink__payload[8] ;
 wire \inst$top.soc.cpu.sink__payload[9] ;
 wire \inst$top.soc.cpu.x.source__valid ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__0._storage[0] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__0._storage[1] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__1._storage[0] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__1._storage[1] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__2._storage[0] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__2._storage[1] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__3._storage[0] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__3._storage[1] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__4._storage[0] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__4._storage[1] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__5._storage[0] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__5._storage[1] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__6._storage[0] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__6._storage[1] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__7._storage[0] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__7._storage[1] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__0._storage ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__0.port__w_data ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__1._storage ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__1.port__w_data ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__2._storage ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__2.port__w_data ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__3._storage ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__3.port__w_data ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__4._storage ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__4.port__w_data ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__5._storage ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__5.port__w_data ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__6._storage ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__6.port__w_data ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__7._storage ;
 wire \inst$top.soc.gpio_0._gpio.bridge.Output.pin__7.port__w_data ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb$20 ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb$21 ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[0] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[1] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[2] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[3] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[4] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[5] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[6] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[7] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__r_en ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[0] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[1] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[2] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[3] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[4] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[5] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[6] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[7] ;
 wire \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__r_en ;
 wire \inst$top.soc.gpio_0._gpio.pin_0_i_sync_ff_0 ;
 wire \inst$top.soc.gpio_0._gpio.pin_1_i_sync_ff_0 ;
 wire \inst$top.soc.gpio_0._gpio.pin_2_i_sync_ff_0 ;
 wire \inst$top.soc.gpio_0._gpio.pin_3_i_sync_ff_0 ;
 wire \inst$top.soc.gpio_0._gpio.pin_4_i_sync_ff_0 ;
 wire \inst$top.soc.gpio_0._gpio.pin_5_i_sync_ff_0 ;
 wire \inst$top.soc.gpio_0._gpio.pin_6_i_sync_ff_0 ;
 wire \inst$top.soc.gpio_0._gpio.pin_7_i_sync_ff_0 ;
 wire net653;
 wire net652;
 wire net651;
 wire net650;
 wire net649;
 wire net648;
 wire net647;
 wire net646;
 wire \inst$top.soc.gpio_0._gpio.r_data ;
 wire \inst$top.soc.gpio_0._gpio.r_data$23 ;
 wire \inst$top.soc.gpio_0._gpio.r_data$35 ;
 wire \inst$top.soc.gpio_0._gpio.r_data$47 ;
 wire \inst$top.soc.gpio_0._gpio.r_data$59 ;
 wire \inst$top.soc.gpio_0._gpio.r_data$71 ;
 wire \inst$top.soc.gpio_0._gpio.r_data$83 ;
 wire \inst$top.soc.gpio_0._gpio.r_data$95 ;
 wire \inst$top.soc.gpio_0._gpio.w_data ;
 wire \inst$top.soc.gpio_0._gpio.w_data$16 ;
 wire \inst$top.soc.gpio_0._gpio.w_data$26 ;
 wire \inst$top.soc.gpio_0._gpio.w_data$29 ;
 wire \inst$top.soc.gpio_0._gpio.w_data$38 ;
 wire \inst$top.soc.gpio_0._gpio.w_data$41 ;
 wire \inst$top.soc.gpio_0._gpio.w_data$50 ;
 wire \inst$top.soc.gpio_0._gpio.w_data$53 ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__0._storage[0] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__0._storage[1] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__1._storage[0] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__1._storage[1] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__2._storage[0] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__2._storage[1] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__3._storage[0] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__3._storage[1] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__0._storage ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__0.port__w_data ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__1._storage ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__1.port__w_data ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__2._storage ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__2.port__w_data ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__3._storage ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__3.port__w_data ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$14 ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$15 ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[0] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[1] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[2] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[3] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[4] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[5] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[6] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[7] ;
 wire \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__r_en ;
 wire \inst$top.soc.gpio_open_drain._gpio.pin_0_i_sync_ff_0 ;
 wire \inst$top.soc.gpio_open_drain._gpio.pin_1_i_sync_ff_0 ;
 wire \inst$top.soc.gpio_open_drain._gpio.pin_2_i_sync_ff_0 ;
 wire \inst$top.soc.gpio_open_drain._gpio.pin_3_i_sync_ff_0 ;
 wire net636;
 wire net635;
 wire net634;
 wire net633;
 wire \inst$top.soc.gpio_open_drain._gpio.r_data ;
 wire \inst$top.soc.gpio_open_drain._gpio.r_data$23 ;
 wire \inst$top.soc.gpio_open_drain._gpio.r_data$35 ;
 wire \inst$top.soc.gpio_open_drain._gpio.r_data$47 ;
 wire \inst$top.soc.gpio_open_drain._gpio.w_data$38 ;
 wire \inst$top.soc.gpio_open_drain._gpio.w_data$41 ;
 wire \inst$top.soc.gpio_open_drain._gpio.w_data$50 ;
 wire \inst$top.soc.gpio_open_drain._gpio.w_data$53 ;
 wire \inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[0] ;
 wire \inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[1] ;
 wire \inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[6] ;
 wire \inst$top.soc.soc_id.bridge.mux.r_shadow__0__r_en ;
 wire \inst$top.soc.soc_id.bridge.mux.r_shadow__1__r_en ;
 wire \inst$top.soc.soc_id.bridge.mux.r_shadow__2__r_en ;
 wire \inst$top.soc.soc_id.bridge.mux.r_shadow__3__r_en ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[0] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[1] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.Config.port__w_data ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.Config.raw_enable._storage ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[0] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[1] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.RawControl.port__w_data ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[0] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[1] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[2] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[3] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[4] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[5] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[6] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[7] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12.w_stb ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb$16 ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb$17 ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[0] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[1] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[2] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[3] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[4] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[5] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[6] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[7] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__r_en ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[2] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[3] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[4] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[5] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[6] ;
 wire \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[7] ;
 wire \inst$top.soc.spiflash.ctrl.fsm_state[0] ;
 wire \inst$top.soc.spiflash.ctrl.fsm_state[1] ;
 wire \inst$top.soc.spiflash.ctrl.fsm_state[2] ;
 wire \inst$top.soc.spiflash.ctrl.fsm_state[3] ;
 wire \inst$top.soc.spiflash.ctrl.i_data_count[0] ;
 wire \inst$top.soc.spiflash.ctrl.i_data_count[1] ;
 wire \inst$top.soc.spiflash.ctrl.i_data_count[2] ;
 wire \inst$top.soc.spiflash.ctrl.o_addr_count[0] ;
 wire \inst$top.soc.spiflash.ctrl.o_addr_count[1] ;
 wire \inst$top.soc.spiflash.ctrl.o_data_count[0] ;
 wire \inst$top.soc.spiflash.ctrl.o_data_count[1] ;
 wire \inst$top.soc.spiflash.ctrl.o_data_count[2] ;
 wire \inst$top.soc.spiflash.ctrl.o_dummy_count[0] ;
 wire \inst$top.soc.spiflash.ctrl.o_dummy_count[1] ;
 wire \inst$top.soc.spiflash.ctrl.r_data[0] ;
 wire \inst$top.soc.spiflash.ctrl.r_data[1] ;
 wire \inst$top.soc.spiflash.ctrl.r_data[2] ;
 wire \inst$top.soc.spiflash.ctrl.r_data[3] ;
 wire \inst$top.soc.spiflash.ctrl.r_data[4] ;
 wire \inst$top.soc.spiflash.ctrl.r_data[5] ;
 wire \inst$top.soc.spiflash.ctrl.r_data[6] ;
 wire \inst$top.soc.spiflash.ctrl.r_data[7] ;
 wire \inst$top.soc.spiflash.ctrl.raw_tx_data[0] ;
 wire \inst$top.soc.spiflash.ctrl.raw_tx_data[1] ;
 wire \inst$top.soc.spiflash.ctrl.raw_tx_data[2] ;
 wire \inst$top.soc.spiflash.ctrl.raw_tx_data[3] ;
 wire \inst$top.soc.spiflash.ctrl.raw_tx_data[4] ;
 wire \inst$top.soc.spiflash.ctrl.raw_tx_data[5] ;
 wire \inst$top.soc.spiflash.ctrl.raw_tx_data[6] ;
 wire \inst$top.soc.spiflash.ctrl.raw_tx_data[7] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__ack ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[0] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[10] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[11] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[12] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[13] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[14] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[15] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[16] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[17] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[18] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[19] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[1] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[20] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[21] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[22] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[23] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[24] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[25] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[26] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[27] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[28] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[29] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[2] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[30] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[31] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[3] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[4] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[5] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[6] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[7] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[8] ;
 wire \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[9] ;
 wire \inst$top.soc.spiflash.phy.deframer.cycle[0] ;
 wire \inst$top.soc.spiflash.phy.deframer.cycle[1] ;
 wire \inst$top.soc.spiflash.phy.deframer.cycle[2] ;
 wire \inst$top.soc.spiflash.phy.deframer.data_reg[0] ;
 wire \inst$top.soc.spiflash.phy.deframer.data_reg[1] ;
 wire \inst$top.soc.spiflash.phy.deframer.data_reg[2] ;
 wire \inst$top.soc.spiflash.phy.deframer.data_reg[3] ;
 wire \inst$top.soc.spiflash.phy.deframer.data_reg[4] ;
 wire \inst$top.soc.spiflash.phy.deframer.data_reg[5] ;
 wire \inst$top.soc.spiflash.phy.deframer.data_reg[6] ;
 wire \inst$top.soc.spiflash.phy.enframer.cycle[0] ;
 wire \inst$top.soc.spiflash.phy.enframer.cycle[1] ;
 wire \inst$top.soc.spiflash.phy.enframer.cycle[2] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.fsm_state ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[0] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[10] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[11] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[12] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[13] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[14] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[15] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[1] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[2] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[3] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[4] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[5] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[6] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[7] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[8] ;
 wire \inst$top.soc.spiflash.phy.io_clocker.timer[9] ;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_cs.o ;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_cs.o_ff ;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_io0.i_ff ;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_io0.o ;
 wire net659;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_io0.oe ;
 wire net747;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_io1.i_ff ;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_io1.o ;
 wire net658;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_io1.oe ;
 wire net746;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_io2.i_ff ;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_io2.o ;
 wire net657;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_io2.oe ;
 wire net745;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_io3.i_ff ;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_io3.o ;
 wire net656;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_io3.oe ;
 wire net744;
 wire \inst$top.soc.spiflash.phy.io_streamer.buffer_sck.o ;
 wire net661;
 wire \inst$top.soc.spiflash.phy.io_streamer.i_en_0 ;
 wire \inst$top.soc.spiflash.phy.io_streamer.meta_0[0] ;
 wire \inst$top.soc.spiflash.phy.io_streamer.meta_0[1] ;
 wire \inst$top.soc.spiflash.phy.io_streamer.meta_0[2] ;
 wire \inst$top.soc.spiflash.phy.io_streamer.o_latch.cs.o ;
 wire \inst$top.soc.spiflash.phy.io_streamer.o_latch.io0.o ;
 wire \inst$top.soc.spiflash.phy.io_streamer.o_latch.io0.oe ;
 wire \inst$top.soc.spiflash.phy.io_streamer.o_latch.io1.o ;
 wire \inst$top.soc.spiflash.phy.io_streamer.o_latch.io1.oe ;
 wire \inst$top.soc.spiflash.phy.io_streamer.o_latch.io2.o ;
 wire \inst$top.soc.spiflash.phy.io_streamer.o_latch.io2.oe ;
 wire \inst$top.soc.spiflash.phy.io_streamer.o_latch.io3.o ;
 wire \inst$top.soc.spiflash.phy.io_streamer.o_latch.io3.oe ;
 wire \inst$top.soc.spiflash.phy.io_streamer.o_latch.sck.o ;
 wire \inst$top.soc.spiflash.phy.io_streamer.skid_1.meta[0] ;
 wire \inst$top.soc.spiflash.phy.io_streamer.skid_1.meta[1] ;
 wire \inst$top.soc.spiflash.phy.io_streamer.skid_1.meta[2] ;
 wire \inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io0 ;
 wire \inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io1 ;
 wire \inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io2 ;
 wire \inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io3 ;
 wire \inst$top.soc.spiflash.phy.io_streamer.skid_at ;
 wire \inst$top.soc.sram.read_port__data[0] ;
 wire \inst$top.soc.sram.read_port__data[10] ;
 wire \inst$top.soc.sram.read_port__data[11] ;
 wire \inst$top.soc.sram.read_port__data[12] ;
 wire \inst$top.soc.sram.read_port__data[13] ;
 wire \inst$top.soc.sram.read_port__data[14] ;
 wire \inst$top.soc.sram.read_port__data[15] ;
 wire \inst$top.soc.sram.read_port__data[16] ;
 wire \inst$top.soc.sram.read_port__data[17] ;
 wire \inst$top.soc.sram.read_port__data[18] ;
 wire \inst$top.soc.sram.read_port__data[19] ;
 wire \inst$top.soc.sram.read_port__data[1] ;
 wire \inst$top.soc.sram.read_port__data[20] ;
 wire \inst$top.soc.sram.read_port__data[21] ;
 wire \inst$top.soc.sram.read_port__data[22] ;
 wire \inst$top.soc.sram.read_port__data[23] ;
 wire \inst$top.soc.sram.read_port__data[24] ;
 wire \inst$top.soc.sram.read_port__data[25] ;
 wire \inst$top.soc.sram.read_port__data[26] ;
 wire \inst$top.soc.sram.read_port__data[27] ;
 wire \inst$top.soc.sram.read_port__data[28] ;
 wire \inst$top.soc.sram.read_port__data[29] ;
 wire \inst$top.soc.sram.read_port__data[2] ;
 wire \inst$top.soc.sram.read_port__data[30] ;
 wire \inst$top.soc.sram.read_port__data[31] ;
 wire \inst$top.soc.sram.read_port__data[3] ;
 wire \inst$top.soc.sram.read_port__data[4] ;
 wire \inst$top.soc.sram.read_port__data[5] ;
 wire \inst$top.soc.sram.read_port__data[6] ;
 wire \inst$top.soc.sram.read_port__data[7] ;
 wire \inst$top.soc.sram.read_port__data[8] ;
 wire \inst$top.soc.sram.read_port__data[9] ;
 wire \inst$top.soc.sram.read_port__en ;
 wire \inst$top.soc.sram.wb_bus__ack ;
 wire \inst$top.soc.sram.write_port__en[0] ;
 wire \inst$top.soc.sram.write_port__en[1] ;
 wire \inst$top.soc.sram.write_port__en[2] ;
 wire \inst$top.soc.sram.write_port__en[3] ;
 wire \inst$top.soc.uart_0._phy.rx.err.frame ;
 wire \inst$top.soc.uart_0._phy.rx.lower.bitno[0] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.bitno[1] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.bitno[2] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.bitno[3] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.data[0] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.data[1] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.data[2] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.data[3] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.data[4] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.data[5] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.data[6] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.data[7] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.fsm_state[0] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.fsm_state[1] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.rdy ;
 wire \inst$top.soc.uart_0._phy.rx.lower.shreg.start ;
 wire \inst$top.soc.uart_0._phy.rx.lower.shreg.stop ;
 wire \inst$top.soc.uart_0._phy.rx.lower.shreg[1] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.shreg[2] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.shreg[3] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.shreg[4] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.shreg[5] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.shreg[6] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.shreg[7] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.shreg[8] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[0] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[10] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[11] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[12] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[13] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[14] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[15] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[16] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[17] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[18] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[19] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[1] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[20] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[21] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[22] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[23] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[2] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[3] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[4] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[5] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[6] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[7] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[8] ;
 wire \inst$top.soc.uart_0._phy.rx.lower.timer[9] ;
 wire \inst$top.soc.uart_0._phy.rx.overflow ;
 wire \inst$top.soc.uart_0._phy.rx.symbols__payload[0] ;
 wire \inst$top.soc.uart_0._phy.rx.symbols__payload[1] ;
 wire \inst$top.soc.uart_0._phy.rx.symbols__payload[2] ;
 wire \inst$top.soc.uart_0._phy.rx.symbols__payload[3] ;
 wire \inst$top.soc.uart_0._phy.rx.symbols__payload[4] ;
 wire \inst$top.soc.uart_0._phy.rx.symbols__payload[5] ;
 wire \inst$top.soc.uart_0._phy.rx.symbols__payload[6] ;
 wire \inst$top.soc.uart_0._phy.rx.symbols__payload[7] ;
 wire \inst$top.soc.uart_0._phy.rx.symbols__valid ;
 wire \inst$top.soc.uart_0._phy.tx.lower.bitno[0] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.bitno[1] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.bitno[2] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.bitno[3] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.fsm_state ;
 wire net655;
 wire \inst$top.soc.uart_0._phy.tx.lower.shreg.start ;
 wire \inst$top.soc.uart_0._phy.tx.lower.shreg.stop ;
 wire \inst$top.soc.uart_0._phy.tx.lower.shreg[1] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.shreg[2] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.shreg[3] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.shreg[4] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.shreg[5] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.shreg[6] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.shreg[7] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.shreg[8] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[0] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[10] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[11] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[12] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[13] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[14] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[15] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[16] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[17] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[18] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[19] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[1] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[20] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[21] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[22] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[23] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[2] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[3] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[4] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[5] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[6] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[7] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[8] ;
 wire \inst$top.soc.uart_0._phy.tx.lower.timer[9] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.Config.enable._storage ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.Config.enable.port__w_data ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[0] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[10] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[11] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[12] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[13] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[14] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[15] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[16] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[17] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[18] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[19] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[1] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[20] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[21] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[22] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[23] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[2] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[3] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[4] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[5] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[6] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[7] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[8] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[9] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.Status.error._storage ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.Status.error.port__w_data ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.Status.overflow._storage ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.Status.overflow.port__w_data ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb$25 ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb$34 ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[0] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[1] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[2] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[3] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[4] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[5] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[6] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[7] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__r_en ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[0] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[1] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[2] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[3] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[4] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[5] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[6] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[7] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__r_en ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[0] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[1] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[2] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[3] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[4] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[5] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[6] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[7] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__r_en ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[3] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[4] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[5] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[6] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[7] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[0] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[1] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[2] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[3] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[4] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[5] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[6] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[7] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[0] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[1] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[2] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[3] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[4] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[5] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[6] ;
 wire \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[7] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.Config.enable._storage ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.Config.enable.port__w_data ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[0] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[10] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[11] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[12] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[13] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[14] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[15] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[16] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[17] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[18] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[19] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[1] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[20] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[21] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[22] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[23] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[2] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[3] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[4] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[5] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[6] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[7] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[8] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[9] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb$27 ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb$32 ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[0] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[1] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[2] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[3] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[4] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[5] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[6] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[7] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__r_en ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[0] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[1] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[2] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[3] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[4] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[5] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[6] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[7] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__r_en ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[0] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[1] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[2] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[3] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[4] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[5] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[6] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[7] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__r_en ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[1] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[2] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[3] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[4] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[5] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[6] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[7] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[0] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[1] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[2] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[3] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[4] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[5] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[6] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[7] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[0] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[1] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[2] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[3] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[4] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[5] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[6] ;
 wire \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[7] ;
 wire \inst$top.soc.wb_arbiter.grant ;
 wire \inst$top.soc.wb_to_csr.cycle[0] ;
 wire \inst$top.soc.wb_to_csr.cycle[1] ;
 wire \inst$top.soc.wb_to_csr.cycle[2] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__ack ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[0] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[10] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[11] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[12] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[13] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[14] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[15] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[16] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[17] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[18] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[19] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[1] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[20] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[21] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[22] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[23] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[24] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[25] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[26] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[27] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[28] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[29] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[2] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[30] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[31] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[3] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[4] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[5] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[6] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[7] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[8] ;
 wire \inst$top.soc.wb_to_csr.wb_bus__dat_r[9] ;
 wire net1101;
 wire net1100;
 wire net1099;
 wire net1098;
 wire net1097;
 wire net1096;
 wire net1095;
 wire net1094;
 wire net1093;
 wire net1092;
 wire net1091;
 wire net1090;
 wire net1089;
 wire net1088;
 wire net1087;
 wire net1086;
 wire net1085;
 wire net1084;
 wire net1083;
 wire net1082;
 wire net1081;
 wire net1080;
 wire net1079;
 wire net1078;
 wire net1077;
 wire net1076;
 wire net1075;
 wire net1074;
 wire net1073;
 wire net1072;
 wire net1071;
 wire net1070;
 wire net1069;
 wire net1068;
 wire net1067;
 wire net1066;
 wire net1065;
 wire net1064;
 wire net1063;
 wire net1062;
 wire net1061;
 wire net1060;
 wire net1059;
 wire net1058;
 wire net1057;
 wire net1056;
 wire net1055;
 wire net1054;
 wire net1053;
 wire net1052;
 wire net1051;
 wire net1050;
 wire net1049;
 wire net1048;
 wire net1047;
 wire net1046;
 wire net1045;
 wire net1044;
 wire net1043;
 wire net1042;
 wire net1041;
 wire net1040;
 wire net1039;
 wire net1038;
 wire net1037;
 wire net1036;
 wire net1035;
 wire net1034;
 wire net1033;
 wire net1032;
 wire net1031;
 wire net1030;
 wire net1029;
 wire net1028;
 wire net1027;
 wire net1026;
 wire net1025;
 wire net1024;
 wire net1023;
 wire net1022;
 wire net1021;
 wire net1020;
 wire net1019;
 wire net1018;
 wire net1017;
 wire net1016;
 wire net1015;
 wire net1014;
 wire net1013;
 wire net1012;
 wire net1011;
 wire net1010;
 wire net1009;
 wire net1008;
 wire net1007;
 wire net1006;
 wire net1005;
 wire net1004;
 wire net1003;
 wire net1002;
 wire net1001;
 wire net1000;
 wire net999;
 wire net998;
 wire net997;
 wire net996;
 wire net995;
 wire net994;
 wire net993;
 wire net992;
 wire net991;
 wire net990;
 wire net989;
 wire net988;
 wire net987;
 wire net986;
 wire net985;
 wire net984;
 wire net983;
 wire net982;
 wire net981;
 wire net980;
 wire net979;
 wire net978;
 wire net977;
 wire net976;
 wire net975;
 wire net974;
 wire net973;
 wire net972;
 wire net971;
 wire net970;
 wire net962;
 wire net953;
 wire net952;
 wire net951;
 wire net950;
 wire net949;
 wire net948;
 wire net947;
 wire net946;
 wire net945;
 wire net940;
 wire net939;
 wire net938;
 wire net937;
 wire net936;
 wire net935;
 wire net934;
 wire net933;
 wire net932;
 wire net931;
 wire net930;
 wire net929;
 wire net928;
 wire net927;
 wire net926;
 wire net918;
 wire net909;
 wire net908;
 wire net907;
 wire net906;
 wire net905;
 wire net904;
 wire net903;
 wire net902;
 wire net901;
 wire net896;
 wire net895;
 wire net894;
 wire net893;
 wire net892;
 wire net891;
 wire net890;
 wire net889;
 wire net888;
 wire net887;
 wire net886;
 wire net885;
 wire net884;
 wire net883;
 wire net882;
 wire net881;
 wire net880;
 wire net879;
 wire net878;
 wire net877;
 wire net876;
 wire net875;
 wire net874;
 wire net873;
 wire net872;
 wire net871;
 wire net870;
 wire net869;
 wire net868;
 wire net867;
 wire net866;
 wire net865;
 wire net864;
 wire net863;
 wire net862;
 wire net861;
 wire net860;
 wire net859;
 wire net858;
 wire net857;
 wire net856;
 wire net855;
 wire net854;
 wire net853;
 wire net852;
 wire net851;
 wire net850;
 wire net849;
 wire net848;
 wire net847;
 wire net846;
 wire net845;
 wire net844;
 wire net843;
 wire net842;
 wire net841;
 wire net840;
 wire net839;
 wire net838;
 wire net837;
 wire net836;
 wire net835;
 wire net834;
 wire net833;
 wire net832;
 wire net831;
 wire net830;
 wire net829;
 wire net828;
 wire net827;
 wire net826;
 wire net825;
 wire net824;
 wire net823;
 wire net822;
 wire net821;
 wire net820;
 wire net819;
 wire net818;
 wire net817;
 wire net816;
 wire net815;
 wire net814;
 wire net813;
 wire net812;
 wire net811;
 wire net810;
 wire net809;
 wire net808;
 wire net807;
 wire net806;
 wire net805;
 wire net804;
 wire net803;
 wire net802;
 wire net801;
 wire net800;
 wire net799;
 wire net798;
 wire net797;
 wire net796;
 wire net795;
 wire net794;
 wire net793;
 wire net792;
 wire net791;
 wire net790;
 wire net789;
 wire net788;
 wire net787;
 wire net786;
 wire net785;
 wire net784;
 wire net783;
 wire net782;
 wire net781;
 wire net780;
 wire net779;
 wire net778;
 wire net777;
 wire net776;
 wire net775;
 wire net774;
 wire net773;
 wire net772;
 wire net771;
 wire net770;
 wire net769;
 wire net768;
 wire net767;
 wire net766;
 wire net765;
 wire net764;
 wire net763;
 wire net762;
 wire net761;
 wire net760;
 wire net759;
 wire net758;
 wire net757;
 wire net756;
 wire net755;
 wire net754;
 wire net753;
 wire net752;
 wire net751;
 wire net750;
 wire net742;
 wire net711;
 wire net709;
 wire net705;
 wire net704;
 wire net699;
 wire net654;
 wire net645;
 wire net644;
 wire net643;
 wire net642;
 wire net641;
 wire net640;
 wire net639;
 wire net638;
 wire net637;
 wire net632;
 wire net631;
 wire net630;
 wire net629;
 wire net628;
 wire net627;
 wire net626;
 wire net625;
 wire net624;
 wire net623;
 wire net622;
 wire net621;
 wire net620;
 wire net619;
 wire net618;
 wire net617;
 wire net616;
 wire net615;
 wire net614;
 wire net613;
 wire net612;
 wire net611;
 wire net610;
 wire net609;
 wire net608;
 wire net607;
 wire net606;
 wire net605;
 wire net604;
 wire net603;
 wire net602;
 wire net601;
 wire net549;
 wire net548;
 wire net547;
 wire net546;
 wire net545;
 wire net544;
 wire net543;
 wire net542;
 wire net541;
 wire net540;
 wire net539;
 wire net538;
 wire net537;
 wire net536;
 wire net535;
 wire net534;
 wire net533;
 wire net532;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net968;
 wire net967;
 wire net966;
 wire net965;
 wire net964;
 wire net963;
 wire net961;
 wire net960;
 wire net959;
 wire net958;
 wire net957;
 wire net956;
 wire net955;
 wire net954;
 wire net944;
 wire net943;
 wire net942;
 wire net941;
 wire net925;
 wire net924;
 wire net923;
 wire net922;
 wire net921;
 wire net920;
 wire net919;
 wire net917;
 wire net916;
 wire net915;
 wire net914;
 wire net913;
 wire net912;
 wire net911;
 wire net910;
 wire net900;
 wire net899;
 wire net898;
 wire net897;
 wire net749;
 wire net748;
 wire net743;
 wire net733;
 wire net732;
 wire net731;
 wire net730;
 wire net729;
 wire net728;
 wire net727;
 wire net726;
 wire net725;
 wire net720;
 wire net719;
 wire net718;
 wire net717;
 wire net716;
 wire net715;
 wire net714;
 wire net713;
 wire net712;
 wire net710;
 wire net708;
 wire net707;
 wire net706;
 wire net698;
 wire net689;
 wire net688;
 wire net687;
 wire net686;
 wire net685;
 wire net684;
 wire net683;
 wire net682;
 wire net681;
 wire net676;
 wire net675;
 wire net674;
 wire net673;
 wire net672;
 wire net671;
 wire net670;
 wire net669;
 wire net668;
 wire net667;
 wire net666;
 wire net665;
 wire net664;
 wire net663;
 wire net662;
 wire net529;
 wire net530;
 wire net531;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire clk_in_regs;
 wire clknet_0_clk_in;
 wire clknet_1_0__leaf_clk_in;
 wire clknet_leaf_0_clk_in_regs;
 wire clknet_leaf_1_clk_in_regs;
 wire clknet_leaf_2_clk_in_regs;
 wire clknet_leaf_4_clk_in_regs;
 wire clknet_leaf_5_clk_in_regs;
 wire clknet_leaf_6_clk_in_regs;
 wire clknet_leaf_8_clk_in_regs;
 wire clknet_leaf_9_clk_in_regs;
 wire clknet_leaf_10_clk_in_regs;
 wire clknet_leaf_11_clk_in_regs;
 wire clknet_leaf_12_clk_in_regs;
 wire clknet_leaf_13_clk_in_regs;
 wire clknet_leaf_14_clk_in_regs;
 wire clknet_leaf_15_clk_in_regs;
 wire clknet_leaf_16_clk_in_regs;
 wire clknet_leaf_17_clk_in_regs;
 wire clknet_leaf_18_clk_in_regs;
 wire clknet_leaf_19_clk_in_regs;
 wire clknet_leaf_21_clk_in_regs;
 wire clknet_leaf_22_clk_in_regs;
 wire clknet_leaf_23_clk_in_regs;
 wire clknet_leaf_24_clk_in_regs;
 wire clknet_leaf_25_clk_in_regs;
 wire clknet_leaf_26_clk_in_regs;
 wire clknet_leaf_27_clk_in_regs;
 wire clknet_leaf_28_clk_in_regs;
 wire clknet_leaf_29_clk_in_regs;
 wire clknet_leaf_30_clk_in_regs;
 wire clknet_leaf_31_clk_in_regs;
 wire clknet_leaf_32_clk_in_regs;
 wire clknet_leaf_33_clk_in_regs;
 wire clknet_leaf_34_clk_in_regs;
 wire clknet_leaf_35_clk_in_regs;
 wire clknet_leaf_36_clk_in_regs;
 wire clknet_leaf_37_clk_in_regs;
 wire clknet_leaf_38_clk_in_regs;
 wire clknet_leaf_39_clk_in_regs;
 wire clknet_leaf_40_clk_in_regs;
 wire clknet_leaf_41_clk_in_regs;
 wire clknet_leaf_42_clk_in_regs;
 wire clknet_leaf_43_clk_in_regs;
 wire clknet_leaf_44_clk_in_regs;
 wire clknet_leaf_45_clk_in_regs;
 wire clknet_leaf_46_clk_in_regs;
 wire clknet_leaf_47_clk_in_regs;
 wire clknet_leaf_48_clk_in_regs;
 wire clknet_leaf_49_clk_in_regs;
 wire clknet_leaf_50_clk_in_regs;
 wire clknet_leaf_51_clk_in_regs;
 wire clknet_leaf_52_clk_in_regs;
 wire clknet_leaf_53_clk_in_regs;
 wire clknet_leaf_54_clk_in_regs;
 wire clknet_leaf_55_clk_in_regs;
 wire clknet_leaf_56_clk_in_regs;
 wire clknet_leaf_57_clk_in_regs;
 wire clknet_leaf_58_clk_in_regs;
 wire clknet_leaf_59_clk_in_regs;
 wire clknet_leaf_60_clk_in_regs;
 wire clknet_leaf_61_clk_in_regs;
 wire clknet_leaf_62_clk_in_regs;
 wire clknet_leaf_63_clk_in_regs;
 wire clknet_leaf_64_clk_in_regs;
 wire clknet_leaf_65_clk_in_regs;
 wire clknet_leaf_66_clk_in_regs;
 wire clknet_leaf_67_clk_in_regs;
 wire clknet_leaf_68_clk_in_regs;
 wire clknet_leaf_69_clk_in_regs;
 wire clknet_leaf_70_clk_in_regs;
 wire clknet_leaf_71_clk_in_regs;
 wire clknet_leaf_72_clk_in_regs;
 wire clknet_leaf_73_clk_in_regs;
 wire clknet_leaf_74_clk_in_regs;
 wire clknet_leaf_75_clk_in_regs;
 wire clknet_leaf_76_clk_in_regs;
 wire clknet_leaf_77_clk_in_regs;
 wire clknet_leaf_78_clk_in_regs;
 wire clknet_leaf_79_clk_in_regs;
 wire clknet_leaf_80_clk_in_regs;
 wire clknet_leaf_81_clk_in_regs;
 wire clknet_leaf_82_clk_in_regs;
 wire clknet_leaf_83_clk_in_regs;
 wire clknet_leaf_84_clk_in_regs;
 wire clknet_leaf_85_clk_in_regs;
 wire clknet_leaf_86_clk_in_regs;
 wire clknet_leaf_87_clk_in_regs;
 wire clknet_leaf_89_clk_in_regs;
 wire clknet_leaf_90_clk_in_regs;
 wire clknet_leaf_91_clk_in_regs;
 wire clknet_leaf_92_clk_in_regs;
 wire clknet_leaf_93_clk_in_regs;
 wire clknet_leaf_94_clk_in_regs;
 wire clknet_leaf_95_clk_in_regs;
 wire clknet_leaf_96_clk_in_regs;
 wire clknet_leaf_97_clk_in_regs;
 wire clknet_leaf_98_clk_in_regs;
 wire clknet_leaf_99_clk_in_regs;
 wire clknet_leaf_100_clk_in_regs;
 wire clknet_leaf_102_clk_in_regs;
 wire clknet_leaf_103_clk_in_regs;
 wire clknet_leaf_104_clk_in_regs;
 wire clknet_leaf_105_clk_in_regs;
 wire clknet_leaf_106_clk_in_regs;
 wire clknet_leaf_107_clk_in_regs;
 wire clknet_leaf_108_clk_in_regs;
 wire clknet_leaf_109_clk_in_regs;
 wire clknet_leaf_110_clk_in_regs;
 wire clknet_leaf_111_clk_in_regs;
 wire clknet_leaf_113_clk_in_regs;
 wire clknet_leaf_114_clk_in_regs;
 wire clknet_leaf_115_clk_in_regs;
 wire clknet_leaf_116_clk_in_regs;
 wire clknet_leaf_117_clk_in_regs;
 wire clknet_leaf_118_clk_in_regs;
 wire clknet_leaf_119_clk_in_regs;
 wire clknet_leaf_121_clk_in_regs;
 wire clknet_leaf_123_clk_in_regs;
 wire clknet_leaf_124_clk_in_regs;
 wire clknet_leaf_127_clk_in_regs;
 wire clknet_leaf_128_clk_in_regs;
 wire clknet_leaf_129_clk_in_regs;
 wire clknet_leaf_130_clk_in_regs;
 wire clknet_leaf_131_clk_in_regs;
 wire clknet_leaf_132_clk_in_regs;
 wire clknet_leaf_134_clk_in_regs;
 wire clknet_leaf_135_clk_in_regs;
 wire clknet_leaf_138_clk_in_regs;
 wire clknet_leaf_140_clk_in_regs;
 wire clknet_leaf_143_clk_in_regs;
 wire clknet_leaf_144_clk_in_regs;
 wire clknet_leaf_145_clk_in_regs;
 wire clknet_leaf_146_clk_in_regs;
 wire clknet_leaf_147_clk_in_regs;
 wire clknet_leaf_148_clk_in_regs;
 wire clknet_leaf_149_clk_in_regs;
 wire clknet_leaf_150_clk_in_regs;
 wire clknet_leaf_151_clk_in_regs;
 wire clknet_leaf_152_clk_in_regs;
 wire clknet_leaf_153_clk_in_regs;
 wire clknet_leaf_154_clk_in_regs;
 wire clknet_leaf_155_clk_in_regs;
 wire clknet_leaf_156_clk_in_regs;
 wire clknet_leaf_157_clk_in_regs;
 wire clknet_leaf_158_clk_in_regs;
 wire clknet_leaf_159_clk_in_regs;
 wire clknet_leaf_160_clk_in_regs;
 wire clknet_leaf_161_clk_in_regs;
 wire clknet_leaf_162_clk_in_regs;
 wire clknet_leaf_163_clk_in_regs;
 wire clknet_leaf_164_clk_in_regs;
 wire clknet_leaf_165_clk_in_regs;
 wire clknet_leaf_166_clk_in_regs;
 wire clknet_leaf_167_clk_in_regs;
 wire clknet_leaf_168_clk_in_regs;
 wire clknet_leaf_169_clk_in_regs;
 wire clknet_leaf_170_clk_in_regs;
 wire clknet_leaf_171_clk_in_regs;
 wire clknet_leaf_172_clk_in_regs;
 wire clknet_leaf_173_clk_in_regs;
 wire clknet_leaf_174_clk_in_regs;
 wire clknet_leaf_175_clk_in_regs;
 wire clknet_leaf_176_clk_in_regs;
 wire clknet_leaf_177_clk_in_regs;
 wire clknet_leaf_178_clk_in_regs;
 wire clknet_leaf_179_clk_in_regs;
 wire clknet_leaf_180_clk_in_regs;
 wire clknet_leaf_181_clk_in_regs;
 wire clknet_leaf_182_clk_in_regs;
 wire clknet_leaf_183_clk_in_regs;
 wire clknet_leaf_184_clk_in_regs;
 wire clknet_leaf_185_clk_in_regs;
 wire clknet_leaf_186_clk_in_regs;
 wire clknet_leaf_187_clk_in_regs;
 wire clknet_leaf_188_clk_in_regs;
 wire clknet_leaf_189_clk_in_regs;
 wire clknet_leaf_190_clk_in_regs;
 wire clknet_leaf_191_clk_in_regs;
 wire clknet_leaf_192_clk_in_regs;
 wire clknet_leaf_193_clk_in_regs;
 wire clknet_leaf_194_clk_in_regs;
 wire clknet_leaf_195_clk_in_regs;
 wire clknet_leaf_196_clk_in_regs;
 wire clknet_leaf_197_clk_in_regs;
 wire clknet_leaf_198_clk_in_regs;
 wire clknet_leaf_199_clk_in_regs;
 wire clknet_leaf_200_clk_in_regs;
 wire clknet_leaf_201_clk_in_regs;
 wire clknet_leaf_202_clk_in_regs;
 wire clknet_leaf_203_clk_in_regs;
 wire clknet_leaf_204_clk_in_regs;
 wire clknet_leaf_205_clk_in_regs;
 wire clknet_leaf_206_clk_in_regs;
 wire clknet_leaf_207_clk_in_regs;
 wire clknet_leaf_208_clk_in_regs;
 wire clknet_leaf_209_clk_in_regs;
 wire clknet_leaf_210_clk_in_regs;
 wire clknet_leaf_211_clk_in_regs;
 wire clknet_leaf_212_clk_in_regs;
 wire clknet_leaf_213_clk_in_regs;
 wire clknet_leaf_214_clk_in_regs;
 wire clknet_leaf_215_clk_in_regs;
 wire clknet_leaf_216_clk_in_regs;
 wire clknet_leaf_217_clk_in_regs;
 wire clknet_leaf_218_clk_in_regs;
 wire clknet_leaf_219_clk_in_regs;
 wire clknet_leaf_220_clk_in_regs;
 wire clknet_leaf_221_clk_in_regs;
 wire clknet_leaf_222_clk_in_regs;
 wire clknet_leaf_223_clk_in_regs;
 wire clknet_leaf_224_clk_in_regs;
 wire clknet_leaf_225_clk_in_regs;
 wire clknet_leaf_226_clk_in_regs;
 wire clknet_leaf_227_clk_in_regs;
 wire clknet_leaf_228_clk_in_regs;
 wire clknet_leaf_229_clk_in_regs;
 wire clknet_leaf_231_clk_in_regs;
 wire clknet_leaf_232_clk_in_regs;
 wire clknet_leaf_233_clk_in_regs;
 wire clknet_leaf_236_clk_in_regs;
 wire clknet_leaf_237_clk_in_regs;
 wire clknet_leaf_238_clk_in_regs;
 wire clknet_leaf_239_clk_in_regs;
 wire clknet_leaf_240_clk_in_regs;
 wire clknet_leaf_241_clk_in_regs;
 wire clknet_leaf_242_clk_in_regs;
 wire clknet_leaf_243_clk_in_regs;
 wire clknet_leaf_244_clk_in_regs;
 wire clknet_leaf_245_clk_in_regs;
 wire clknet_leaf_246_clk_in_regs;
 wire clknet_leaf_247_clk_in_regs;
 wire clknet_leaf_248_clk_in_regs;
 wire clknet_leaf_249_clk_in_regs;
 wire clknet_leaf_250_clk_in_regs;
 wire clknet_leaf_251_clk_in_regs;
 wire clknet_leaf_252_clk_in_regs;
 wire clknet_leaf_253_clk_in_regs;
 wire clknet_leaf_254_clk_in_regs;
 wire clknet_leaf_255_clk_in_regs;
 wire clknet_leaf_256_clk_in_regs;
 wire clknet_leaf_257_clk_in_regs;
 wire clknet_leaf_258_clk_in_regs;
 wire clknet_leaf_259_clk_in_regs;
 wire clknet_leaf_260_clk_in_regs;
 wire clknet_leaf_261_clk_in_regs;
 wire clknet_leaf_262_clk_in_regs;
 wire clknet_leaf_263_clk_in_regs;
 wire clknet_leaf_264_clk_in_regs;
 wire clknet_leaf_265_clk_in_regs;
 wire clknet_leaf_266_clk_in_regs;
 wire clknet_leaf_267_clk_in_regs;
 wire clknet_leaf_268_clk_in_regs;
 wire clknet_leaf_269_clk_in_regs;
 wire clknet_leaf_270_clk_in_regs;
 wire clknet_leaf_271_clk_in_regs;
 wire clknet_leaf_272_clk_in_regs;
 wire clknet_leaf_273_clk_in_regs;
 wire clknet_leaf_274_clk_in_regs;
 wire clknet_leaf_275_clk_in_regs;
 wire clknet_leaf_276_clk_in_regs;
 wire clknet_leaf_277_clk_in_regs;
 wire clknet_leaf_278_clk_in_regs;
 wire clknet_leaf_279_clk_in_regs;
 wire clknet_leaf_280_clk_in_regs;
 wire clknet_leaf_281_clk_in_regs;
 wire clknet_leaf_282_clk_in_regs;
 wire clknet_leaf_283_clk_in_regs;
 wire clknet_leaf_284_clk_in_regs;
 wire clknet_leaf_285_clk_in_regs;
 wire clknet_leaf_286_clk_in_regs;
 wire clknet_leaf_287_clk_in_regs;
 wire clknet_leaf_288_clk_in_regs;
 wire clknet_leaf_289_clk_in_regs;
 wire clknet_leaf_290_clk_in_regs;
 wire clknet_leaf_291_clk_in_regs;
 wire clknet_leaf_292_clk_in_regs;
 wire clknet_leaf_293_clk_in_regs;
 wire clknet_leaf_294_clk_in_regs;
 wire clknet_leaf_295_clk_in_regs;
 wire clknet_leaf_296_clk_in_regs;
 wire clknet_leaf_297_clk_in_regs;
 wire clknet_leaf_298_clk_in_regs;
 wire clknet_leaf_299_clk_in_regs;
 wire clknet_leaf_300_clk_in_regs;
 wire clknet_leaf_302_clk_in_regs;
 wire clknet_leaf_303_clk_in_regs;
 wire clknet_leaf_304_clk_in_regs;
 wire clknet_leaf_305_clk_in_regs;
 wire clknet_leaf_308_clk_in_regs;
 wire clknet_leaf_309_clk_in_regs;
 wire clknet_leaf_310_clk_in_regs;
 wire clknet_leaf_311_clk_in_regs;
 wire clknet_leaf_312_clk_in_regs;
 wire clknet_leaf_313_clk_in_regs;
 wire clknet_leaf_314_clk_in_regs;
 wire clknet_leaf_315_clk_in_regs;
 wire clknet_leaf_316_clk_in_regs;
 wire clknet_leaf_317_clk_in_regs;
 wire clknet_leaf_318_clk_in_regs;
 wire clknet_leaf_319_clk_in_regs;
 wire clknet_leaf_320_clk_in_regs;
 wire clknet_leaf_321_clk_in_regs;
 wire clknet_leaf_322_clk_in_regs;
 wire clknet_leaf_323_clk_in_regs;
 wire clknet_leaf_324_clk_in_regs;
 wire clknet_leaf_325_clk_in_regs;
 wire clknet_leaf_327_clk_in_regs;
 wire clknet_leaf_328_clk_in_regs;
 wire clknet_leaf_329_clk_in_regs;
 wire clknet_leaf_330_clk_in_regs;
 wire clknet_leaf_331_clk_in_regs;
 wire clknet_leaf_332_clk_in_regs;
 wire clknet_leaf_333_clk_in_regs;
 wire clknet_leaf_334_clk_in_regs;
 wire clknet_leaf_335_clk_in_regs;
 wire clknet_leaf_337_clk_in_regs;
 wire clknet_leaf_338_clk_in_regs;
 wire clknet_leaf_339_clk_in_regs;
 wire clknet_leaf_340_clk_in_regs;
 wire clknet_leaf_341_clk_in_regs;
 wire clknet_leaf_342_clk_in_regs;
 wire clknet_leaf_343_clk_in_regs;
 wire clknet_leaf_344_clk_in_regs;
 wire clknet_leaf_345_clk_in_regs;
 wire clknet_leaf_346_clk_in_regs;
 wire clknet_leaf_347_clk_in_regs;
 wire clknet_leaf_348_clk_in_regs;
 wire clknet_leaf_349_clk_in_regs;
 wire clknet_leaf_350_clk_in_regs;
 wire clknet_leaf_351_clk_in_regs;
 wire clknet_leaf_352_clk_in_regs;
 wire clknet_leaf_353_clk_in_regs;
 wire clknet_leaf_354_clk_in_regs;
 wire clknet_leaf_355_clk_in_regs;
 wire clknet_leaf_356_clk_in_regs;
 wire clknet_leaf_357_clk_in_regs;
 wire clknet_leaf_358_clk_in_regs;
 wire clknet_leaf_359_clk_in_regs;
 wire clknet_leaf_360_clk_in_regs;
 wire clknet_leaf_361_clk_in_regs;
 wire clknet_leaf_362_clk_in_regs;
 wire clknet_leaf_363_clk_in_regs;
 wire clknet_leaf_364_clk_in_regs;
 wire clknet_leaf_365_clk_in_regs;
 wire clknet_leaf_366_clk_in_regs;
 wire clknet_leaf_367_clk_in_regs;
 wire clknet_leaf_368_clk_in_regs;
 wire clknet_leaf_369_clk_in_regs;
 wire clknet_leaf_370_clk_in_regs;
 wire clknet_leaf_371_clk_in_regs;
 wire clknet_leaf_372_clk_in_regs;
 wire clknet_leaf_373_clk_in_regs;
 wire clknet_leaf_374_clk_in_regs;
 wire clknet_leaf_375_clk_in_regs;
 wire clknet_leaf_376_clk_in_regs;
 wire clknet_leaf_377_clk_in_regs;
 wire clknet_leaf_378_clk_in_regs;
 wire clknet_leaf_379_clk_in_regs;
 wire clknet_leaf_381_clk_in_regs;
 wire clknet_leaf_383_clk_in_regs;
 wire clknet_leaf_384_clk_in_regs;
 wire clknet_leaf_385_clk_in_regs;
 wire clknet_leaf_387_clk_in_regs;
 wire clknet_leaf_388_clk_in_regs;
 wire clknet_leaf_389_clk_in_regs;
 wire clknet_leaf_390_clk_in_regs;
 wire clknet_leaf_391_clk_in_regs;
 wire clknet_leaf_392_clk_in_regs;
 wire clknet_leaf_393_clk_in_regs;
 wire clknet_leaf_394_clk_in_regs;
 wire clknet_leaf_395_clk_in_regs;
 wire clknet_leaf_396_clk_in_regs;
 wire clknet_leaf_397_clk_in_regs;
 wire clknet_leaf_398_clk_in_regs;
 wire clknet_leaf_399_clk_in_regs;
 wire clknet_leaf_400_clk_in_regs;
 wire clknet_leaf_401_clk_in_regs;
 wire clknet_leaf_402_clk_in_regs;
 wire clknet_leaf_403_clk_in_regs;
 wire clknet_leaf_404_clk_in_regs;
 wire clknet_leaf_405_clk_in_regs;
 wire clknet_leaf_406_clk_in_regs;
 wire clknet_leaf_407_clk_in_regs;
 wire clknet_leaf_408_clk_in_regs;
 wire clknet_leaf_409_clk_in_regs;
 wire clknet_leaf_410_clk_in_regs;
 wire clknet_leaf_411_clk_in_regs;
 wire clknet_leaf_412_clk_in_regs;
 wire clknet_leaf_413_clk_in_regs;
 wire clknet_leaf_414_clk_in_regs;
 wire clknet_leaf_415_clk_in_regs;
 wire clknet_leaf_416_clk_in_regs;
 wire clknet_leaf_417_clk_in_regs;
 wire clknet_leaf_418_clk_in_regs;
 wire clknet_leaf_419_clk_in_regs;
 wire clknet_leaf_421_clk_in_regs;
 wire clknet_leaf_423_clk_in_regs;
 wire clknet_leaf_424_clk_in_regs;
 wire clknet_leaf_425_clk_in_regs;
 wire clknet_leaf_426_clk_in_regs;
 wire clknet_leaf_427_clk_in_regs;
 wire clknet_leaf_428_clk_in_regs;
 wire clknet_leaf_429_clk_in_regs;
 wire clknet_leaf_430_clk_in_regs;
 wire clknet_leaf_431_clk_in_regs;
 wire clknet_leaf_432_clk_in_regs;
 wire clknet_leaf_433_clk_in_regs;
 wire clknet_leaf_434_clk_in_regs;
 wire clknet_leaf_435_clk_in_regs;
 wire clknet_leaf_436_clk_in_regs;
 wire clknet_leaf_437_clk_in_regs;
 wire clknet_leaf_438_clk_in_regs;
 wire clknet_leaf_439_clk_in_regs;
 wire clknet_leaf_440_clk_in_regs;
 wire clknet_leaf_441_clk_in_regs;
 wire clknet_leaf_442_clk_in_regs;
 wire clknet_leaf_443_clk_in_regs;
 wire clknet_leaf_444_clk_in_regs;
 wire clknet_leaf_445_clk_in_regs;
 wire clknet_leaf_446_clk_in_regs;
 wire clknet_leaf_447_clk_in_regs;
 wire clknet_leaf_448_clk_in_regs;
 wire clknet_leaf_449_clk_in_regs;
 wire clknet_leaf_450_clk_in_regs;
 wire clknet_leaf_451_clk_in_regs;
 wire clknet_leaf_452_clk_in_regs;
 wire clknet_leaf_453_clk_in_regs;
 wire clknet_leaf_454_clk_in_regs;
 wire clknet_leaf_455_clk_in_regs;
 wire clknet_leaf_456_clk_in_regs;
 wire clknet_leaf_457_clk_in_regs;
 wire clknet_leaf_458_clk_in_regs;
 wire clknet_leaf_459_clk_in_regs;
 wire clknet_leaf_460_clk_in_regs;
 wire clknet_leaf_461_clk_in_regs;
 wire clknet_leaf_462_clk_in_regs;
 wire clknet_leaf_463_clk_in_regs;
 wire clknet_leaf_464_clk_in_regs;
 wire clknet_leaf_465_clk_in_regs;
 wire clknet_leaf_466_clk_in_regs;
 wire clknet_leaf_467_clk_in_regs;
 wire clknet_leaf_468_clk_in_regs;
 wire clknet_leaf_469_clk_in_regs;
 wire clknet_leaf_470_clk_in_regs;
 wire clknet_leaf_471_clk_in_regs;
 wire clknet_leaf_472_clk_in_regs;
 wire clknet_leaf_473_clk_in_regs;
 wire clknet_leaf_474_clk_in_regs;
 wire clknet_leaf_475_clk_in_regs;
 wire clknet_leaf_476_clk_in_regs;
 wire clknet_leaf_477_clk_in_regs;
 wire clknet_leaf_478_clk_in_regs;
 wire clknet_leaf_479_clk_in_regs;
 wire clknet_leaf_480_clk_in_regs;
 wire clknet_leaf_481_clk_in_regs;
 wire clknet_leaf_482_clk_in_regs;
 wire clknet_leaf_483_clk_in_regs;
 wire clknet_leaf_484_clk_in_regs;
 wire clknet_leaf_485_clk_in_regs;
 wire clknet_leaf_486_clk_in_regs;
 wire clknet_leaf_487_clk_in_regs;
 wire clknet_leaf_488_clk_in_regs;
 wire clknet_leaf_489_clk_in_regs;
 wire clknet_leaf_490_clk_in_regs;
 wire clknet_leaf_491_clk_in_regs;
 wire clknet_leaf_492_clk_in_regs;
 wire clknet_leaf_493_clk_in_regs;
 wire clknet_leaf_494_clk_in_regs;
 wire clknet_leaf_495_clk_in_regs;
 wire clknet_leaf_496_clk_in_regs;
 wire clknet_leaf_497_clk_in_regs;
 wire clknet_leaf_498_clk_in_regs;
 wire clknet_leaf_499_clk_in_regs;
 wire clknet_leaf_500_clk_in_regs;
 wire clknet_leaf_501_clk_in_regs;
 wire clknet_leaf_502_clk_in_regs;
 wire clknet_leaf_503_clk_in_regs;
 wire clknet_leaf_504_clk_in_regs;
 wire clknet_leaf_505_clk_in_regs;
 wire clknet_leaf_506_clk_in_regs;
 wire clknet_leaf_507_clk_in_regs;
 wire clknet_leaf_508_clk_in_regs;
 wire clknet_leaf_509_clk_in_regs;
 wire clknet_leaf_510_clk_in_regs;
 wire clknet_leaf_511_clk_in_regs;
 wire clknet_leaf_512_clk_in_regs;
 wire clknet_leaf_513_clk_in_regs;
 wire clknet_leaf_515_clk_in_regs;
 wire clknet_leaf_519_clk_in_regs;
 wire clknet_leaf_520_clk_in_regs;
 wire clknet_leaf_525_clk_in_regs;
 wire clknet_leaf_527_clk_in_regs;
 wire clknet_leaf_528_clk_in_regs;
 wire clknet_leaf_529_clk_in_regs;
 wire clknet_leaf_530_clk_in_regs;
 wire clknet_leaf_531_clk_in_regs;
 wire clknet_leaf_532_clk_in_regs;
 wire clknet_leaf_533_clk_in_regs;
 wire clknet_leaf_534_clk_in_regs;
 wire clknet_leaf_535_clk_in_regs;
 wire clknet_leaf_536_clk_in_regs;
 wire clknet_leaf_537_clk_in_regs;
 wire clknet_leaf_538_clk_in_regs;
 wire clknet_leaf_542_clk_in_regs;
 wire clknet_leaf_543_clk_in_regs;
 wire clknet_leaf_544_clk_in_regs;
 wire clknet_leaf_545_clk_in_regs;
 wire clknet_leaf_546_clk_in_regs;
 wire clknet_leaf_547_clk_in_regs;
 wire clknet_leaf_549_clk_in_regs;
 wire clknet_leaf_550_clk_in_regs;
 wire clknet_leaf_551_clk_in_regs;
 wire clknet_leaf_554_clk_in_regs;
 wire clknet_leaf_555_clk_in_regs;
 wire clknet_leaf_557_clk_in_regs;
 wire clknet_leaf_559_clk_in_regs;
 wire clknet_leaf_560_clk_in_regs;
 wire clknet_leaf_561_clk_in_regs;
 wire clknet_leaf_562_clk_in_regs;
 wire clknet_leaf_564_clk_in_regs;
 wire clknet_leaf_565_clk_in_regs;
 wire clknet_leaf_566_clk_in_regs;
 wire clknet_leaf_567_clk_in_regs;
 wire clknet_leaf_568_clk_in_regs;
 wire clknet_leaf_570_clk_in_regs;
 wire clknet_leaf_572_clk_in_regs;
 wire clknet_leaf_573_clk_in_regs;
 wire clknet_leaf_574_clk_in_regs;
 wire clknet_leaf_575_clk_in_regs;
 wire clknet_leaf_576_clk_in_regs;
 wire clknet_leaf_577_clk_in_regs;
 wire clknet_leaf_578_clk_in_regs;
 wire clknet_leaf_579_clk_in_regs;
 wire clknet_leaf_580_clk_in_regs;
 wire clknet_leaf_584_clk_in_regs;
 wire clknet_leaf_585_clk_in_regs;
 wire clknet_leaf_586_clk_in_regs;
 wire clknet_leaf_587_clk_in_regs;
 wire clknet_leaf_588_clk_in_regs;
 wire clknet_leaf_589_clk_in_regs;
 wire clknet_leaf_590_clk_in_regs;
 wire clknet_leaf_591_clk_in_regs;
 wire clknet_leaf_592_clk_in_regs;
 wire clknet_leaf_593_clk_in_regs;
 wire clknet_leaf_594_clk_in_regs;
 wire clknet_leaf_595_clk_in_regs;
 wire clknet_leaf_596_clk_in_regs;
 wire clknet_leaf_597_clk_in_regs;
 wire clknet_leaf_598_clk_in_regs;
 wire clknet_leaf_599_clk_in_regs;
 wire clknet_leaf_600_clk_in_regs;
 wire clknet_leaf_601_clk_in_regs;
 wire clknet_leaf_602_clk_in_regs;
 wire clknet_leaf_603_clk_in_regs;
 wire clknet_leaf_604_clk_in_regs;
 wire clknet_leaf_605_clk_in_regs;
 wire clknet_leaf_606_clk_in_regs;
 wire clknet_leaf_607_clk_in_regs;
 wire clknet_leaf_608_clk_in_regs;
 wire clknet_leaf_609_clk_in_regs;
 wire clknet_leaf_610_clk_in_regs;
 wire clknet_leaf_611_clk_in_regs;
 wire clknet_leaf_612_clk_in_regs;
 wire clknet_leaf_613_clk_in_regs;
 wire clknet_leaf_614_clk_in_regs;
 wire clknet_leaf_615_clk_in_regs;
 wire clknet_leaf_616_clk_in_regs;
 wire clknet_leaf_617_clk_in_regs;
 wire clknet_leaf_618_clk_in_regs;
 wire clknet_leaf_619_clk_in_regs;
 wire clknet_leaf_620_clk_in_regs;
 wire clknet_leaf_621_clk_in_regs;
 wire clknet_leaf_622_clk_in_regs;
 wire clknet_leaf_623_clk_in_regs;
 wire clknet_leaf_624_clk_in_regs;
 wire clknet_leaf_625_clk_in_regs;
 wire clknet_leaf_626_clk_in_regs;
 wire clknet_leaf_627_clk_in_regs;
 wire clknet_leaf_628_clk_in_regs;
 wire clknet_leaf_629_clk_in_regs;
 wire clknet_leaf_630_clk_in_regs;
 wire clknet_leaf_632_clk_in_regs;
 wire clknet_leaf_633_clk_in_regs;
 wire clknet_leaf_634_clk_in_regs;
 wire clknet_leaf_635_clk_in_regs;
 wire clknet_leaf_636_clk_in_regs;
 wire clknet_leaf_637_clk_in_regs;
 wire clknet_leaf_638_clk_in_regs;
 wire clknet_leaf_640_clk_in_regs;
 wire clknet_leaf_641_clk_in_regs;
 wire clknet_leaf_642_clk_in_regs;
 wire clknet_leaf_643_clk_in_regs;
 wire clknet_leaf_644_clk_in_regs;
 wire clknet_leaf_645_clk_in_regs;
 wire clknet_leaf_646_clk_in_regs;
 wire clknet_leaf_647_clk_in_regs;
 wire clknet_leaf_648_clk_in_regs;
 wire clknet_leaf_649_clk_in_regs;
 wire clknet_leaf_650_clk_in_regs;
 wire clknet_leaf_651_clk_in_regs;
 wire clknet_leaf_652_clk_in_regs;
 wire clknet_leaf_653_clk_in_regs;
 wire clknet_leaf_654_clk_in_regs;
 wire clknet_leaf_655_clk_in_regs;
 wire clknet_leaf_656_clk_in_regs;
 wire clknet_leaf_657_clk_in_regs;
 wire clknet_leaf_658_clk_in_regs;
 wire clknet_leaf_659_clk_in_regs;
 wire clknet_leaf_660_clk_in_regs;
 wire clknet_leaf_661_clk_in_regs;
 wire clknet_leaf_662_clk_in_regs;
 wire clknet_leaf_663_clk_in_regs;
 wire clknet_leaf_664_clk_in_regs;
 wire clknet_leaf_665_clk_in_regs;
 wire clknet_leaf_666_clk_in_regs;
 wire clknet_leaf_667_clk_in_regs;
 wire clknet_leaf_669_clk_in_regs;
 wire clknet_leaf_671_clk_in_regs;
 wire clknet_leaf_672_clk_in_regs;
 wire clknet_leaf_673_clk_in_regs;
 wire clknet_leaf_675_clk_in_regs;
 wire clknet_leaf_678_clk_in_regs;
 wire clknet_leaf_679_clk_in_regs;
 wire clknet_leaf_680_clk_in_regs;
 wire clknet_leaf_681_clk_in_regs;
 wire clknet_leaf_682_clk_in_regs;
 wire clknet_leaf_683_clk_in_regs;
 wire clknet_leaf_684_clk_in_regs;
 wire clknet_leaf_685_clk_in_regs;
 wire clknet_leaf_686_clk_in_regs;
 wire clknet_leaf_687_clk_in_regs;
 wire clknet_leaf_688_clk_in_regs;
 wire clknet_leaf_689_clk_in_regs;
 wire clknet_leaf_690_clk_in_regs;
 wire clknet_leaf_691_clk_in_regs;
 wire clknet_leaf_692_clk_in_regs;
 wire clknet_leaf_694_clk_in_regs;
 wire clknet_leaf_695_clk_in_regs;
 wire clknet_leaf_696_clk_in_regs;
 wire clknet_leaf_697_clk_in_regs;
 wire clknet_leaf_698_clk_in_regs;
 wire clknet_leaf_700_clk_in_regs;
 wire clknet_leaf_701_clk_in_regs;
 wire clknet_leaf_702_clk_in_regs;
 wire clknet_leaf_703_clk_in_regs;
 wire clknet_leaf_704_clk_in_regs;
 wire clknet_leaf_705_clk_in_regs;
 wire clknet_leaf_706_clk_in_regs;
 wire clknet_leaf_707_clk_in_regs;
 wire clknet_leaf_708_clk_in_regs;
 wire clknet_leaf_709_clk_in_regs;
 wire clknet_leaf_711_clk_in_regs;
 wire clknet_leaf_712_clk_in_regs;
 wire clknet_leaf_715_clk_in_regs;
 wire clknet_leaf_716_clk_in_regs;
 wire clknet_leaf_717_clk_in_regs;
 wire clknet_leaf_718_clk_in_regs;
 wire clknet_leaf_719_clk_in_regs;
 wire clknet_leaf_720_clk_in_regs;
 wire clknet_leaf_721_clk_in_regs;
 wire clknet_leaf_722_clk_in_regs;
 wire clknet_leaf_723_clk_in_regs;
 wire clknet_leaf_724_clk_in_regs;
 wire clknet_leaf_725_clk_in_regs;
 wire clknet_leaf_726_clk_in_regs;
 wire clknet_leaf_727_clk_in_regs;
 wire clknet_leaf_728_clk_in_regs;
 wire clknet_leaf_729_clk_in_regs;
 wire clknet_leaf_730_clk_in_regs;
 wire clknet_leaf_731_clk_in_regs;
 wire clknet_leaf_732_clk_in_regs;
 wire clknet_leaf_733_clk_in_regs;
 wire clknet_leaf_734_clk_in_regs;
 wire clknet_leaf_735_clk_in_regs;
 wire clknet_leaf_736_clk_in_regs;
 wire clknet_leaf_737_clk_in_regs;
 wire clknet_leaf_738_clk_in_regs;
 wire clknet_leaf_739_clk_in_regs;
 wire clknet_leaf_740_clk_in_regs;
 wire clknet_leaf_741_clk_in_regs;
 wire clknet_leaf_742_clk_in_regs;
 wire clknet_leaf_743_clk_in_regs;
 wire clknet_leaf_744_clk_in_regs;
 wire clknet_leaf_745_clk_in_regs;
 wire clknet_leaf_746_clk_in_regs;
 wire clknet_leaf_748_clk_in_regs;
 wire clknet_leaf_749_clk_in_regs;
 wire clknet_leaf_750_clk_in_regs;
 wire clknet_leaf_751_clk_in_regs;
 wire clknet_leaf_752_clk_in_regs;
 wire clknet_leaf_753_clk_in_regs;
 wire clknet_leaf_754_clk_in_regs;
 wire clknet_leaf_755_clk_in_regs;
 wire clknet_leaf_756_clk_in_regs;
 wire clknet_leaf_757_clk_in_regs;
 wire clknet_leaf_758_clk_in_regs;
 wire clknet_leaf_759_clk_in_regs;
 wire clknet_leaf_760_clk_in_regs;
 wire clknet_leaf_761_clk_in_regs;
 wire clknet_leaf_762_clk_in_regs;
 wire clknet_leaf_763_clk_in_regs;
 wire clknet_leaf_764_clk_in_regs;
 wire clknet_leaf_765_clk_in_regs;
 wire clknet_leaf_766_clk_in_regs;
 wire clknet_leaf_767_clk_in_regs;
 wire clknet_leaf_768_clk_in_regs;
 wire clknet_leaf_769_clk_in_regs;
 wire clknet_leaf_770_clk_in_regs;
 wire clknet_leaf_771_clk_in_regs;
 wire clknet_leaf_772_clk_in_regs;
 wire clknet_leaf_773_clk_in_regs;
 wire clknet_leaf_774_clk_in_regs;
 wire clknet_leaf_776_clk_in_regs;
 wire clknet_leaf_777_clk_in_regs;
 wire clknet_leaf_778_clk_in_regs;
 wire clknet_leaf_779_clk_in_regs;
 wire clknet_leaf_781_clk_in_regs;
 wire clknet_leaf_783_clk_in_regs;
 wire clknet_leaf_784_clk_in_regs;
 wire clknet_leaf_785_clk_in_regs;
 wire clknet_leaf_786_clk_in_regs;
 wire clknet_leaf_787_clk_in_regs;
 wire clknet_leaf_788_clk_in_regs;
 wire clknet_leaf_789_clk_in_regs;
 wire clknet_leaf_790_clk_in_regs;
 wire clknet_0_clk_in_regs;
 wire clknet_1_0_0_clk_in_regs;
 wire clknet_1_1_0_clk_in_regs;
 wire clknet_3_0_0_clk_in_regs;
 wire clknet_3_1_0_clk_in_regs;
 wire clknet_3_2_0_clk_in_regs;
 wire clknet_3_3_0_clk_in_regs;
 wire clknet_3_4_0_clk_in_regs;
 wire clknet_3_5_0_clk_in_regs;
 wire clknet_3_6_0_clk_in_regs;
 wire clknet_3_7_0_clk_in_regs;
 wire clknet_5_0_0_clk_in_regs;
 wire clknet_5_1_0_clk_in_regs;
 wire clknet_5_2_0_clk_in_regs;
 wire clknet_5_3_0_clk_in_regs;
 wire clknet_5_4_0_clk_in_regs;
 wire clknet_5_5_0_clk_in_regs;
 wire clknet_5_6_0_clk_in_regs;
 wire clknet_5_7_0_clk_in_regs;
 wire clknet_5_8_0_clk_in_regs;
 wire clknet_5_9_0_clk_in_regs;
 wire clknet_5_10_0_clk_in_regs;
 wire clknet_5_11_0_clk_in_regs;
 wire clknet_5_12_0_clk_in_regs;
 wire clknet_5_13_0_clk_in_regs;
 wire clknet_5_14_0_clk_in_regs;
 wire clknet_5_15_0_clk_in_regs;
 wire clknet_5_16_0_clk_in_regs;
 wire clknet_5_17_0_clk_in_regs;
 wire clknet_5_18_0_clk_in_regs;
 wire clknet_5_19_0_clk_in_regs;
 wire clknet_5_20_0_clk_in_regs;
 wire clknet_5_21_0_clk_in_regs;
 wire clknet_5_22_0_clk_in_regs;
 wire clknet_5_23_0_clk_in_regs;
 wire clknet_5_24_0_clk_in_regs;
 wire clknet_5_25_0_clk_in_regs;
 wire clknet_5_26_0_clk_in_regs;
 wire clknet_5_27_0_clk_in_regs;
 wire clknet_5_28_0_clk_in_regs;
 wire clknet_5_29_0_clk_in_regs;
 wire clknet_5_30_0_clk_in_regs;
 wire clknet_5_31_0_clk_in_regs;
 wire clknet_6_0__leaf_clk_in_regs;
 wire clknet_6_1__leaf_clk_in_regs;
 wire clknet_6_2__leaf_clk_in_regs;
 wire clknet_6_3__leaf_clk_in_regs;
 wire clknet_6_4__leaf_clk_in_regs;
 wire clknet_6_5__leaf_clk_in_regs;
 wire clknet_6_6__leaf_clk_in_regs;
 wire clknet_6_7__leaf_clk_in_regs;
 wire clknet_6_8__leaf_clk_in_regs;
 wire clknet_6_9__leaf_clk_in_regs;
 wire clknet_6_10__leaf_clk_in_regs;
 wire clknet_6_11__leaf_clk_in_regs;
 wire clknet_6_12__leaf_clk_in_regs;
 wire clknet_6_13__leaf_clk_in_regs;
 wire clknet_6_14__leaf_clk_in_regs;
 wire clknet_6_15__leaf_clk_in_regs;
 wire clknet_6_16__leaf_clk_in_regs;
 wire clknet_6_17__leaf_clk_in_regs;
 wire clknet_6_18__leaf_clk_in_regs;
 wire clknet_6_19__leaf_clk_in_regs;
 wire clknet_6_20__leaf_clk_in_regs;
 wire clknet_6_21__leaf_clk_in_regs;
 wire clknet_6_22__leaf_clk_in_regs;
 wire clknet_6_23__leaf_clk_in_regs;
 wire clknet_6_24__leaf_clk_in_regs;
 wire clknet_6_25__leaf_clk_in_regs;
 wire clknet_6_26__leaf_clk_in_regs;
 wire clknet_6_27__leaf_clk_in_regs;
 wire clknet_6_28__leaf_clk_in_regs;
 wire clknet_6_29__leaf_clk_in_regs;
 wire clknet_6_30__leaf_clk_in_regs;
 wire clknet_6_31__leaf_clk_in_regs;
 wire clknet_6_32__leaf_clk_in_regs;
 wire clknet_6_33__leaf_clk_in_regs;
 wire clknet_6_34__leaf_clk_in_regs;
 wire clknet_6_35__leaf_clk_in_regs;
 wire clknet_6_36__leaf_clk_in_regs;
 wire clknet_6_37__leaf_clk_in_regs;
 wire clknet_6_38__leaf_clk_in_regs;
 wire clknet_6_39__leaf_clk_in_regs;
 wire clknet_6_40__leaf_clk_in_regs;
 wire clknet_6_41__leaf_clk_in_regs;
 wire clknet_6_42__leaf_clk_in_regs;
 wire clknet_6_43__leaf_clk_in_regs;
 wire clknet_6_44__leaf_clk_in_regs;
 wire clknet_6_45__leaf_clk_in_regs;
 wire clknet_6_46__leaf_clk_in_regs;
 wire clknet_6_47__leaf_clk_in_regs;
 wire clknet_6_48__leaf_clk_in_regs;
 wire clknet_6_49__leaf_clk_in_regs;
 wire clknet_6_50__leaf_clk_in_regs;
 wire clknet_6_51__leaf_clk_in_regs;
 wire clknet_6_52__leaf_clk_in_regs;
 wire clknet_6_53__leaf_clk_in_regs;
 wire clknet_6_54__leaf_clk_in_regs;
 wire clknet_6_55__leaf_clk_in_regs;
 wire clknet_6_56__leaf_clk_in_regs;
 wire clknet_6_57__leaf_clk_in_regs;
 wire clknet_6_58__leaf_clk_in_regs;
 wire clknet_6_59__leaf_clk_in_regs;
 wire clknet_6_60__leaf_clk_in_regs;
 wire clknet_6_61__leaf_clk_in_regs;
 wire clknet_6_62__leaf_clk_in_regs;
 wire clknet_6_63__leaf_clk_in_regs;
 wire delaynet_0_sys_clk_in;
 wire delaynet_1_sys_clk_in;
 wire delaynet_2_sys_clk_in;
 wire delaynet_3_sys_clk_in;
 wire delaynet_4_sys_clk_in;
 wire delaynet_5_sys_clk_in;
 wire delaynet_6_sys_clk_in;
 wire delaynet_7_sys_clk_in;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;

 sky130_fd_sc_hd__inv_1 _22645_ (.A(\inst$top.soc.cpu.sink__payload$24[36] ),
    .Y(_19826_));
 sky130_fd_sc_hd__nand3_1 _22646_ (.A(_19826_),
    .B(\inst$top.soc.cpu.sink__payload$24[34] ),
    .C(\inst$top.soc.cpu.sink__payload$24[35] ),
    .Y(_19827_));
 sky130_fd_sc_hd__clkinv_1 _22647_ (.A(\inst$top.soc.cpu.exception.w_trap ),
    .Y(_19828_));
 sky130_fd_sc_hd__nand3_1 _22648_ (.A(_19828_),
    .B(\inst$top.soc.cpu.d.sink__payload$16.rd_we ),
    .C(\inst$top.soc.cpu.m.source__valid ),
    .Y(_19829_));
 sky130_fd_sc_hd__clkinv_1 _22649_ (.A(_19829_),
    .Y(_19830_));
 sky130_fd_sc_hd__inv_1 _22650_ (.A(\inst$top.soc.cpu.sink__payload$24[33] ),
    .Y(_19831_));
 sky130_fd_sc_hd__nand3_1 _22651_ (.A(_19830_),
    .B(\inst$top.soc.cpu.sink__payload$24[32] ),
    .C(_19831_),
    .Y(_19832_));
 sky130_fd_sc_hd__nor2_1 _22652_ (.A(_19827_),
    .B(_19832_),
    .Y(_00133_));
 sky130_fd_sc_hd__inv_1 _22653_ (.A(\inst$top.soc.cpu.sink__payload$24[34] ),
    .Y(_19833_));
 sky130_fd_sc_hd__inv_1 _22654_ (.A(\inst$top.soc.cpu.sink__payload$24[35] ),
    .Y(_19834_));
 sky130_fd_sc_hd__nand3_1 _22655_ (.A(_19833_),
    .B(_19826_),
    .C(_19834_),
    .Y(_19835_));
 sky130_fd_sc_hd__inv_1 _22656_ (.A(\inst$top.soc.cpu.sink__payload$24[32] ),
    .Y(_19836_));
 sky130_fd_sc_hd__nand3_1 _22657_ (.A(_19830_),
    .B(_19836_),
    .C(\inst$top.soc.cpu.sink__payload$24[33] ),
    .Y(_19837_));
 sky130_fd_sc_hd__nor2_1 _22658_ (.A(_19835_),
    .B(_19837_),
    .Y(_00151_));
 sky130_fd_sc_hd__nor2_1 _22659_ (.A(_19827_),
    .B(_19837_),
    .Y(_00134_));
 sky130_fd_sc_hd__nand3_1 _22660_ (.A(_19833_),
    .B(_19826_),
    .C(\inst$top.soc.cpu.sink__payload$24[35] ),
    .Y(_19838_));
 sky130_fd_sc_hd__nand3_1 _22661_ (.A(_19830_),
    .B(_19836_),
    .C(_19831_),
    .Y(_19839_));
 sky130_fd_sc_hd__nor2_1 _22662_ (.A(_19838_),
    .B(_19839_),
    .Y(_00159_));
 sky130_fd_sc_hd__nor2_1 _22663_ (.A(_19827_),
    .B(_19839_),
    .Y(_00132_));
 sky130_fd_sc_hd__nor2_2 _22664_ (.A(_19835_),
    .B(_19832_),
    .Y(_00140_));
 sky130_fd_sc_hd__nor2_1 _22665_ (.A(_19838_),
    .B(_19832_),
    .Y(_00160_));
 sky130_fd_sc_hd__nand3_1 _22666_ (.A(_19826_),
    .B(_19834_),
    .C(\inst$top.soc.cpu.sink__payload$24[34] ),
    .Y(_19840_));
 sky130_fd_sc_hd__nand3_1 _22667_ (.A(_19830_),
    .B(\inst$top.soc.cpu.sink__payload$24[32] ),
    .C(\inst$top.soc.cpu.sink__payload$24[33] ),
    .Y(_19841_));
 sky130_fd_sc_hd__nor2_2 _22668_ (.A(_19840_),
    .B(_19841_),
    .Y(_00158_));
 sky130_fd_sc_hd__nor2_1 _22669_ (.A(_19838_),
    .B(_19837_),
    .Y(_00130_));
 sky130_fd_sc_hd__nor2_1 _22670_ (.A(_19838_),
    .B(_19841_),
    .Y(_00131_));
 sky130_fd_sc_hd__nor2_2 _22671_ (.A(_19835_),
    .B(_19841_),
    .Y(_00154_));
 sky130_fd_sc_hd__nor2_1 _22672_ (.A(_19827_),
    .B(_19841_),
    .Y(_00135_));
 sky130_fd_sc_hd__nor2_2 _22673_ (.A(_19840_),
    .B(_19837_),
    .Y(_00157_));
 sky130_fd_sc_hd__nand3_1 _22674_ (.A(\inst$top.soc.cpu.sink__payload$24[34] ),
    .B(\inst$top.soc.cpu.sink__payload$24[36] ),
    .C(\inst$top.soc.cpu.sink__payload$24[35] ),
    .Y(_19842_));
 sky130_fd_sc_hd__nor2_1 _22675_ (.A(_19842_),
    .B(_19841_),
    .Y(_00153_));
 sky130_fd_sc_hd__nor2_1 _22676_ (.A(_19842_),
    .B(_19837_),
    .Y(_00152_));
 sky130_fd_sc_hd__nor2_1 _22677_ (.A(_19842_),
    .B(_19832_),
    .Y(_00150_));
 sky130_fd_sc_hd__nor2_1 _22678_ (.A(_19842_),
    .B(_19839_),
    .Y(_00149_));
 sky130_fd_sc_hd__nand3_1 _22679_ (.A(_19833_),
    .B(\inst$top.soc.cpu.sink__payload$24[36] ),
    .C(\inst$top.soc.cpu.sink__payload$24[35] ),
    .Y(_19843_));
 sky130_fd_sc_hd__nor2_1 _22680_ (.A(_19843_),
    .B(_19841_),
    .Y(_00148_));
 sky130_fd_sc_hd__nor2_1 _22681_ (.A(_19843_),
    .B(_19837_),
    .Y(_00147_));
 sky130_fd_sc_hd__nor2_1 _22682_ (.A(_19843_),
    .B(_19832_),
    .Y(_00146_));
 sky130_fd_sc_hd__nor2_1 _22683_ (.A(_19843_),
    .B(_19839_),
    .Y(_00145_));
 sky130_fd_sc_hd__nand3_1 _22684_ (.A(_19834_),
    .B(\inst$top.soc.cpu.sink__payload$24[34] ),
    .C(\inst$top.soc.cpu.sink__payload$24[36] ),
    .Y(_19844_));
 sky130_fd_sc_hd__nor2_2 _22685_ (.A(_19844_),
    .B(_19841_),
    .Y(_00144_));
 sky130_fd_sc_hd__nor2_4 _22686_ (.A(_19844_),
    .B(_19837_),
    .Y(_00143_));
 sky130_fd_sc_hd__nor2_4 _22687_ (.A(_19844_),
    .B(_19832_),
    .Y(_00142_));
 sky130_fd_sc_hd__nor2_4 _22688_ (.A(_19844_),
    .B(_19839_),
    .Y(_00141_));
 sky130_fd_sc_hd__nand3_1 _22689_ (.A(_19833_),
    .B(_19834_),
    .C(\inst$top.soc.cpu.sink__payload$24[36] ),
    .Y(_19845_));
 sky130_fd_sc_hd__nor2_2 _22690_ (.A(_19845_),
    .B(_19841_),
    .Y(_00139_));
 sky130_fd_sc_hd__nor2_2 _22691_ (.A(_19845_),
    .B(_19837_),
    .Y(_00138_));
 sky130_fd_sc_hd__inv_2 _22693_ (.A(net2561),
    .Y(_19847_));
 sky130_fd_sc_hd__or2_2 _22695_ (.A(\inst$top.soc.cpu.loadstore.dbus__adr[1] ),
    .B(net2555),
    .X(_19849_));
 sky130_fd_sc_hd__o21ai_2 _22696_ (.A1(net2558),
    .A2(\inst$top.soc.cpu.fetch.ibus__adr[1] ),
    .B1(_19849_),
    .Y(_19850_));
 sky130_fd_sc_hd__inv_2 _22697_ (.A(_19850_),
    .Y(\inst$top.soc.bus__addr[3] ));
 sky130_fd_sc_hd__nand2_1 _22699_ (.A(net2555),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[0] ),
    .Y(_19852_));
 sky130_fd_sc_hd__nand2_1 _22701_ (.A(net2558),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[0] ),
    .Y(_19854_));
 sky130_fd_sc_hd__nand2_2 _22702_ (.A(_19852_),
    .B(_19854_),
    .Y(\inst$top.soc.bus__addr[2] ));
 sky130_fd_sc_hd__nand2_1 _22703_ (.A(net2555),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[4] ),
    .Y(_19855_));
 sky130_fd_sc_hd__nand2_1 _22704_ (.A(net2558),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[4] ),
    .Y(_19856_));
 sky130_fd_sc_hd__nand2_2 _22705_ (.A(_19855_),
    .B(_19856_),
    .Y(\inst$top.soc.bus__adr[4] ));
 sky130_fd_sc_hd__nand2_1 _22706_ (.A(net2555),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[3] ),
    .Y(_19857_));
 sky130_fd_sc_hd__nand2_1 _22707_ (.A(net2558),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[3] ),
    .Y(_19858_));
 sky130_fd_sc_hd__nand2_2 _22708_ (.A(_19857_),
    .B(_19858_),
    .Y(\inst$top.soc.bus__adr[3] ));
 sky130_fd_sc_hd__mux2i_1 _22709_ (.A0(\inst$top.soc.cpu.fetch.ibus__adr[6] ),
    .A1(\inst$top.soc.cpu.loadstore.dbus__adr[6] ),
    .S(net2559),
    .Y(_19859_));
 sky130_fd_sc_hd__inv_2 _22710_ (.A(_19859_),
    .Y(\inst$top.soc.bus__adr[6] ));
 sky130_fd_sc_hd__nand2_1 _22711_ (.A(net2555),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[5] ),
    .Y(_19860_));
 sky130_fd_sc_hd__nand2_1 _22712_ (.A(net2558),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[5] ),
    .Y(_19861_));
 sky130_fd_sc_hd__nand2_2 _22713_ (.A(_19860_),
    .B(_19861_),
    .Y(\inst$top.soc.bus__adr[5] ));
 sky130_fd_sc_hd__nand2_1 _22715_ (.A(net2556),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[7] ),
    .Y(_19863_));
 sky130_fd_sc_hd__nand2_1 _22717_ (.A(net2559),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[7] ),
    .Y(_19865_));
 sky130_fd_sc_hd__nand2_2 _22718_ (.A(_19863_),
    .B(_19865_),
    .Y(\inst$top.soc.bus__adr[7] ));
 sky130_fd_sc_hd__inv_2 _22719_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[0] ),
    .Y(_02706_));
 sky130_fd_sc_hd__nor2_2 _22720_ (.A(_19845_),
    .B(_19832_),
    .Y(_00137_));
 sky130_fd_sc_hd__nor2_2 _22721_ (.A(_19840_),
    .B(_19839_),
    .Y(_00155_));
 sky130_fd_sc_hd__or2_1 _22723_ (.A(\inst$top.soc.cpu.loadstore.dbus__adr[2] ),
    .B(net2555),
    .X(_19867_));
 sky130_fd_sc_hd__o21ai_4 _22724_ (.A1(net2558),
    .A2(\inst$top.soc.cpu.fetch.ibus__adr[2] ),
    .B1(_19867_),
    .Y(_19868_));
 sky130_fd_sc_hd__inv_2 _22725_ (.A(_19868_),
    .Y(\inst$top.soc.bus__adr[2] ));
 sky130_fd_sc_hd__inv_1 _22726_ (.A(\inst$top.soc.cpu.sink__payload$12[31] ),
    .Y(_19869_));
 sky130_fd_sc_hd__inv_2 _22727_ (.A(\inst$top.soc.cpu.d.sink__payload.auipc ),
    .Y(_19870_));
 sky130_fd_sc_hd__nor2_4 _22728_ (.A(\inst$top.soc.cpu.d.sink__payload.lui ),
    .B(_19870_),
    .Y(_19871_));
 sky130_fd_sc_hd__inv_2 _22729_ (.A(_19871_),
    .Y(_19872_));
 sky130_fd_sc_hd__inv_1 _22732_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[31] ),
    .Y(_19875_));
 sky130_fd_sc_hd__nand2_1 _22734_ (.A(_19875_),
    .B(net2886),
    .Y(_19877_));
 sky130_fd_sc_hd__nor2_1 _22735_ (.A(\inst$top.soc.cpu.d.sink__payload.auipc ),
    .B(\inst$top.soc.cpu.d.sink__payload.lui ),
    .Y(_19878_));
 sky130_fd_sc_hd__nand2_2 _22736_ (.A(net2850),
    .B(net2842),
    .Y(_19879_));
 sky130_fd_sc_hd__nand2_1 _22737_ (.A(_19878_),
    .B(_19879_),
    .Y(_19880_));
 sky130_fd_sc_hd__inv_2 _22738_ (.A(_19880_),
    .Y(_19881_));
 sky130_fd_sc_hd__o211ai_1 _22739_ (.A1(\inst$top.soc.cpu.gprf.mem_rp1__data[31] ),
    .A2(net2887),
    .B1(_19877_),
    .C1(net1828),
    .Y(_19882_));
 sky130_fd_sc_hd__o21ai_2 _22740_ (.A1(_19869_),
    .A2(net1832),
    .B1(_19882_),
    .Y(_19883_));
 sky130_fd_sc_hd__inv_2 _22741_ (.A(net1481),
    .Y(_19884_));
 sky130_fd_sc_hd__inv_2 _22743_ (.A(\inst$top.soc.cpu.d.sink__payload.rs2_re ),
    .Y(_19885_));
 sky130_fd_sc_hd__nor2_4 _22744_ (.A(\inst$top.soc.cpu.d.sink__payload.store ),
    .B(_19885_),
    .Y(_19886_));
 sky130_fd_sc_hd__inv_2 _22747_ (.A(net2884),
    .Y(_19889_));
 sky130_fd_sc_hd__nand2_1 _22751_ (.A(net2554),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[31] ),
    .Y(_19893_));
 sky130_fd_sc_hd__nand2_1 _22754_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[31] ),
    .B(net2883),
    .Y(_19896_));
 sky130_fd_sc_hd__nand3_1 _22755_ (.A(net1989),
    .B(_19893_),
    .C(_19896_),
    .Y(_19897_));
 sky130_fd_sc_hd__o21ai_2 _22756_ (.A1(\inst$top.soc.cpu.sink__payload$12[140] ),
    .A2(net1989),
    .B1(_19897_),
    .Y(_19898_));
 sky130_fd_sc_hd__inv_2 _22757_ (.A(net1739),
    .Y(_19899_));
 sky130_fd_sc_hd__inv_1 _22759_ (.A(\inst$top.soc.cpu.sink__payload$12[30] ),
    .Y(_19900_));
 sky130_fd_sc_hd__inv_2 _22761_ (.A(net2888),
    .Y(_19902_));
 sky130_fd_sc_hd__inv_1 _22764_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[30] ),
    .Y(_19905_));
 sky130_fd_sc_hd__nand2_1 _22765_ (.A(net2546),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[30] ),
    .Y(_19906_));
 sky130_fd_sc_hd__o21ai_0 _22766_ (.A1(net2546),
    .A2(_19905_),
    .B1(_19906_),
    .Y(_19907_));
 sky130_fd_sc_hd__nand2_1 _22768_ (.A(_19907_),
    .B(net1830),
    .Y(_19909_));
 sky130_fd_sc_hd__o21ai_2 _22769_ (.A1(_19900_),
    .A2(net1831),
    .B1(_19909_),
    .Y(_19910_));
 sky130_fd_sc_hd__inv_1 _22771_ (.A(\inst$top.soc.cpu.sink__payload$12[139] ),
    .Y(_19911_));
 sky130_fd_sc_hd__inv_1 _22774_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[30] ),
    .Y(_19914_));
 sky130_fd_sc_hd__nand2_1 _22775_ (.A(net2552),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[30] ),
    .Y(_19915_));
 sky130_fd_sc_hd__o21ai_2 _22776_ (.A1(net2551),
    .A2(_19914_),
    .B1(_19915_),
    .Y(_19916_));
 sky130_fd_sc_hd__nand2_1 _22777_ (.A(_19916_),
    .B(net1986),
    .Y(_19917_));
 sky130_fd_sc_hd__o21ai_2 _22778_ (.A1(_19911_),
    .A2(net1986),
    .B1(_19917_),
    .Y(_19918_));
 sky130_fd_sc_hd__inv_1 _22779_ (.A(net1473),
    .Y(_19919_));
 sky130_fd_sc_hd__inv_1 _22781_ (.A(\inst$top.soc.cpu.sink__payload$12[29] ),
    .Y(_19920_));
 sky130_fd_sc_hd__inv_1 _22782_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[29] ),
    .Y(_19921_));
 sky130_fd_sc_hd__nand2_1 _22783_ (.A(_19921_),
    .B(net2888),
    .Y(_19922_));
 sky130_fd_sc_hd__o211ai_1 _22784_ (.A1(net2888),
    .A2(\inst$top.soc.cpu.gprf.mem_rp1__data[29] ),
    .B1(_19922_),
    .C1(net1829),
    .Y(_19923_));
 sky130_fd_sc_hd__o21ai_2 _22785_ (.A1(_19920_),
    .A2(_19872_),
    .B1(_19923_),
    .Y(_19924_));
 sky130_fd_sc_hd__inv_1 _22787_ (.A(\inst$top.soc.cpu.sink__payload$12[138] ),
    .Y(_19925_));
 sky130_fd_sc_hd__inv_1 _22788_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[29] ),
    .Y(_19926_));
 sky130_fd_sc_hd__nand2_1 _22789_ (.A(net2554),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[29] ),
    .Y(_19927_));
 sky130_fd_sc_hd__o21ai_4 _22790_ (.A1(net2553),
    .A2(_19926_),
    .B1(_19927_),
    .Y(_19928_));
 sky130_fd_sc_hd__nand2_1 _22791_ (.A(_19928_),
    .B(net1986),
    .Y(_19929_));
 sky130_fd_sc_hd__o21ai_1 _22792_ (.A1(_19925_),
    .A2(net1986),
    .B1(_19929_),
    .Y(_19930_));
 sky130_fd_sc_hd__inv_1 _22794_ (.A(net1465),
    .Y(_19932_));
 sky130_fd_sc_hd__nand2_1 _22797_ (.A(net2549),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[28] ),
    .Y(_19934_));
 sky130_fd_sc_hd__nand2_1 _22798_ (.A(net2888),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[28] ),
    .Y(_19935_));
 sky130_fd_sc_hd__nand2_1 _22799_ (.A(_19934_),
    .B(_19935_),
    .Y(_19936_));
 sky130_fd_sc_hd__a22oi_2 _22800_ (.A1(\inst$top.soc.cpu.sink__payload$12[28] ),
    .A2(_19871_),
    .B1(net1828),
    .B2(_19936_),
    .Y(_19937_));
 sky130_fd_sc_hd__inv_2 _22801_ (.A(net1735),
    .Y(_19938_));
 sky130_fd_sc_hd__inv_1 _22803_ (.A(\inst$top.soc.cpu.sink__payload$12[137] ),
    .Y(_19939_));
 sky130_fd_sc_hd__nand2_1 _22804_ (.A(net2553),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[28] ),
    .Y(_19940_));
 sky130_fd_sc_hd__nand2_1 _22805_ (.A(net2884),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[28] ),
    .Y(_19941_));
 sky130_fd_sc_hd__nand2_1 _22806_ (.A(_19940_),
    .B(_19941_),
    .Y(_19942_));
 sky130_fd_sc_hd__nand2_1 _22807_ (.A(_19942_),
    .B(net1987),
    .Y(_19943_));
 sky130_fd_sc_hd__o21ai_0 _22808_ (.A1(_19939_),
    .A2(net1987),
    .B1(_19943_),
    .Y(_19944_));
 sky130_fd_sc_hd__inv_2 _22810_ (.A(net1457),
    .Y(_19946_));
 sky130_fd_sc_hd__inv_1 _22812_ (.A(\inst$top.soc.cpu.sink__payload$12[27] ),
    .Y(_19947_));
 sky130_fd_sc_hd__inv_1 _22813_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[27] ),
    .Y(_19948_));
 sky130_fd_sc_hd__nand2_1 _22814_ (.A(net2549),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[27] ),
    .Y(_19949_));
 sky130_fd_sc_hd__o21ai_0 _22815_ (.A1(net2549),
    .A2(_19948_),
    .B1(_19949_),
    .Y(_19950_));
 sky130_fd_sc_hd__nand2_1 _22816_ (.A(_19950_),
    .B(net1829),
    .Y(_19951_));
 sky130_fd_sc_hd__o21ai_4 _22817_ (.A1(_19947_),
    .A2(net1831),
    .B1(_19951_),
    .Y(_19952_));
 sky130_fd_sc_hd__nand2_1 _22820_ (.A(net2553),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[27] ),
    .Y(_19954_));
 sky130_fd_sc_hd__nand2_1 _22821_ (.A(net2882),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[27] ),
    .Y(_19955_));
 sky130_fd_sc_hd__nand3_1 _22822_ (.A(net1988),
    .B(_19954_),
    .C(_19955_),
    .Y(_19956_));
 sky130_fd_sc_hd__o21a_1 _22823_ (.A1(\inst$top.soc.cpu.sink__payload$12[136] ),
    .A2(net1989),
    .B1(_19956_),
    .X(_19957_));
 sky130_fd_sc_hd__nand2_1 _22826_ (.A(net2551),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[26] ),
    .Y(_19959_));
 sky130_fd_sc_hd__nand2_1 _22827_ (.A(net2882),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[26] ),
    .Y(_19960_));
 sky130_fd_sc_hd__nand3_1 _22828_ (.A(net1987),
    .B(_19959_),
    .C(_19960_),
    .Y(_19961_));
 sky130_fd_sc_hd__o21a_1 _22829_ (.A1(\inst$top.soc.cpu.sink__payload$12[135] ),
    .A2(net1987),
    .B1(_19961_),
    .X(_19962_));
 sky130_fd_sc_hd__nand2_1 _22832_ (.A(net2551),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[25] ),
    .Y(_19964_));
 sky130_fd_sc_hd__nand2_1 _22833_ (.A(net2882),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[25] ),
    .Y(_19965_));
 sky130_fd_sc_hd__nand3_1 _22834_ (.A(net1988),
    .B(_19964_),
    .C(_19965_),
    .Y(_19966_));
 sky130_fd_sc_hd__o21a_1 _22835_ (.A1(\inst$top.soc.cpu.sink__payload$12[134] ),
    .A2(net1988),
    .B1(_19966_),
    .X(_19967_));
 sky130_fd_sc_hd__inv_2 _22838_ (.A(_02616_),
    .Y(_02196_));
 sky130_fd_sc_hd__nand2_1 _22839_ (.A(net2553),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[24] ),
    .Y(_19969_));
 sky130_fd_sc_hd__nand2_1 _22840_ (.A(net2884),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[24] ),
    .Y(_19970_));
 sky130_fd_sc_hd__and2_2 _22841_ (.A(_19969_),
    .B(_19970_),
    .X(_19971_));
 sky130_fd_sc_hd__nand2_1 _22842_ (.A(_19971_),
    .B(net1986),
    .Y(_19972_));
 sky130_fd_sc_hd__o21ai_4 _22843_ (.A1(\inst$top.soc.cpu.sink__payload$12[133] ),
    .A2(net1986),
    .B1(_19972_),
    .Y(_19973_));
 sky130_fd_sc_hd__inv_1 _22844_ (.A(net1450),
    .Y(_19974_));
 sky130_fd_sc_hd__inv_2 _22847_ (.A(net1989),
    .Y(_19976_));
 sky130_fd_sc_hd__inv_1 _22850_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[23] ),
    .Y(_19979_));
 sky130_fd_sc_hd__nand2_1 _22851_ (.A(_19979_),
    .B(net2885),
    .Y(_19980_));
 sky130_fd_sc_hd__o21ai_1 _22852_ (.A1(net2883),
    .A2(\inst$top.soc.cpu.gprf.mem_rp2__data[23] ),
    .B1(_19980_),
    .Y(_19981_));
 sky130_fd_sc_hd__nand2_1 _22853_ (.A(net1825),
    .B(\inst$top.soc.cpu.sink__payload$12[132] ),
    .Y(_19982_));
 sky130_fd_sc_hd__o21ai_1 _22854_ (.A1(net1825),
    .A2(net1824),
    .B1(_19982_),
    .Y(_19983_));
 sky130_fd_sc_hd__inv_1 _22855_ (.A(net1447),
    .Y(_19984_));
 sky130_fd_sc_hd__inv_1 _22858_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[22] ),
    .Y(_19986_));
 sky130_fd_sc_hd__nand2_1 _22859_ (.A(_19986_),
    .B(net2885),
    .Y(_19987_));
 sky130_fd_sc_hd__o21ai_1 _22860_ (.A1(net2885),
    .A2(\inst$top.soc.cpu.gprf.mem_rp2__data[22] ),
    .B1(_19987_),
    .Y(_19988_));
 sky130_fd_sc_hd__nand2_1 _22861_ (.A(net1826),
    .B(\inst$top.soc.cpu.sink__payload$12[131] ),
    .Y(_19989_));
 sky130_fd_sc_hd__o21ai_1 _22862_ (.A1(net1826),
    .A2(net1823),
    .B1(_19989_),
    .Y(_19990_));
 sky130_fd_sc_hd__inv_1 _22864_ (.A(net1443),
    .Y(_19992_));
 sky130_fd_sc_hd__inv_1 _22866_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[21] ),
    .Y(_19993_));
 sky130_fd_sc_hd__nand2_1 _22867_ (.A(_19993_),
    .B(net2884),
    .Y(_19994_));
 sky130_fd_sc_hd__o21ai_2 _22868_ (.A1(net2884),
    .A2(\inst$top.soc.cpu.gprf.mem_rp2__data[21] ),
    .B1(_19994_),
    .Y(_19995_));
 sky130_fd_sc_hd__nand2_1 _22869_ (.A(_19995_),
    .B(net1987),
    .Y(_19996_));
 sky130_fd_sc_hd__o21ai_2 _22870_ (.A1(\inst$top.soc.cpu.sink__payload$12[130] ),
    .A2(net1987),
    .B1(_19996_),
    .Y(_19997_));
 sky130_fd_sc_hd__inv_2 _22871_ (.A(net1437),
    .Y(_19998_));
 sky130_fd_sc_hd__inv_1 _22873_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[20] ),
    .Y(_19999_));
 sky130_fd_sc_hd__nand2_1 _22874_ (.A(_19999_),
    .B(net2884),
    .Y(_20000_));
 sky130_fd_sc_hd__o21ai_1 _22875_ (.A1(net2884),
    .A2(\inst$top.soc.cpu.gprf.mem_rp2__data[20] ),
    .B1(_20000_),
    .Y(_20001_));
 sky130_fd_sc_hd__nand2_1 _22876_ (.A(net1827),
    .B(\inst$top.soc.cpu.sink__payload$12[129] ),
    .Y(_20002_));
 sky130_fd_sc_hd__o21a_2 _22877_ (.A1(net1827),
    .A2(net1822),
    .B1(_20002_),
    .X(_20003_));
 sky130_fd_sc_hd__inv_1 _22880_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[19] ),
    .Y(_20005_));
 sky130_fd_sc_hd__nand2_1 _22881_ (.A(_20005_),
    .B(net2883),
    .Y(_20006_));
 sky130_fd_sc_hd__o21ai_1 _22882_ (.A1(net2883),
    .A2(\inst$top.soc.cpu.gprf.mem_rp2__data[19] ),
    .B1(_20006_),
    .Y(_20007_));
 sky130_fd_sc_hd__nand2_1 _22883_ (.A(net1826),
    .B(\inst$top.soc.cpu.sink__payload$12[128] ),
    .Y(_20008_));
 sky130_fd_sc_hd__o21ai_1 _22884_ (.A1(net1826),
    .A2(_20007_),
    .B1(_20008_),
    .Y(_20009_));
 sky130_fd_sc_hd__inv_2 _22885_ (.A(net1435),
    .Y(_02983_));
 sky130_fd_sc_hd__or2_2 _22886_ (.A(net2884),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[18] ),
    .X(_20010_));
 sky130_fd_sc_hd__o21ai_1 _22887_ (.A1(\inst$top.soc.cpu.gprf.x_bypass2_data[18] ),
    .A2(net2551),
    .B1(_20010_),
    .Y(_20011_));
 sky130_fd_sc_hd__nand2_1 _22888_ (.A(_20011_),
    .B(net1988),
    .Y(_20012_));
 sky130_fd_sc_hd__o21ai_4 _22889_ (.A1(\inst$top.soc.cpu.sink__payload$12[127] ),
    .A2(net1988),
    .B1(_20012_),
    .Y(_20013_));
 sky130_fd_sc_hd__inv_2 _22891_ (.A(net1722),
    .Y(_20014_));
 sky130_fd_sc_hd__or2_2 _22893_ (.A(net2884),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[17] ),
    .X(_20015_));
 sky130_fd_sc_hd__o21ai_2 _22894_ (.A1(\inst$top.soc.cpu.gprf.x_bypass2_data[17] ),
    .A2(net2553),
    .B1(_20015_),
    .Y(_20016_));
 sky130_fd_sc_hd__nand2_1 _22895_ (.A(_20016_),
    .B(net1989),
    .Y(_20017_));
 sky130_fd_sc_hd__o21ai_2 _22896_ (.A1(\inst$top.soc.cpu.sink__payload$12[126] ),
    .A2(net1988),
    .B1(_20017_),
    .Y(_20018_));
 sky130_fd_sc_hd__clkinv_1 _22897_ (.A(net1717),
    .Y(_20019_));
 sky130_fd_sc_hd__or2_2 _22899_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_raw ),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[16] ),
    .X(_20020_));
 sky130_fd_sc_hd__o21ai_2 _22900_ (.A1(\inst$top.soc.cpu.gprf.x_bypass2_data[16] ),
    .A2(net2554),
    .B1(_20020_),
    .Y(_20021_));
 sky130_fd_sc_hd__nand2_1 _22901_ (.A(_20021_),
    .B(net1988),
    .Y(_20022_));
 sky130_fd_sc_hd__o21ai_2 _22902_ (.A1(\inst$top.soc.cpu.sink__payload$12[125] ),
    .A2(net1988),
    .B1(_20022_),
    .Y(_20023_));
 sky130_fd_sc_hd__clkinv_1 _22903_ (.A(net1716),
    .Y(_20024_));
 sky130_fd_sc_hd__nand2_1 _22905_ (.A(net2551),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[15] ),
    .Y(_20025_));
 sky130_fd_sc_hd__nand2_1 _22906_ (.A(net2882),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[15] ),
    .Y(_20026_));
 sky130_fd_sc_hd__nand2_1 _22907_ (.A(_20025_),
    .B(_20026_),
    .Y(_20027_));
 sky130_fd_sc_hd__or2_2 _22908_ (.A(\inst$top.soc.cpu.sink__payload$12[124] ),
    .B(net1988),
    .X(_20028_));
 sky130_fd_sc_hd__o21ai_2 _22909_ (.A1(_20027_),
    .A2(net1826),
    .B1(_20028_),
    .Y(_20029_));
 sky130_fd_sc_hd__inv_2 _22910_ (.A(net1710),
    .Y(_20030_));
 sky130_fd_sc_hd__inv_1 _22912_ (.A(\inst$top.soc.cpu.sink__payload$12[123] ),
    .Y(_20031_));
 sky130_fd_sc_hd__nand2_1 _22913_ (.A(net2551),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[14] ),
    .Y(_20032_));
 sky130_fd_sc_hd__nand2_1 _22914_ (.A(net2883),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[14] ),
    .Y(_20033_));
 sky130_fd_sc_hd__nand2_1 _22915_ (.A(_20032_),
    .B(_20033_),
    .Y(_20034_));
 sky130_fd_sc_hd__nand2_1 _22916_ (.A(_20034_),
    .B(net1986),
    .Y(_20035_));
 sky130_fd_sc_hd__o21ai_2 _22917_ (.A1(_20031_),
    .A2(net1986),
    .B1(_20035_),
    .Y(_20036_));
 sky130_fd_sc_hd__inv_2 _22918_ (.A(net1424),
    .Y(_03011_));
 sky130_fd_sc_hd__inv_1 _22919_ (.A(\inst$top.soc.cpu.sink__payload$12[122] ),
    .Y(_20037_));
 sky130_fd_sc_hd__nand2_1 _22920_ (.A(net2551),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[13] ),
    .Y(_20038_));
 sky130_fd_sc_hd__nand2_1 _22921_ (.A(net2883),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[13] ),
    .Y(_20039_));
 sky130_fd_sc_hd__nand2_1 _22922_ (.A(_20038_),
    .B(_20039_),
    .Y(_20040_));
 sky130_fd_sc_hd__nand2_1 _22923_ (.A(_20040_),
    .B(net1987),
    .Y(_20041_));
 sky130_fd_sc_hd__o21ai_2 _22924_ (.A1(_20037_),
    .A2(net1987),
    .B1(_20041_),
    .Y(_20042_));
 sky130_fd_sc_hd__clkinv_2 _22925_ (.A(net1420),
    .Y(_03017_));
 sky130_fd_sc_hd__inv_1 _22926_ (.A(\inst$top.soc.cpu.sink__payload$12[121] ),
    .Y(_20043_));
 sky130_fd_sc_hd__nand2_1 _22927_ (.A(net2553),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[12] ),
    .Y(_20044_));
 sky130_fd_sc_hd__nand2_1 _22928_ (.A(net2884),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[12] ),
    .Y(_20045_));
 sky130_fd_sc_hd__nand2_1 _22929_ (.A(_20044_),
    .B(_20045_),
    .Y(_20046_));
 sky130_fd_sc_hd__nand2_1 _22930_ (.A(_20046_),
    .B(_19886_),
    .Y(_20047_));
 sky130_fd_sc_hd__o21ai_0 _22931_ (.A1(_20043_),
    .A2(net1989),
    .B1(_20047_),
    .Y(_20048_));
 sky130_fd_sc_hd__inv_1 _22934_ (.A(\inst$top.soc.cpu.sink__payload$12[120] ),
    .Y(_20050_));
 sky130_fd_sc_hd__nand2_1 _22935_ (.A(net2553),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[11] ),
    .Y(_20051_));
 sky130_fd_sc_hd__nand2_1 _22936_ (.A(net2882),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[11] ),
    .Y(_20052_));
 sky130_fd_sc_hd__nand2_1 _22937_ (.A(_20051_),
    .B(_20052_),
    .Y(_20053_));
 sky130_fd_sc_hd__nand2_1 _22938_ (.A(_20053_),
    .B(net1989),
    .Y(_20054_));
 sky130_fd_sc_hd__o21ai_1 _22939_ (.A1(_20050_),
    .A2(net1989),
    .B1(_20054_),
    .Y(_20055_));
 sky130_fd_sc_hd__nand2_1 _22941_ (.A(net2553),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[10] ),
    .Y(_20056_));
 sky130_fd_sc_hd__nand2_1 _22942_ (.A(net2883),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[10] ),
    .Y(_20057_));
 sky130_fd_sc_hd__nand2_1 _22943_ (.A(_20056_),
    .B(_20057_),
    .Y(_20058_));
 sky130_fd_sc_hd__inv_1 _22944_ (.A(\inst$top.soc.cpu.sink__payload$12[119] ),
    .Y(_20059_));
 sky130_fd_sc_hd__nand2_1 _22945_ (.A(net1827),
    .B(_20059_),
    .Y(_20060_));
 sky130_fd_sc_hd__o21ai_4 _22946_ (.A1(net1827),
    .A2(_20058_),
    .B1(_20060_),
    .Y(_20061_));
 sky130_fd_sc_hd__inv_2 _22948_ (.A(_20061_),
    .Y(_20062_));
 sky130_fd_sc_hd__nand2_1 _22950_ (.A(net2554),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[9] ),
    .Y(_20063_));
 sky130_fd_sc_hd__nand2_1 _22951_ (.A(net2885),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[9] ),
    .Y(_20064_));
 sky130_fd_sc_hd__nand2_2 _22952_ (.A(_20063_),
    .B(_20064_),
    .Y(_20065_));
 sky130_fd_sc_hd__or2_2 _22953_ (.A(\inst$top.soc.cpu.sink__payload$12[118] ),
    .B(net1986),
    .X(_20066_));
 sky130_fd_sc_hd__o21ai_4 _22954_ (.A1(_20065_),
    .A2(net1826),
    .B1(_20066_),
    .Y(_20067_));
 sky130_fd_sc_hd__inv_2 _22956_ (.A(net1709),
    .Y(_20068_));
 sky130_fd_sc_hd__nand2_1 _22958_ (.A(net2553),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[8] ),
    .Y(_20069_));
 sky130_fd_sc_hd__nand2_1 _22959_ (.A(net2885),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[8] ),
    .Y(_20070_));
 sky130_fd_sc_hd__nand2_1 _22960_ (.A(_20069_),
    .B(_20070_),
    .Y(_20071_));
 sky130_fd_sc_hd__inv_1 _22961_ (.A(\inst$top.soc.cpu.sink__payload$12[117] ),
    .Y(_20072_));
 sky130_fd_sc_hd__nand2_1 _22962_ (.A(net1825),
    .B(_20072_),
    .Y(_20073_));
 sky130_fd_sc_hd__o21ai_2 _22963_ (.A1(net1825),
    .A2(_20071_),
    .B1(_20073_),
    .Y(_20074_));
 sky130_fd_sc_hd__inv_2 _22964_ (.A(net1400),
    .Y(_03045_));
 sky130_fd_sc_hd__nand2_1 _22965_ (.A(net2552),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[7] ),
    .Y(_20075_));
 sky130_fd_sc_hd__nand2_1 _22966_ (.A(net2882),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[7] ),
    .Y(_20076_));
 sky130_fd_sc_hd__nand2_1 _22967_ (.A(_20075_),
    .B(_20076_),
    .Y(_20077_));
 sky130_fd_sc_hd__inv_1 _22968_ (.A(_20077_),
    .Y(_20078_));
 sky130_fd_sc_hd__nand2_1 _22969_ (.A(net1825),
    .B(\inst$top.soc.cpu.sink__payload$12[116] ),
    .Y(_20079_));
 sky130_fd_sc_hd__o21ai_4 _22970_ (.A1(net1825),
    .A2(_20078_),
    .B1(_20079_),
    .Y(_20080_));
 sky130_fd_sc_hd__nand2_1 _22972_ (.A(net2552),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[6] ),
    .Y(_20081_));
 sky130_fd_sc_hd__nand2_1 _22973_ (.A(net2885),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[6] ),
    .Y(_20082_));
 sky130_fd_sc_hd__nand2_1 _22974_ (.A(_20081_),
    .B(_20082_),
    .Y(_20083_));
 sky130_fd_sc_hd__inv_1 _22975_ (.A(_20083_),
    .Y(_20084_));
 sky130_fd_sc_hd__nand2_1 _22976_ (.A(net1825),
    .B(\inst$top.soc.cpu.sink__payload$12[115] ),
    .Y(_20085_));
 sky130_fd_sc_hd__o21ai_4 _22977_ (.A1(net1825),
    .A2(_20084_),
    .B1(_20085_),
    .Y(_20086_));
 sky130_fd_sc_hd__nand2_1 _22979_ (.A(net2551),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[5] ),
    .Y(_20087_));
 sky130_fd_sc_hd__nand2_1 _22980_ (.A(net2883),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[5] ),
    .Y(_20088_));
 sky130_fd_sc_hd__nand2_1 _22981_ (.A(_20087_),
    .B(_20088_),
    .Y(_20089_));
 sky130_fd_sc_hd__inv_1 _22982_ (.A(_20089_),
    .Y(_20090_));
 sky130_fd_sc_hd__nand2_1 _22983_ (.A(net1825),
    .B(\inst$top.soc.cpu.sink__payload$12[114] ),
    .Y(_20091_));
 sky130_fd_sc_hd__o21ai_1 _22984_ (.A1(net1825),
    .A2(_20090_),
    .B1(_20091_),
    .Y(_20092_));
 sky130_fd_sc_hd__nand2_1 _22987_ (.A(net2553),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[4] ),
    .Y(_20094_));
 sky130_fd_sc_hd__nand2_1 _22988_ (.A(net2882),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[4] ),
    .Y(_20095_));
 sky130_fd_sc_hd__nand2_1 _22989_ (.A(_20094_),
    .B(_20095_),
    .Y(_20096_));
 sky130_fd_sc_hd__inv_2 _22990_ (.A(_20096_),
    .Y(_20097_));
 sky130_fd_sc_hd__nand2_1 _22991_ (.A(_20097_),
    .B(net1987),
    .Y(_20098_));
 sky130_fd_sc_hd__o21ai_2 _22992_ (.A1(\inst$top.soc.cpu.sink__payload$12[113] ),
    .A2(net1987),
    .B1(_20098_),
    .Y(_20099_));
 sky130_fd_sc_hd__inv_2 _22993_ (.A(net1199),
    .Y(_20100_));
 sky130_fd_sc_hd__nand2_1 _22996_ (.A(net2551),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[3] ),
    .Y(_20102_));
 sky130_fd_sc_hd__nand2_1 _22997_ (.A(net2882),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[3] ),
    .Y(_20103_));
 sky130_fd_sc_hd__nand2_1 _22998_ (.A(_20102_),
    .B(_20103_),
    .Y(_20104_));
 sky130_fd_sc_hd__nand2_1 _22999_ (.A(_20104_),
    .B(net1988),
    .Y(_20105_));
 sky130_fd_sc_hd__nand2_1 _23000_ (.A(net1826),
    .B(\inst$top.soc.cpu.sink__payload$12[112] ),
    .Y(_20106_));
 sky130_fd_sc_hd__nand2_1 _23001_ (.A(_20105_),
    .B(_20106_),
    .Y(_20107_));
 sky130_fd_sc_hd__nand2_1 _23005_ (.A(net2552),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[2] ),
    .Y(_20110_));
 sky130_fd_sc_hd__nand2_1 _23006_ (.A(net2882),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[2] ),
    .Y(_20111_));
 sky130_fd_sc_hd__nand2_1 _23007_ (.A(_20110_),
    .B(_20111_),
    .Y(_20112_));
 sky130_fd_sc_hd__inv_1 _23008_ (.A(_20112_),
    .Y(_20113_));
 sky130_fd_sc_hd__nand2_1 _23009_ (.A(net1826),
    .B(\inst$top.soc.cpu.sink__payload$12[111] ),
    .Y(_20114_));
 sky130_fd_sc_hd__o21ai_1 _23010_ (.A1(net1826),
    .A2(_20113_),
    .B1(_20114_),
    .Y(_20115_));
 sky130_fd_sc_hd__inv_1 _23013_ (.A(_19879_),
    .Y(_20117_));
 sky130_fd_sc_hd__inv_1 _23014_ (.A(\inst$top.soc.cpu.sink__payload$12[102] ),
    .Y(_20118_));
 sky130_fd_sc_hd__inv_1 _23015_ (.A(_19878_),
    .Y(_20119_));
 sky130_fd_sc_hd__a21oi_1 _23016_ (.A1(_20117_),
    .A2(_20118_),
    .B1(_20119_),
    .Y(_20120_));
 sky130_fd_sc_hd__nand2_1 _23017_ (.A(net2546),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[1] ),
    .Y(_20121_));
 sky130_fd_sc_hd__nand2_1 _23018_ (.A(net2886),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[1] ),
    .Y(_20122_));
 sky130_fd_sc_hd__nand3_1 _23019_ (.A(_20121_),
    .B(_19879_),
    .C(_20122_),
    .Y(_20123_));
 sky130_fd_sc_hd__nand2_2 _23020_ (.A(_20120_),
    .B(_20123_),
    .Y(_20124_));
 sky130_fd_sc_hd__nand2_1 _23022_ (.A(net2552),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[1] ),
    .Y(_20125_));
 sky130_fd_sc_hd__nand2_1 _23023_ (.A(net2882),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[1] ),
    .Y(_20126_));
 sky130_fd_sc_hd__nand2_1 _23024_ (.A(_20125_),
    .B(_20126_),
    .Y(_20127_));
 sky130_fd_sc_hd__or2_2 _23025_ (.A(\inst$top.soc.cpu.sink__payload$12[110] ),
    .B(_19886_),
    .X(_20128_));
 sky130_fd_sc_hd__o21ai_4 _23026_ (.A1(_20127_),
    .A2(net1827),
    .B1(_20128_),
    .Y(_20129_));
 sky130_fd_sc_hd__clkinv_1 _23027_ (.A(net1703),
    .Y(_20130_));
 sky130_fd_sc_hd__nand2_1 _23030_ (.A(net2546),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[0] ),
    .Y(_20132_));
 sky130_fd_sc_hd__nand2_1 _23031_ (.A(net2886),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[0] ),
    .Y(_20133_));
 sky130_fd_sc_hd__nand2_1 _23032_ (.A(_20132_),
    .B(_20133_),
    .Y(_20134_));
 sky130_fd_sc_hd__nor2_1 _23033_ (.A(\inst$top.soc.cpu.sink__payload$12[101] ),
    .B(_19879_),
    .Y(_20135_));
 sky130_fd_sc_hd__nor2_1 _23034_ (.A(_20119_),
    .B(_20135_),
    .Y(_20136_));
 sky130_fd_sc_hd__o21ai_1 _23035_ (.A1(_20117_),
    .A2(_20134_),
    .B1(_20136_),
    .Y(_20137_));
 sky130_fd_sc_hd__inv_1 _23037_ (.A(\inst$top.soc.cpu.d.sink__payload.rd_we ),
    .Y(_20138_));
 sky130_fd_sc_hd__nand3_1 _23039_ (.A(net2891),
    .B(\inst$top.soc.cpu.exception.m_mip.meip ),
    .C(\inst$top.soc.cpu.exception.m_mie.meie ),
    .Y(_20140_));
 sky130_fd_sc_hd__inv_2 _23040_ (.A(_20140_),
    .Y(_20141_));
 sky130_fd_sc_hd__nand3_1 _23041_ (.A(\inst$top.soc.cpu.exception.m_mip[3] ),
    .B(\inst$top.soc.cpu.exception.m_mie[3] ),
    .C(net2891),
    .Y(_20142_));
 sky130_fd_sc_hd__nand3_1 _23042_ (.A(net2890),
    .B(\inst$top.soc.cpu.exception.m_mip[4] ),
    .C(\inst$top.soc.cpu.exception.m_mie[4] ),
    .Y(_20143_));
 sky130_fd_sc_hd__nand2_1 _23043_ (.A(_20142_),
    .B(_20143_),
    .Y(_20144_));
 sky130_fd_sc_hd__nor2_1 _23044_ (.A(_20141_),
    .B(_20144_),
    .Y(_20145_));
 sky130_fd_sc_hd__nand3_1 _23045_ (.A(net2891),
    .B(\inst$top.soc.cpu.exception.m_mip.msip ),
    .C(\inst$top.soc.cpu.exception.m_mie.msie ),
    .Y(_20146_));
 sky130_fd_sc_hd__nand3_1 _23046_ (.A(net2891),
    .B(\inst$top.soc.cpu.exception.m_mip.mtip ),
    .C(\inst$top.soc.cpu.exception.m_mie.mtie ),
    .Y(_20147_));
 sky130_fd_sc_hd__nand2_1 _23047_ (.A(_20146_),
    .B(_20147_),
    .Y(_20148_));
 sky130_fd_sc_hd__inv_2 _23048_ (.A(_20148_),
    .Y(_20149_));
 sky130_fd_sc_hd__nand2_2 _23049_ (.A(_20145_),
    .B(_20149_),
    .Y(_20150_));
 sky130_fd_sc_hd__nand3_1 _23050_ (.A(net2891),
    .B(\inst$top.soc.cpu.exception.m_mip[5] ),
    .C(\inst$top.soc.cpu.exception.m_mie[5] ),
    .Y(_20151_));
 sky130_fd_sc_hd__nand3_1 _23051_ (.A(net2890),
    .B(\inst$top.soc.cpu.exception.m_mip[6] ),
    .C(\inst$top.soc.cpu.exception.m_mie[6] ),
    .Y(_20152_));
 sky130_fd_sc_hd__nand2_1 _23052_ (.A(_20151_),
    .B(_20152_),
    .Y(_20153_));
 sky130_fd_sc_hd__nand3_1 _23053_ (.A(net2891),
    .B(\inst$top.soc.cpu.exception.m_mip[7] ),
    .C(\inst$top.soc.cpu.exception.m_mie[7] ),
    .Y(_20154_));
 sky130_fd_sc_hd__nand3_1 _23054_ (.A(net2890),
    .B(\inst$top.soc.cpu.exception.m_mip[8] ),
    .C(\inst$top.soc.cpu.exception.m_mie[8] ),
    .Y(_20155_));
 sky130_fd_sc_hd__nand2_1 _23055_ (.A(_20154_),
    .B(_20155_),
    .Y(_20156_));
 sky130_fd_sc_hd__nor2_1 _23056_ (.A(_20153_),
    .B(_20156_),
    .Y(_20157_));
 sky130_fd_sc_hd__nand3_1 _23057_ (.A(net2890),
    .B(\inst$top.soc.cpu.exception.m_mip[9] ),
    .C(\inst$top.soc.cpu.exception.m_mie[9] ),
    .Y(_20158_));
 sky130_fd_sc_hd__nand3_1 _23058_ (.A(net2890),
    .B(\inst$top.soc.cpu.exception.m_mip[10] ),
    .C(\inst$top.soc.cpu.exception.m_mie[10] ),
    .Y(_20159_));
 sky130_fd_sc_hd__nand2_1 _23059_ (.A(_20158_),
    .B(_20159_),
    .Y(_20160_));
 sky130_fd_sc_hd__nand3_1 _23061_ (.A(\inst$top.soc.cpu.exception.m_mstatus.mie ),
    .B(\inst$top.soc.cpu.exception.m_mip[11] ),
    .C(\inst$top.soc.cpu.exception.m_mie[11] ),
    .Y(_20162_));
 sky130_fd_sc_hd__nand3_1 _23062_ (.A(net2891),
    .B(\inst$top.soc.cpu.exception.m_mip[12] ),
    .C(\inst$top.soc.cpu.exception.m_mie[12] ),
    .Y(_20163_));
 sky130_fd_sc_hd__nand2_1 _23063_ (.A(_20162_),
    .B(_20163_),
    .Y(_20164_));
 sky130_fd_sc_hd__nor2_1 _23064_ (.A(_20160_),
    .B(_20164_),
    .Y(_20165_));
 sky130_fd_sc_hd__nand2_1 _23065_ (.A(_20157_),
    .B(_20165_),
    .Y(_20166_));
 sky130_fd_sc_hd__nor2_2 _23066_ (.A(_20150_),
    .B(_20166_),
    .Y(_20167_));
 sky130_fd_sc_hd__nand3_1 _23067_ (.A(net2890),
    .B(\inst$top.soc.cpu.exception.m_mip[17] ),
    .C(\inst$top.soc.cpu.exception.m_mie[17] ),
    .Y(_20168_));
 sky130_fd_sc_hd__nand3_1 _23068_ (.A(net2891),
    .B(\inst$top.soc.cpu.exception.m_mip[18] ),
    .C(\inst$top.soc.cpu.exception.m_mie[18] ),
    .Y(_20169_));
 sky130_fd_sc_hd__nand2_1 _23069_ (.A(_20168_),
    .B(_20169_),
    .Y(_20170_));
 sky130_fd_sc_hd__nand3_1 _23070_ (.A(net2890),
    .B(\inst$top.soc.cpu.exception.m_mip[14] ),
    .C(\inst$top.soc.cpu.exception.m_mie[14] ),
    .Y(_20171_));
 sky130_fd_sc_hd__nand3_1 _23071_ (.A(net2890),
    .B(\inst$top.soc.cpu.exception.m_mip[13] ),
    .C(\inst$top.soc.cpu.exception.m_mie[13] ),
    .Y(_20172_));
 sky130_fd_sc_hd__nand2_1 _23072_ (.A(_20171_),
    .B(_20172_),
    .Y(_20173_));
 sky130_fd_sc_hd__nand3_1 _23073_ (.A(net2890),
    .B(\inst$top.soc.cpu.exception.m_mip[15] ),
    .C(\inst$top.soc.cpu.exception.m_mie[15] ),
    .Y(_20174_));
 sky130_fd_sc_hd__nand3_1 _23074_ (.A(net2890),
    .B(\inst$top.soc.cpu.exception.m_mip[16] ),
    .C(\inst$top.soc.cpu.exception.m_mie[16] ),
    .Y(_20175_));
 sky130_fd_sc_hd__nand2_1 _23075_ (.A(_20174_),
    .B(_20175_),
    .Y(_20176_));
 sky130_fd_sc_hd__nor2_1 _23076_ (.A(_20173_),
    .B(_20176_),
    .Y(_20177_));
 sky130_fd_sc_hd__inv_1 _23077_ (.A(_20177_),
    .Y(_20178_));
 sky130_fd_sc_hd__nor2_1 _23078_ (.A(_20170_),
    .B(_20178_),
    .Y(_20179_));
 sky130_fd_sc_hd__nand2_1 _23079_ (.A(\inst$top.soc.cpu.d.sink__payload$6.loadstore_misaligned ),
    .B(\inst$top.soc.cpu.d.sink__payload$6.load ),
    .Y(_20180_));
 sky130_fd_sc_hd__o21ai_0 _23080_ (.A1(\inst$top.soc.cpu.sink__payload$18[181] ),
    .A2(\inst$top.soc.cpu.sink__payload$18[180] ),
    .B1(\inst$top.soc.cpu.d.sink__payload$6.branch_taken ),
    .Y(_20181_));
 sky130_fd_sc_hd__nor2_2 _23081_ (.A(\inst$top.soc.cpu.d.sink__payload$6.illegal ),
    .B(\inst$top.soc.cpu.d.sink__payload$6.ebreak ),
    .Y(_20182_));
 sky130_fd_sc_hd__nand2_1 _23082_ (.A(_20181_),
    .B(_20182_),
    .Y(_20183_));
 sky130_fd_sc_hd__nor2_1 _23083_ (.A(_20180_),
    .B(_20183_),
    .Y(_20184_));
 sky130_fd_sc_hd__nand3_1 _23084_ (.A(net1381),
    .B(_20179_),
    .C(_20184_),
    .Y(_20185_));
 sky130_fd_sc_hd__inv_1 _23086_ (.A(\inst$top.soc.cpu.d.sink__payload$6.load ),
    .Y(_20187_));
 sky130_fd_sc_hd__nand4_1 _23087_ (.A(_20182_),
    .B(\inst$top.soc.cpu.d.sink__payload$6.loadstore_misaligned ),
    .C(_20187_),
    .D(\inst$top.soc.cpu.d.sink__payload$6.store ),
    .Y(_20188_));
 sky130_fd_sc_hd__inv_2 _23088_ (.A(\inst$top.soc.cpu.d.sink__payload$6.branch_taken ),
    .Y(_02861_));
 sky130_fd_sc_hd__nor2_1 _23089_ (.A(\inst$top.soc.cpu.sink__payload$18[181] ),
    .B(\inst$top.soc.cpu.sink__payload$18[180] ),
    .Y(_20189_));
 sky130_fd_sc_hd__nor2_1 _23090_ (.A(_02861_),
    .B(_20189_),
    .Y(_20190_));
 sky130_fd_sc_hd__nor2_1 _23091_ (.A(_20190_),
    .B(_20170_),
    .Y(_20191_));
 sky130_fd_sc_hd__nand2_1 _23092_ (.A(_20177_),
    .B(_20191_),
    .Y(_20192_));
 sky130_fd_sc_hd__nor2_1 _23093_ (.A(_20188_),
    .B(_20192_),
    .Y(_20193_));
 sky130_fd_sc_hd__nand2_1 _23094_ (.A(net1381),
    .B(_20193_),
    .Y(_20194_));
 sky130_fd_sc_hd__nand2_1 _23095_ (.A(_20185_),
    .B(_20194_),
    .Y(_20195_));
 sky130_fd_sc_hd__nand2_1 _23096_ (.A(\inst$top.soc.cpu.d.sink__payload$6.loadstore_misaligned ),
    .B(\inst$top.soc.cpu.d.sink__payload$6.store ),
    .Y(_20196_));
 sky130_fd_sc_hd__nand3_1 _23097_ (.A(_20196_),
    .B(_20180_),
    .C(\inst$top.soc.cpu.d.sink__payload$6.ecall ),
    .Y(_20197_));
 sky130_fd_sc_hd__nor2_1 _23098_ (.A(_20197_),
    .B(_20183_),
    .Y(_20198_));
 sky130_fd_sc_hd__nand3_1 _23099_ (.A(_20167_),
    .B(_20179_),
    .C(_20198_),
    .Y(_20199_));
 sky130_fd_sc_hd__nand2_1 _23100_ (.A(_20140_),
    .B(_20142_),
    .Y(_20200_));
 sky130_fd_sc_hd__nand2_1 _23101_ (.A(_20143_),
    .B(_20151_),
    .Y(_20201_));
 sky130_fd_sc_hd__nor2_1 _23102_ (.A(_20200_),
    .B(_20201_),
    .Y(_20202_));
 sky130_fd_sc_hd__nand2_1 _23103_ (.A(_20202_),
    .B(_20149_),
    .Y(_20203_));
 sky130_fd_sc_hd__nand2_1 _23104_ (.A(_20152_),
    .B(_20154_),
    .Y(_20204_));
 sky130_fd_sc_hd__nand2_1 _23105_ (.A(_20158_),
    .B(_20155_),
    .Y(_20205_));
 sky130_fd_sc_hd__nor2_1 _23106_ (.A(_20204_),
    .B(_20205_),
    .Y(_20206_));
 sky130_fd_sc_hd__nand2_1 _23107_ (.A(_20159_),
    .B(_20162_),
    .Y(_20207_));
 sky130_fd_sc_hd__nand2_1 _23108_ (.A(_20163_),
    .B(_20172_),
    .Y(_20208_));
 sky130_fd_sc_hd__nor2_1 _23109_ (.A(_20207_),
    .B(_20208_),
    .Y(_20209_));
 sky130_fd_sc_hd__nand2_1 _23110_ (.A(_20206_),
    .B(_20209_),
    .Y(_20210_));
 sky130_fd_sc_hd__nor2_1 _23111_ (.A(_20203_),
    .B(_20210_),
    .Y(_20211_));
 sky130_fd_sc_hd__inv_1 _23112_ (.A(\inst$top.soc.cpu.d.sink__payload$6.illegal ),
    .Y(_20212_));
 sky130_fd_sc_hd__nand4_1 _23113_ (.A(_20181_),
    .B(_20212_),
    .C(\inst$top.soc.cpu.d.sink__payload$6.ebreak ),
    .D(_20169_),
    .Y(_20213_));
 sky130_fd_sc_hd__nand2_1 _23114_ (.A(_20171_),
    .B(_20174_),
    .Y(_20214_));
 sky130_fd_sc_hd__inv_1 _23115_ (.A(_20214_),
    .Y(_20215_));
 sky130_fd_sc_hd__nand3_1 _23116_ (.A(_20215_),
    .B(_20168_),
    .C(_20175_),
    .Y(_20216_));
 sky130_fd_sc_hd__nor2_1 _23117_ (.A(_20213_),
    .B(_20216_),
    .Y(_20217_));
 sky130_fd_sc_hd__nand2_1 _23118_ (.A(_20211_),
    .B(_20217_),
    .Y(_20218_));
 sky130_fd_sc_hd__nor2_1 _23119_ (.A(_20212_),
    .B(_20192_),
    .Y(_20219_));
 sky130_fd_sc_hd__nand2_1 _23120_ (.A(net1381),
    .B(_20219_),
    .Y(_20220_));
 sky130_fd_sc_hd__nand3_1 _23121_ (.A(_20199_),
    .B(_20218_),
    .C(net1192),
    .Y(_20221_));
 sky130_fd_sc_hd__nor2_1 _23122_ (.A(net1068),
    .B(_20221_),
    .Y(_20222_));
 sky130_fd_sc_hd__inv_1 _23123_ (.A(\inst$top.soc.cpu.d.sink__payload$6.mret ),
    .Y(_20223_));
 sky130_fd_sc_hd__nand2_1 _23124_ (.A(net1381),
    .B(_20179_),
    .Y(_20224_));
 sky130_fd_sc_hd__inv_1 _23125_ (.A(_20224_),
    .Y(_20225_));
 sky130_fd_sc_hd__nand2_1 _23126_ (.A(_20225_),
    .B(_20190_),
    .Y(_20226_));
 sky130_fd_sc_hd__nand4_1 _23127_ (.A(_20222_),
    .B(net2538),
    .C(_20225_),
    .D(net1018),
    .Y(_20227_));
 sky130_fd_sc_hd__nand2_1 _23128_ (.A(_20227_),
    .B(\inst$top.soc.cpu.x.source__valid ),
    .Y(_20228_));
 sky130_fd_sc_hd__nand2_1 _23130_ (.A(\inst$top.soc.cpu.x.source__valid ),
    .B(net1839),
    .Y(_20230_));
 sky130_fd_sc_hd__nand3_2 _23131_ (.A(_20228_),
    .B(\inst$top.soc.cpu.d.source__valid ),
    .C(_20230_),
    .Y(_20231_));
 sky130_fd_sc_hd__nor2_1 _23132_ (.A(_20138_),
    .B(_20231_),
    .Y(_20232_));
 sky130_fd_sc_hd__nor2_2 _23135_ (.A(net2637),
    .B(net2677),
    .Y(_20235_));
 sky130_fd_sc_hd__inv_2 _23136_ (.A(net2511),
    .Y(_20236_));
 sky130_fd_sc_hd__nor2_1 _23137_ (.A(net2611),
    .B(net2603),
    .Y(_20237_));
 sky130_fd_sc_hd__inv_1 _23138_ (.A(net2496),
    .Y(_20238_));
 sky130_fd_sc_hd__nor3_1 _23139_ (.A(net2591),
    .B(_20236_),
    .C(_20238_),
    .Y(_20239_));
 sky130_fd_sc_hd__inv_1 _23140_ (.A(_20239_),
    .Y(_20240_));
 sky130_fd_sc_hd__xor2_1 _23141_ (.A(\inst$top.soc.cpu.sink__payload$12[100] ),
    .B(net2590),
    .X(_20241_));
 sky130_fd_sc_hd__xor2_1 _23142_ (.A(\inst$top.soc.cpu.sink__payload$12[42] ),
    .B(net2597),
    .X(_20242_));
 sky130_fd_sc_hd__xnor2_1 _23143_ (.A(net2687),
    .B(\inst$top.soc.cpu.sink__payload$12[39] ),
    .Y(_20243_));
 sky130_fd_sc_hd__xnor2_1 _23144_ (.A(net2620),
    .B(\inst$top.soc.cpu.sink__payload$12[40] ),
    .Y(_20244_));
 sky130_fd_sc_hd__nand2_1 _23145_ (.A(_20243_),
    .B(_20244_),
    .Y(_20245_));
 sky130_fd_sc_hd__nor3_1 _23146_ (.A(_20241_),
    .B(_20242_),
    .C(_20245_),
    .Y(_20246_));
 sky130_fd_sc_hd__xnor2_1 _23147_ (.A(net2608),
    .B(\inst$top.soc.cpu.sink__payload$12[41] ),
    .Y(_20247_));
 sky130_fd_sc_hd__and2_0 _23148_ (.A(_20246_),
    .B(_20247_),
    .X(_20248_));
 sky130_fd_sc_hd__nand4_1 _23149_ (.A(_20232_),
    .B(\inst$top.soc.cpu.d.sink__payload.bypass_x ),
    .C(_20240_),
    .D(_20248_),
    .Y(_20249_));
 sky130_fd_sc_hd__nand2_1 _23150_ (.A(_20218_),
    .B(net1192),
    .Y(_20250_));
 sky130_fd_sc_hd__inv_1 _23151_ (.A(_20199_),
    .Y(_20251_));
 sky130_fd_sc_hd__nor2_1 _23152_ (.A(_20250_),
    .B(_20251_),
    .Y(_20252_));
 sky130_fd_sc_hd__inv_1 _23153_ (.A(net1068),
    .Y(_20253_));
 sky130_fd_sc_hd__nand3_2 _23154_ (.A(_20252_),
    .B(_20253_),
    .C(net1018),
    .Y(_20254_));
 sky130_fd_sc_hd__nor2_4 _23155_ (.A(_20224_),
    .B(_20254_),
    .Y(_20255_));
 sky130_fd_sc_hd__inv_1 _23157_ (.A(net1838),
    .Y(_20257_));
 sky130_fd_sc_hd__nand3_2 _23158_ (.A(net874),
    .B(net2539),
    .C(_20257_),
    .Y(_20258_));
 sky130_fd_sc_hd__nand2_1 _23159_ (.A(_20258_),
    .B(\inst$top.soc.cpu.x.source__valid ),
    .Y(_20259_));
 sky130_fd_sc_hd__nand4_2 _23160_ (.A(_20259_),
    .B(\inst$top.soc.cpu.d.sink__payload.rd_we ),
    .C(\inst$top.soc.cpu.d.source__valid ),
    .D(_20248_),
    .Y(_20260_));
 sky130_fd_sc_hd__clkinv_1 _23161_ (.A(net2620),
    .Y(_20261_));
 sky130_fd_sc_hd__nand2_1 _23162_ (.A(\inst$top.soc.cpu.d.sink__payload$6.rd_we ),
    .B(\inst$top.soc.cpu.x.source__valid ),
    .Y(_20262_));
 sky130_fd_sc_hd__inv_2 _23163_ (.A(net2680),
    .Y(_20263_));
 sky130_fd_sc_hd__clkinv_1 _23164_ (.A(net2611),
    .Y(_20264_));
 sky130_fd_sc_hd__o22ai_1 _23165_ (.A1(\inst$top.soc.cpu.sink__payload$18[39] ),
    .A2(net2465),
    .B1(net2460),
    .B2(\inst$top.soc.cpu.sink__payload$18[101] ),
    .Y(_20265_));
 sky130_fd_sc_hd__a211oi_1 _23166_ (.A1(_20261_),
    .A2(\inst$top.soc.cpu.sink__payload$18[100] ),
    .B1(_20262_),
    .C1(_20265_),
    .Y(_20266_));
 sky130_fd_sc_hd__inv_2 _23167_ (.A(\inst$top.soc.cpu.sink__payload$18[101] ),
    .Y(_20267_));
 sky130_fd_sc_hd__o22ai_1 _23168_ (.A1(net2608),
    .A2(_20267_),
    .B1(_20261_),
    .B2(\inst$top.soc.cpu.sink__payload$18[100] ),
    .Y(_20268_));
 sky130_fd_sc_hd__a21oi_1 _23169_ (.A1(net2465),
    .A2(\inst$top.soc.cpu.sink__payload$18[39] ),
    .B1(_20268_),
    .Y(_20269_));
 sky130_fd_sc_hd__nand2_1 _23170_ (.A(\inst$top.soc.cpu.sink__payload$18[103] ),
    .B(net2590),
    .Y(_20270_));
 sky130_fd_sc_hd__inv_1 _23171_ (.A(\inst$top.soc.cpu.sink__payload$18[103] ),
    .Y(_20271_));
 sky130_fd_sc_hd__inv_1 _23172_ (.A(net2590),
    .Y(_20272_));
 sky130_fd_sc_hd__nand2_1 _23173_ (.A(_20271_),
    .B(net2450),
    .Y(_20273_));
 sky130_fd_sc_hd__xor2_1 _23174_ (.A(\inst$top.soc.cpu.sink__payload$18[102] ),
    .B(net2597),
    .X(_20274_));
 sky130_fd_sc_hd__a21oi_1 _23175_ (.A1(_20270_),
    .A2(_20273_),
    .B1(_20274_),
    .Y(_20275_));
 sky130_fd_sc_hd__nand3_1 _23176_ (.A(_20266_),
    .B(_20269_),
    .C(_20275_),
    .Y(_20276_));
 sky130_fd_sc_hd__inv_1 _23177_ (.A(_20276_),
    .Y(_20277_));
 sky130_fd_sc_hd__inv_1 _23178_ (.A(\inst$top.soc.cpu.d.sink__payload$6.bypass_m ),
    .Y(_20278_));
 sky130_fd_sc_hd__nand2_1 _23179_ (.A(_20277_),
    .B(_20278_),
    .Y(_20279_));
 sky130_fd_sc_hd__nand3_1 _23180_ (.A(_20260_),
    .B(_20240_),
    .C(_20279_),
    .Y(_20280_));
 sky130_fd_sc_hd__nand2_1 _23181_ (.A(\inst$top.soc.cpu.sink__payload$6[34] ),
    .B(\inst$top.soc.cpu.sink__payload$6[35] ),
    .Y(_20281_));
 sky130_fd_sc_hd__inv_1 _23182_ (.A(\inst$top.soc.cpu.sink__payload$6[37] ),
    .Y(_20282_));
 sky130_fd_sc_hd__nor2_1 _23183_ (.A(\inst$top.soc.cpu.sink__payload$6[36] ),
    .B(_20282_),
    .Y(_20283_));
 sky130_fd_sc_hd__nand2_1 _23184_ (.A(_20283_),
    .B(net2821),
    .Y(_20284_));
 sky130_fd_sc_hd__nor2_1 _23185_ (.A(_20281_),
    .B(_20284_),
    .Y(_20285_));
 sky130_fd_sc_hd__nor2_1 _23187_ (.A(\inst$top.soc.cpu.sink__payload$6[37] ),
    .B(\inst$top.soc.cpu.sink__payload$6[36] ),
    .Y(_20287_));
 sky130_fd_sc_hd__nor2_1 _23188_ (.A(\inst$top.soc.cpu.sink__payload$6[34] ),
    .B(\inst$top.soc.cpu.sink__payload$6[35] ),
    .Y(_20288_));
 sky130_fd_sc_hd__nand2_1 _23189_ (.A(_20287_),
    .B(_20288_),
    .Y(_20289_));
 sky130_fd_sc_hd__nor2_1 _23190_ (.A(\inst$top.soc.cpu.sink__payload$6[38] ),
    .B(_20289_),
    .Y(_20290_));
 sky130_fd_sc_hd__inv_1 _23191_ (.A(net2821),
    .Y(_20291_));
 sky130_fd_sc_hd__nand2_1 _23192_ (.A(\inst$top.soc.cpu.sink__payload$6[37] ),
    .B(\inst$top.soc.cpu.sink__payload$6[36] ),
    .Y(_20292_));
 sky130_fd_sc_hd__inv_1 _23193_ (.A(_20288_),
    .Y(_20293_));
 sky130_fd_sc_hd__nor3_1 _23194_ (.A(_20291_),
    .B(_20292_),
    .C(_20293_),
    .Y(_20294_));
 sky130_fd_sc_hd__inv_1 _23195_ (.A(_20294_),
    .Y(_20295_));
 sky130_fd_sc_hd__nand3_1 _23196_ (.A(_20283_),
    .B(net2821),
    .C(_20288_),
    .Y(_20296_));
 sky130_fd_sc_hd__nand2_1 _23197_ (.A(_20295_),
    .B(_20296_),
    .Y(_20297_));
 sky130_fd_sc_hd__nor3_1 _23198_ (.A(_20285_),
    .B(_20290_),
    .C(_20297_),
    .Y(_20298_));
 sky130_fd_sc_hd__nand3_1 _23199_ (.A(_20287_),
    .B(\inst$top.soc.cpu.sink__payload$6[34] ),
    .C(\inst$top.soc.cpu.sink__payload$6[35] ),
    .Y(_20299_));
 sky130_fd_sc_hd__nor2_1 _23200_ (.A(net2821),
    .B(_20299_),
    .Y(_20300_));
 sky130_fd_sc_hd__inv_1 _23201_ (.A(\inst$top.soc.cpu.sink__payload$6[35] ),
    .Y(_20301_));
 sky130_fd_sc_hd__nand2_1 _23202_ (.A(_20301_),
    .B(\inst$top.soc.cpu.sink__payload$6[34] ),
    .Y(_20302_));
 sky130_fd_sc_hd__nor2_1 _23203_ (.A(_20302_),
    .B(_20284_),
    .Y(_20303_));
 sky130_fd_sc_hd__inv_1 _23204_ (.A(\inst$top.soc.cpu.sink__payload$6[36] ),
    .Y(_20304_));
 sky130_fd_sc_hd__nand2_1 _23205_ (.A(_20288_),
    .B(_20291_),
    .Y(_20305_));
 sky130_fd_sc_hd__nor2_1 _23206_ (.A(_20304_),
    .B(_20305_),
    .Y(_20306_));
 sky130_fd_sc_hd__nand2_1 _23207_ (.A(_20306_),
    .B(_20282_),
    .Y(_20307_));
 sky130_fd_sc_hd__nor3b_1 _23208_ (.A(_20300_),
    .B(_20303_),
    .C_N(_20307_),
    .Y(_20308_));
 sky130_fd_sc_hd__nor3_1 _23209_ (.A(net2821),
    .B(_20292_),
    .C(_20302_),
    .Y(_20309_));
 sky130_fd_sc_hd__nor4_1 _23210_ (.A(\inst$top.soc.cpu.sink__payload$6[37] ),
    .B(net2821),
    .C(_20304_),
    .D(_20302_),
    .Y(_20310_));
 sky130_fd_sc_hd__nor2_1 _23211_ (.A(_20309_),
    .B(_20310_),
    .Y(_20311_));
 sky130_fd_sc_hd__nand3_1 _23212_ (.A(_20298_),
    .B(_20308_),
    .C(_20311_),
    .Y(_20312_));
 sky130_fd_sc_hd__a21oi_1 _23213_ (.A1(_20312_),
    .A2(_20296_),
    .B1(_20239_),
    .Y(_20313_));
 sky130_fd_sc_hd__nand3_1 _23214_ (.A(_20249_),
    .B(_20280_),
    .C(_20313_),
    .Y(_20314_));
 sky130_fd_sc_hd__xor2_1 _23216_ (.A(net2724),
    .B(\inst$top.soc.cpu.sink__payload$12[40] ),
    .X(_20316_));
 sky130_fd_sc_hd__inv_1 _23217_ (.A(\inst$top.soc.cpu.sink__payload$12[41] ),
    .Y(_20317_));
 sky130_fd_sc_hd__clkinv_1 _23218_ (.A(net2691),
    .Y(_20318_));
 sky130_fd_sc_hd__o22ai_1 _23219_ (.A1(net2703),
    .A2(_20317_),
    .B1(net2445),
    .B2(\inst$top.soc.cpu.sink__payload$12[100] ),
    .Y(_20319_));
 sky130_fd_sc_hd__inv_1 _23220_ (.A(net2698),
    .Y(_20320_));
 sky130_fd_sc_hd__inv_1 _23221_ (.A(\inst$top.soc.cpu.sink__payload$12[39] ),
    .Y(_20321_));
 sky130_fd_sc_hd__nand2_1 _23222_ (.A(_20321_),
    .B(net2767),
    .Y(_20322_));
 sky130_fd_sc_hd__o21ai_0 _23223_ (.A1(\inst$top.soc.cpu.sink__payload$12[42] ),
    .A2(net2432),
    .B1(_20322_),
    .Y(_20323_));
 sky130_fd_sc_hd__clkinv_1 _23224_ (.A(net2711),
    .Y(_20324_));
 sky130_fd_sc_hd__nand2_1 _23225_ (.A(net2445),
    .B(\inst$top.soc.cpu.sink__payload$12[100] ),
    .Y(_20325_));
 sky130_fd_sc_hd__nand2_1 _23226_ (.A(net2432),
    .B(\inst$top.soc.cpu.sink__payload$12[42] ),
    .Y(_20326_));
 sky130_fd_sc_hd__inv_2 _23227_ (.A(net2802),
    .Y(_20327_));
 sky130_fd_sc_hd__nand2_1 _23228_ (.A(net2349),
    .B(\inst$top.soc.cpu.sink__payload$12[39] ),
    .Y(_20328_));
 sky130_fd_sc_hd__o2111ai_1 _23229_ (.A1(\inst$top.soc.cpu.sink__payload$12[41] ),
    .A2(net2417),
    .B1(_20325_),
    .C1(_20326_),
    .D1(_20328_),
    .Y(_20329_));
 sky130_fd_sc_hd__nor4_1 _23230_ (.A(_20316_),
    .B(_20319_),
    .C(_20323_),
    .D(_20329_),
    .Y(_20330_));
 sky130_fd_sc_hd__nand4_2 _23231_ (.A(_20259_),
    .B(\inst$top.soc.cpu.d.sink__payload.rd_we ),
    .C(\inst$top.soc.cpu.d.source__valid ),
    .D(_20330_),
    .Y(_20331_));
 sky130_fd_sc_hd__nor2_1 _23232_ (.A(net2690),
    .B(net2696),
    .Y(_20332_));
 sky130_fd_sc_hd__inv_2 _23233_ (.A(net2729),
    .Y(_20333_));
 sky130_fd_sc_hd__nand4_1 _23234_ (.A(_20332_),
    .B(net2322),
    .C(net2349),
    .D(net2417),
    .Y(_20334_));
 sky130_fd_sc_hd__o22ai_1 _23235_ (.A1(\inst$top.soc.cpu.sink__payload$18[39] ),
    .A2(net2349),
    .B1(net2432),
    .B2(\inst$top.soc.cpu.sink__payload$18[102] ),
    .Y(_20335_));
 sky130_fd_sc_hd__a221oi_1 _23236_ (.A1(net2690),
    .A2(_20271_),
    .B1(net2349),
    .B2(\inst$top.soc.cpu.sink__payload$18[39] ),
    .C1(_20335_),
    .Y(_20336_));
 sky130_fd_sc_hd__o22ai_1 _23237_ (.A1(\inst$top.soc.cpu.sink__payload$18[100] ),
    .A2(net2322),
    .B1(net2417),
    .B2(\inst$top.soc.cpu.sink__payload$18[101] ),
    .Y(_20337_));
 sky130_fd_sc_hd__a211oi_1 _23238_ (.A1(net2322),
    .A2(\inst$top.soc.cpu.sink__payload$18[100] ),
    .B1(_20262_),
    .C1(_20337_),
    .Y(_20338_));
 sky130_fd_sc_hd__o22ai_1 _23240_ (.A1(net2690),
    .A2(_20271_),
    .B1(net2703),
    .B2(_20267_),
    .Y(_20340_));
 sky130_fd_sc_hd__a21oi_1 _23241_ (.A1(net2432),
    .A2(\inst$top.soc.cpu.sink__payload$18[102] ),
    .B1(_20340_),
    .Y(_20341_));
 sky130_fd_sc_hd__nand3_1 _23242_ (.A(_20336_),
    .B(_20338_),
    .C(_20341_),
    .Y(_20342_));
 sky130_fd_sc_hd__inv_1 _23243_ (.A(_20342_),
    .Y(_20343_));
 sky130_fd_sc_hd__nand2_1 _23244_ (.A(_20343_),
    .B(_20278_),
    .Y(_20344_));
 sky130_fd_sc_hd__nand3_1 _23245_ (.A(_20331_),
    .B(_20334_),
    .C(_20344_),
    .Y(_20345_));
 sky130_fd_sc_hd__nand3_1 _23246_ (.A(_20232_),
    .B(\inst$top.soc.cpu.d.sink__payload.bypass_x ),
    .C(_20330_),
    .Y(_20346_));
 sky130_fd_sc_hd__inv_1 _23247_ (.A(_20334_),
    .Y(_20347_));
 sky130_fd_sc_hd__inv_1 _23248_ (.A(_20285_),
    .Y(_20348_));
 sky130_fd_sc_hd__nand2_1 _23249_ (.A(_20311_),
    .B(_20348_),
    .Y(_20349_));
 sky130_fd_sc_hd__nor2_1 _23251_ (.A(_20347_),
    .B(_20349_),
    .Y(_20351_));
 sky130_fd_sc_hd__nand3_1 _23252_ (.A(_20345_),
    .B(_20346_),
    .C(_20351_),
    .Y(_20352_));
 sky130_fd_sc_hd__nor2_1 _23253_ (.A(\inst$top.soc.cpu.sink__payload$6[45] ),
    .B(\inst$top.soc.cpu.sink__payload$6[44] ),
    .Y(_20353_));
 sky130_fd_sc_hd__nor2_1 _23254_ (.A(_20353_),
    .B(_20295_),
    .Y(_20354_));
 sky130_fd_sc_hd__o31ai_1 _23255_ (.A1(\inst$top.soc.cpu.m.source__valid ),
    .A2(\inst$top.soc.cpu.x.source__valid ),
    .A3(\inst$top.soc.cpu.d.source__valid ),
    .B1(_20354_),
    .Y(_20355_));
 sky130_fd_sc_hd__nand3_2 _23256_ (.A(_20314_),
    .B(_20352_),
    .C(_20355_),
    .Y(_20356_));
 sky130_fd_sc_hd__inv_2 _23257_ (.A(_02862_),
    .Y(_20357_));
 sky130_fd_sc_hd__nand4_1 _23258_ (.A(net872),
    .B(net2537),
    .C(net1816),
    .D(_20257_),
    .Y(_20358_));
 sky130_fd_sc_hd__nand2_1 _23259_ (.A(_20358_),
    .B(\inst$top.soc.cpu.x.source__valid ),
    .Y(_20359_));
 sky130_fd_sc_hd__nand2_1 _23260_ (.A(_20359_),
    .B(\inst$top.soc.cpu.f.source__valid ),
    .Y(_20360_));
 sky130_fd_sc_hd__inv_1 _23261_ (.A(\inst$top.soc.cpu.d.sink__payload.fence_i ),
    .Y(_20361_));
 sky130_fd_sc_hd__nor2_1 _23262_ (.A(_20361_),
    .B(_20231_),
    .Y(_20362_));
 sky130_fd_sc_hd__nor2_4 _23263_ (.A(_20360_),
    .B(net837),
    .Y(_20363_));
 sky130_fd_sc_hd__inv_2 _23264_ (.A(_20231_),
    .Y(_20364_));
 sky130_fd_sc_hd__nand2_1 _23265_ (.A(_20364_),
    .B(\inst$top.soc.cpu.d.sink__payload.csr_we ),
    .Y(_20365_));
 sky130_fd_sc_hd__nand3_1 _23266_ (.A(net879),
    .B(\inst$top.soc.cpu.x.source__valid ),
    .C(\inst$top.soc.cpu.d.sink__payload$6.csr_we ),
    .Y(_20366_));
 sky130_fd_sc_hd__nor3_2 _23267_ (.A(\inst$top.soc.cpu.fetch.ibus__cyc ),
    .B(net2931),
    .C(\inst$top.soc.cpu.loadstore.dbus__cyc ),
    .Y(_20367_));
 sky130_fd_sc_hd__nand3_1 _23268_ (.A(_19828_),
    .B(\inst$top.soc.cpu.m.source__valid ),
    .C(\inst$top.soc.cpu.d.sink__payload$16.csr_we ),
    .Y(_20368_));
 sky130_fd_sc_hd__nand4_1 _23269_ (.A(_20365_),
    .B(_20366_),
    .C(net2238),
    .D(_20368_),
    .Y(_20369_));
 sky130_fd_sc_hd__a21oi_2 _23270_ (.A1(_20356_),
    .A2(net792),
    .B1(_20369_),
    .Y(_20370_));
 sky130_fd_sc_hd__nor2_1 _23273_ (.A(_19835_),
    .B(_19839_),
    .Y(_00129_));
 sky130_fd_sc_hd__nor2_2 _23274_ (.A(_19840_),
    .B(_19832_),
    .Y(_00156_));
 sky130_fd_sc_hd__nor2_4 _23275_ (.A(_19845_),
    .B(_19839_),
    .Y(_00136_));
 sky130_fd_sc_hd__nand2_1 _23277_ (.A(net2847),
    .B(\inst$top.soc.cpu.d.sink__payload.csr_clear ),
    .Y(_20373_));
 sky130_fd_sc_hd__xor2_1 _23278_ (.A(_20373_),
    .B(net1692),
    .X(_03085_));
 sky130_fd_sc_hd__inv_2 _23279_ (.A(_03085_),
    .Y(_03089_));
 sky130_fd_sc_hd__nand2_1 _23280_ (.A(net2551),
    .B(\inst$top.soc.cpu.gprf.mem_rp2__data[0] ),
    .Y(_20374_));
 sky130_fd_sc_hd__nand2_1 _23281_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_raw ),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[0] ),
    .Y(_20375_));
 sky130_fd_sc_hd__nand2_1 _23282_ (.A(_20374_),
    .B(_20375_),
    .Y(_20376_));
 sky130_fd_sc_hd__or2_2 _23283_ (.A(\inst$top.soc.cpu.sink__payload$12[109] ),
    .B(net1986),
    .X(_20377_));
 sky130_fd_sc_hd__o21ai_2 _23284_ (.A1(_20376_),
    .A2(net1827),
    .B1(_20377_),
    .Y(_20378_));
 sky130_fd_sc_hd__clkinv_1 _23288_ (.A(net2843),
    .Y(_20381_));
 sky130_fd_sc_hd__inv_1 _23290_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa_x_select ),
    .Y(_20383_));
 sky130_fd_sc_hd__inv_1 _23292_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[0] ),
    .Y(_20385_));
 sky130_fd_sc_hd__inv_1 _23293_ (.A(net2892),
    .Y(_20386_));
 sky130_fd_sc_hd__inv_1 _23295_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.mode.x_data[0] ),
    .Y(_20388_));
 sky130_fd_sc_hd__inv_1 _23297_ (.A(net2897),
    .Y(_20390_));
 sky130_fd_sc_hd__inv_1 _23298_ (.A(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[0] ),
    .Y(_20391_));
 sky130_fd_sc_hd__nand2_1 _23299_ (.A(net2893),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[0] ),
    .Y(_20392_));
 sky130_fd_sc_hd__o21ai_0 _23300_ (.A1(_20390_),
    .A2(_20391_),
    .B1(_20392_),
    .Y(_20393_));
 sky130_fd_sc_hd__a21oi_1 _23301_ (.A1(net2915),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[0] ),
    .B1(_20393_),
    .Y(_20394_));
 sky130_fd_sc_hd__o221ai_1 _23302_ (.A1(net2213),
    .A2(_20385_),
    .B1(net2210),
    .B2(_20388_),
    .C1(_20394_),
    .Y(_20395_));
 sky130_fd_sc_hd__nand2_1 _23303_ (.A(_20395_),
    .B(\inst$top.soc.cpu.csrf.bank_300_x_select ),
    .Y(_20396_));
 sky130_fd_sc_hd__nand2_1 _23304_ (.A(_20396_),
    .B(net2845),
    .Y(_20397_));
 sky130_fd_sc_hd__inv_1 _23305_ (.A(_20397_),
    .Y(_20398_));
 sky130_fd_sc_hd__a21oi_1 _23306_ (.A1(net2215),
    .A2(net1682),
    .B1(_20398_),
    .Y(_03084_));
 sky130_fd_sc_hd__inv_2 _23307_ (.A(_03084_),
    .Y(_03088_));
 sky130_fd_sc_hd__inv_2 _23308_ (.A(\inst$top.soc.cpu.divider.quotient[0] ),
    .Y(_02846_));
 sky130_fd_sc_hd__inv_2 _23309_ (.A(\inst$top.soc.cpu.divider.remainder[0] ),
    .Y(_02853_));
 sky130_fd_sc_hd__inv_2 _23310_ (.A(\inst$top.soc.cpu.d.sink__payload$16.load ),
    .Y(_20399_));
 sky130_fd_sc_hd__inv_1 _23313_ (.A(\inst$top.soc.cpu.sink__payload$24[39] ),
    .Y(_20402_));
 sky130_fd_sc_hd__nor3_1 _23314_ (.A(\inst$top.soc.cpu.sink__payload$24[38] ),
    .B(\inst$top.soc.cpu.sink__payload$24[40] ),
    .C(_20402_),
    .Y(_20403_));
 sky130_fd_sc_hd__inv_1 _23317_ (.A(\inst$top.soc.cpu.sink__payload$24[82] ),
    .Y(_20406_));
 sky130_fd_sc_hd__nand2_1 _23318_ (.A(net2823),
    .B(\inst$top.soc.cpu.sink__payload$24[98] ),
    .Y(_20407_));
 sky130_fd_sc_hd__o21ai_0 _23319_ (.A1(net2823),
    .A2(_20406_),
    .B1(_20407_),
    .Y(_20408_));
 sky130_fd_sc_hd__inv_1 _23320_ (.A(\inst$top.soc.cpu.sink__payload$24[41] ),
    .Y(_20409_));
 sky130_fd_sc_hd__nor2_1 _23321_ (.A(\inst$top.soc.cpu.sink__payload$24[38] ),
    .B(\inst$top.soc.cpu.sink__payload$24[39] ),
    .Y(_20410_));
 sky130_fd_sc_hd__inv_1 _23322_ (.A(_20410_),
    .Y(_20411_));
 sky130_fd_sc_hd__nor2_1 _23323_ (.A(_20409_),
    .B(_20411_),
    .Y(_20412_));
 sky130_fd_sc_hd__clkinv_1 _23324_ (.A(net2823),
    .Y(_20413_));
 sky130_fd_sc_hd__nand2_1 _23325_ (.A(_20413_),
    .B(\inst$top.soc.cpu.sink__payload$24[74] ),
    .Y(_20414_));
 sky130_fd_sc_hd__nand2_1 _23327_ (.A(\inst$top.soc.cpu.sink__payload$24[90] ),
    .B(net2824),
    .Y(_20416_));
 sky130_fd_sc_hd__inv_1 _23328_ (.A(\inst$top.soc.cpu.sink__payload$24[38] ),
    .Y(_20417_));
 sky130_fd_sc_hd__a21oi_1 _23329_ (.A1(_20417_),
    .A2(\inst$top.soc.cpu.sink__payload$24[41] ),
    .B1(\inst$top.soc.cpu.sink__payload$24[39] ),
    .Y(_20418_));
 sky130_fd_sc_hd__inv_1 _23330_ (.A(_20418_),
    .Y(_20419_));
 sky130_fd_sc_hd__a21oi_1 _23331_ (.A1(_20414_),
    .A2(_20416_),
    .B1(_20419_),
    .Y(_20420_));
 sky130_fd_sc_hd__a221oi_1 _23332_ (.A1(\inst$top.soc.cpu.sink__payload$24[74] ),
    .A2(net1983),
    .B1(_20408_),
    .B2(_20412_),
    .C1(_20420_),
    .Y(_20421_));
 sky130_fd_sc_hd__clkinv_1 _23333_ (.A(net2827),
    .Y(_20422_));
 sky130_fd_sc_hd__nand2_1 _23336_ (.A(_20409_),
    .B(net2197),
    .Y(_20425_));
 sky130_fd_sc_hd__o211ai_1 _23337_ (.A1(\inst$top.soc.cpu.multiplier.w_result[0] ),
    .A2(net2197),
    .B1(net2202),
    .C1(_20425_),
    .Y(_20426_));
 sky130_fd_sc_hd__o21a_1 _23338_ (.A1(net2201),
    .A2(_20421_),
    .B1(_20426_),
    .X(_20427_));
 sky130_fd_sc_hd__inv_2 _23339_ (.A(_20427_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[0] ));
 sky130_fd_sc_hd__xor2_1 _23340_ (.A(_20373_),
    .B(net1706),
    .X(_03092_));
 sky130_fd_sc_hd__inv_2 _23341_ (.A(_03092_),
    .Y(_03096_));
 sky130_fd_sc_hd__inv_1 _23347_ (.A(\inst$top.soc.cpu.csrf.bank_300_x_select ),
    .Y(_20432_));
 sky130_fd_sc_hd__inv_1 _23348_ (.A(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[1] ),
    .Y(_20433_));
 sky130_fd_sc_hd__nand2_1 _23349_ (.A(net2893),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[1] ),
    .Y(_20434_));
 sky130_fd_sc_hd__o21ai_0 _23350_ (.A1(_20390_),
    .A2(_20433_),
    .B1(_20434_),
    .Y(_20435_));
 sky130_fd_sc_hd__inv_1 _23351_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[1] ),
    .Y(_20436_));
 sky130_fd_sc_hd__inv_1 _23353_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.mode.x_data[1] ),
    .Y(_20438_));
 sky130_fd_sc_hd__o22ai_1 _23354_ (.A1(net2213),
    .A2(_20436_),
    .B1(net2210),
    .B2(_20438_),
    .Y(_20439_));
 sky130_fd_sc_hd__a211oi_2 _23355_ (.A1(net2915),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[1] ),
    .B1(_20435_),
    .C1(_20439_),
    .Y(_20440_));
 sky130_fd_sc_hd__o21ai_0 _23356_ (.A1(_20432_),
    .A2(_20440_),
    .B1(net2845),
    .Y(_20441_));
 sky130_fd_sc_hd__o21ai_1 _23357_ (.A1(net2848),
    .A2(net1385),
    .B1(_20441_),
    .Y(_03095_));
 sky130_fd_sc_hd__inv_1 _23358_ (.A(\inst$top.soc.cpu.sink__payload$24[83] ),
    .Y(_20442_));
 sky130_fd_sc_hd__nand2_1 _23359_ (.A(net2823),
    .B(\inst$top.soc.cpu.sink__payload$24[99] ),
    .Y(_20443_));
 sky130_fd_sc_hd__o21ai_0 _23360_ (.A1(net2823),
    .A2(_20442_),
    .B1(_20443_),
    .Y(_20444_));
 sky130_fd_sc_hd__a32oi_1 _23361_ (.A1(_20418_),
    .A2(net2823),
    .A3(\inst$top.soc.cpu.sink__payload$24[91] ),
    .B1(_20412_),
    .B2(_20444_),
    .Y(_20445_));
 sky130_fd_sc_hd__inv_1 _23363_ (.A(net1982),
    .Y(_20447_));
 sky130_fd_sc_hd__o21ai_0 _23364_ (.A1(net2822),
    .A2(_20419_),
    .B1(_20447_),
    .Y(_20448_));
 sky130_fd_sc_hd__nand2_1 _23365_ (.A(_20448_),
    .B(\inst$top.soc.cpu.sink__payload$24[75] ),
    .Y(_20449_));
 sky130_fd_sc_hd__nand2_1 _23366_ (.A(_20445_),
    .B(_20449_),
    .Y(_20450_));
 sky130_fd_sc_hd__nand2_1 _23368_ (.A(net2197),
    .B(_20413_),
    .Y(_20452_));
 sky130_fd_sc_hd__o211a_1 _23369_ (.A1(\inst$top.soc.cpu.multiplier.w_result[1] ),
    .A2(net2197),
    .B1(net2201),
    .C1(_20452_),
    .X(_20453_));
 sky130_fd_sc_hd__a21oi_1 _23370_ (.A1(_20450_),
    .A2(\inst$top.soc.cpu.d.sink__payload$16.load ),
    .B1(_20453_),
    .Y(_20454_));
 sky130_fd_sc_hd__inv_2 _23371_ (.A(_20454_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[1] ));
 sky130_fd_sc_hd__inv_1 _23372_ (.A(\inst$top.soc.cpu.gprf.mem_rp1__data[2] ),
    .Y(_20455_));
 sky130_fd_sc_hd__nand2_1 _23373_ (.A(net2549),
    .B(_20455_),
    .Y(_20456_));
 sky130_fd_sc_hd__inv_1 _23374_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[2] ),
    .Y(_20457_));
 sky130_fd_sc_hd__nand2_1 _23375_ (.A(_20457_),
    .B(net2886),
    .Y(_20458_));
 sky130_fd_sc_hd__nand3_1 _23376_ (.A(_20456_),
    .B(_20458_),
    .C(_19879_),
    .Y(_20459_));
 sky130_fd_sc_hd__nand2_1 _23377_ (.A(_20117_),
    .B(\inst$top.soc.cpu.sink__payload$12[103] ),
    .Y(_20460_));
 sky130_fd_sc_hd__nand3_1 _23378_ (.A(_20459_),
    .B(_19870_),
    .C(_20460_),
    .Y(_20461_));
 sky130_fd_sc_hd__inv_1 _23379_ (.A(\inst$top.soc.cpu.sink__payload$12[2] ),
    .Y(_20462_));
 sky130_fd_sc_hd__a21oi_1 _23380_ (.A1(_20462_),
    .A2(\inst$top.soc.cpu.d.sink__payload.auipc ),
    .B1(\inst$top.soc.cpu.d.sink__payload.lui ),
    .Y(_20463_));
 sky130_fd_sc_hd__nand2_1 _23381_ (.A(_20461_),
    .B(_20463_),
    .Y(_20464_));
 sky130_fd_sc_hd__xor2_1 _23382_ (.A(_20373_),
    .B(net1366),
    .X(_03099_));
 sky130_fd_sc_hd__inv_2 _23383_ (.A(_03099_),
    .Y(_03103_));
 sky130_fd_sc_hd__clkinv_1 _23384_ (.A(net1386),
    .Y(_20465_));
 sky130_fd_sc_hd__inv_1 _23391_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[2] ),
    .Y(_20471_));
 sky130_fd_sc_hd__inv_1 _23392_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[0] ),
    .Y(_20472_));
 sky130_fd_sc_hd__o22ai_1 _23393_ (.A1(net2211),
    .A2(_20471_),
    .B1(net2210),
    .B2(_20472_),
    .Y(_20473_));
 sky130_fd_sc_hd__a221oi_1 _23394_ (.A1(net2897),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[2] ),
    .B1(net2908),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[0] ),
    .C1(_20473_),
    .Y(_20474_));
 sky130_fd_sc_hd__nand2_1 _23396_ (.A(net2893),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[2] ),
    .Y(_20476_));
 sky130_fd_sc_hd__nand2_1 _23398_ (.A(net2912),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[2] ),
    .Y(_20478_));
 sky130_fd_sc_hd__nand3_1 _23399_ (.A(_20474_),
    .B(_20476_),
    .C(_20478_),
    .Y(_20479_));
 sky130_fd_sc_hd__nand2_1 _23400_ (.A(net2845),
    .B(\inst$top.soc.cpu.csrf.bank_300_x_select ),
    .Y(_20480_));
 sky130_fd_sc_hd__inv_1 _23401_ (.A(_20480_),
    .Y(_20481_));
 sky130_fd_sc_hd__nand2_1 _23403_ (.A(_20479_),
    .B(net1980),
    .Y(_20483_));
 sky130_fd_sc_hd__o21ai_1 _23404_ (.A1(net2847),
    .A2(net1182),
    .B1(_20483_),
    .Y(_03098_));
 sky130_fd_sc_hd__inv_2 _23405_ (.A(_03098_),
    .Y(_03102_));
 sky130_fd_sc_hd__nor2_1 _23406_ (.A(net2822),
    .B(\inst$top.soc.cpu.sink__payload$24[76] ),
    .Y(_20484_));
 sky130_fd_sc_hd__nor2_1 _23407_ (.A(\inst$top.soc.cpu.sink__payload$24[92] ),
    .B(_20413_),
    .Y(_20485_));
 sky130_fd_sc_hd__nand2_1 _23409_ (.A(net1982),
    .B(\inst$top.soc.cpu.sink__payload$24[76] ),
    .Y(_20487_));
 sky130_fd_sc_hd__inv_1 _23410_ (.A(\inst$top.soc.cpu.sink__payload$24[84] ),
    .Y(_20488_));
 sky130_fd_sc_hd__nand2_1 _23411_ (.A(net2824),
    .B(\inst$top.soc.cpu.sink__payload$24[100] ),
    .Y(_20489_));
 sky130_fd_sc_hd__o21ai_0 _23412_ (.A1(net2822),
    .A2(_20488_),
    .B1(_20489_),
    .Y(_20490_));
 sky130_fd_sc_hd__nand2_1 _23413_ (.A(_20412_),
    .B(_20490_),
    .Y(_20491_));
 sky130_fd_sc_hd__o311ai_0 _23414_ (.A1(_20484_),
    .A2(_20485_),
    .A3(_20419_),
    .B1(_20487_),
    .C1(_20491_),
    .Y(_20492_));
 sky130_fd_sc_hd__nor2_1 _23416_ (.A(net2825),
    .B(\inst$top.soc.cpu.sink__payload$24[43] ),
    .Y(_20494_));
 sky130_fd_sc_hd__nor2_1 _23417_ (.A(\inst$top.soc.cpu.multiplier.w_result[2] ),
    .B(net2196),
    .Y(_20495_));
 sky130_fd_sc_hd__nor2_1 _23418_ (.A(_20494_),
    .B(_20495_),
    .Y(_20496_));
 sky130_fd_sc_hd__mux2i_1 _23419_ (.A0(_20492_),
    .A1(_20496_),
    .S(net2201),
    .Y(_20497_));
 sky130_fd_sc_hd__inv_2 _23420_ (.A(_20497_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[2] ));
 sky130_fd_sc_hd__inv_2 _23421_ (.A(_20373_),
    .Y(_20498_));
 sky130_fd_sc_hd__nand2_1 _23423_ (.A(net2549),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[3] ),
    .Y(_20500_));
 sky130_fd_sc_hd__nand2_1 _23424_ (.A(net2887),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[3] ),
    .Y(_20501_));
 sky130_fd_sc_hd__nand3_1 _23425_ (.A(_20500_),
    .B(_19879_),
    .C(_20501_),
    .Y(_20502_));
 sky130_fd_sc_hd__o211ai_1 _23426_ (.A1(\inst$top.soc.cpu.sink__payload$12[104] ),
    .A2(_19879_),
    .B1(_19878_),
    .C1(_20502_),
    .Y(_20503_));
 sky130_fd_sc_hd__nand2_1 _23427_ (.A(_19871_),
    .B(\inst$top.soc.cpu.sink__payload$12[3] ),
    .Y(_20504_));
 sky130_fd_sc_hd__nand2_2 _23428_ (.A(_20503_),
    .B(_20504_),
    .Y(_20505_));
 sky130_fd_sc_hd__xor2_1 _23429_ (.A(net1979),
    .B(net1361),
    .X(_03106_));
 sky130_fd_sc_hd__inv_2 _23430_ (.A(_03106_),
    .Y(_03110_));
 sky130_fd_sc_hd__inv_1 _23431_ (.A(net1393),
    .Y(_20506_));
 sky130_fd_sc_hd__clkinv_1 _23435_ (.A(net2905),
    .Y(_20509_));
 sky130_fd_sc_hd__inv_1 _23436_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.msip.x_data ),
    .Y(_20510_));
 sky130_fd_sc_hd__nand2_1 _23437_ (.A(net2896),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[3] ),
    .Y(_20511_));
 sky130_fd_sc_hd__inv_1 _23438_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[1] ),
    .Y(_20512_));
 sky130_fd_sc_hd__nand2_1 _23440_ (.A(net2897),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[3] ),
    .Y(_20514_));
 sky130_fd_sc_hd__nand2_1 _23442_ (.A(net2908),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[1] ),
    .Y(_20516_));
 sky130_fd_sc_hd__inv_1 _23443_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[3] ),
    .Y(_20517_));
 sky130_fd_sc_hd__nand2_1 _23444_ (.A(\inst$top.soc.cpu.exception.csr_bank.mstatus_x_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.mstatus.mie.x_data ),
    .Y(_20518_));
 sky130_fd_sc_hd__o21ai_0 _23445_ (.A1(net2211),
    .A2(_20517_),
    .B1(_20518_),
    .Y(_20519_));
 sky130_fd_sc_hd__a21oi_1 _23446_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mie_x_select ),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mie.msie.x_data ),
    .B1(_20519_),
    .Y(_20520_));
 sky130_fd_sc_hd__o2111ai_1 _23447_ (.A1(net2210),
    .A2(_20512_),
    .B1(_20514_),
    .C1(_20516_),
    .D1(_20520_),
    .Y(_20521_));
 sky130_fd_sc_hd__a21oi_1 _23448_ (.A1(net2915),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[3] ),
    .B1(_20521_),
    .Y(_20522_));
 sky130_fd_sc_hd__o211ai_1 _23449_ (.A1(_20509_),
    .A2(_20510_),
    .B1(_20511_),
    .C1(_20522_),
    .Y(_20523_));
 sky130_fd_sc_hd__nand2_1 _23450_ (.A(_20523_),
    .B(net1980),
    .Y(_20524_));
 sky130_fd_sc_hd__o21ai_1 _23451_ (.A1(net2847),
    .A2(net1174),
    .B1(_20524_),
    .Y(_03105_));
 sky130_fd_sc_hd__inv_2 _23452_ (.A(_03105_),
    .Y(_03109_));
 sky130_fd_sc_hd__nor2_1 _23453_ (.A(net2822),
    .B(\inst$top.soc.cpu.sink__payload$24[77] ),
    .Y(_20525_));
 sky130_fd_sc_hd__nor2_1 _23454_ (.A(\inst$top.soc.cpu.sink__payload$24[93] ),
    .B(_20413_),
    .Y(_20526_));
 sky130_fd_sc_hd__nand2_1 _23455_ (.A(_20413_),
    .B(\inst$top.soc.cpu.sink__payload$24[85] ),
    .Y(_20527_));
 sky130_fd_sc_hd__nand2_1 _23456_ (.A(net2822),
    .B(\inst$top.soc.cpu.sink__payload$24[101] ),
    .Y(_20528_));
 sky130_fd_sc_hd__nand2_1 _23457_ (.A(_20527_),
    .B(_20528_),
    .Y(_20529_));
 sky130_fd_sc_hd__nand2_1 _23458_ (.A(_20412_),
    .B(_20529_),
    .Y(_20530_));
 sky130_fd_sc_hd__nand2_1 _23459_ (.A(net1982),
    .B(\inst$top.soc.cpu.sink__payload$24[77] ),
    .Y(_20531_));
 sky130_fd_sc_hd__o311ai_0 _23460_ (.A1(_20525_),
    .A2(_20526_),
    .A3(_20419_),
    .B1(_20530_),
    .C1(_20531_),
    .Y(_20532_));
 sky130_fd_sc_hd__nor2_1 _23461_ (.A(net2825),
    .B(\inst$top.soc.cpu.sink__payload$24[44] ),
    .Y(_20533_));
 sky130_fd_sc_hd__nor2_1 _23462_ (.A(\inst$top.soc.cpu.multiplier.w_result[3] ),
    .B(net2196),
    .Y(_20534_));
 sky130_fd_sc_hd__nor2_1 _23463_ (.A(_20533_),
    .B(_20534_),
    .Y(_20535_));
 sky130_fd_sc_hd__mux2i_1 _23465_ (.A0(_20532_),
    .A1(_20535_),
    .S(net2203),
    .Y(_20537_));
 sky130_fd_sc_hd__inv_2 _23466_ (.A(_20537_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[3] ));
 sky130_fd_sc_hd__nand2_1 _23467_ (.A(net2546),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[4] ),
    .Y(_20538_));
 sky130_fd_sc_hd__nand2_1 _23468_ (.A(net2886),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[4] ),
    .Y(_20539_));
 sky130_fd_sc_hd__nand3_1 _23469_ (.A(_20538_),
    .B(_19879_),
    .C(_20539_),
    .Y(_20540_));
 sky130_fd_sc_hd__o211ai_1 _23470_ (.A1(\inst$top.soc.cpu.sink__payload$12[105] ),
    .A2(_19879_),
    .B1(_19878_),
    .C1(_20540_),
    .Y(_20541_));
 sky130_fd_sc_hd__nand2_1 _23471_ (.A(_19871_),
    .B(\inst$top.soc.cpu.sink__payload$12[4] ),
    .Y(_20542_));
 sky130_fd_sc_hd__nand2_1 _23472_ (.A(_20541_),
    .B(_20542_),
    .Y(_20543_));
 sky130_fd_sc_hd__xor2_1 _23473_ (.A(net1979),
    .B(net1356),
    .X(_03115_));
 sky130_fd_sc_hd__inv_2 _23474_ (.A(_03115_),
    .Y(_03119_));
 sky130_fd_sc_hd__inv_1 _23479_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[4] ),
    .Y(_20547_));
 sky130_fd_sc_hd__inv_1 _23480_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[2] ),
    .Y(_20548_));
 sky130_fd_sc_hd__o22ai_1 _23481_ (.A1(net2211),
    .A2(_20547_),
    .B1(net2210),
    .B2(_20548_),
    .Y(_20549_));
 sky130_fd_sc_hd__a221oi_1 _23482_ (.A1(net2897),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[4] ),
    .B1(net2908),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[2] ),
    .C1(_20549_),
    .Y(_20550_));
 sky130_fd_sc_hd__nand2_1 _23483_ (.A(net2893),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[4] ),
    .Y(_20551_));
 sky130_fd_sc_hd__nand2_1 _23484_ (.A(net2912),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[4] ),
    .Y(_20552_));
 sky130_fd_sc_hd__nand3_1 _23485_ (.A(_20550_),
    .B(_20551_),
    .C(_20552_),
    .Y(_20553_));
 sky130_fd_sc_hd__nand2_1 _23486_ (.A(_20553_),
    .B(net1980),
    .Y(_20554_));
 sky130_fd_sc_hd__o21ai_1 _23487_ (.A1(net2847),
    .A2(net1197),
    .B1(_20554_),
    .Y(_03114_));
 sky130_fd_sc_hd__inv_2 _23488_ (.A(_03114_),
    .Y(_03118_));
 sky130_fd_sc_hd__nand2_1 _23489_ (.A(_20448_),
    .B(\inst$top.soc.cpu.sink__payload$24[78] ),
    .Y(_20555_));
 sky130_fd_sc_hd__inv_1 _23490_ (.A(\inst$top.soc.cpu.sink__payload$24[86] ),
    .Y(_20556_));
 sky130_fd_sc_hd__nand2_1 _23491_ (.A(net2822),
    .B(\inst$top.soc.cpu.sink__payload$24[102] ),
    .Y(_20557_));
 sky130_fd_sc_hd__o21ai_0 _23492_ (.A1(net2822),
    .A2(_20556_),
    .B1(_20557_),
    .Y(_20558_));
 sky130_fd_sc_hd__nand2_1 _23493_ (.A(_20412_),
    .B(_20558_),
    .Y(_20559_));
 sky130_fd_sc_hd__nand3_1 _23494_ (.A(_20418_),
    .B(net2824),
    .C(\inst$top.soc.cpu.sink__payload$24[94] ),
    .Y(_20560_));
 sky130_fd_sc_hd__nand3_1 _23495_ (.A(_20555_),
    .B(_20559_),
    .C(_20560_),
    .Y(_20561_));
 sky130_fd_sc_hd__nor2_1 _23496_ (.A(net2825),
    .B(\inst$top.soc.cpu.sink__payload$24[45] ),
    .Y(_20562_));
 sky130_fd_sc_hd__nor2_1 _23497_ (.A(\inst$top.soc.cpu.multiplier.w_result[4] ),
    .B(net2196),
    .Y(_20563_));
 sky130_fd_sc_hd__nor2_1 _23498_ (.A(_20562_),
    .B(_20563_),
    .Y(_20564_));
 sky130_fd_sc_hd__mux2i_1 _23499_ (.A0(_20561_),
    .A1(_20564_),
    .S(net2201),
    .Y(_20565_));
 sky130_fd_sc_hd__inv_2 _23500_ (.A(_20565_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[4] ));
 sky130_fd_sc_hd__inv_1 _23501_ (.A(\inst$top.soc.cpu.sink__payload$12[5] ),
    .Y(_20566_));
 sky130_fd_sc_hd__nand2_1 _23502_ (.A(net2546),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[5] ),
    .Y(_20567_));
 sky130_fd_sc_hd__nand2_1 _23503_ (.A(net2886),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[5] ),
    .Y(_20568_));
 sky130_fd_sc_hd__nand2_1 _23504_ (.A(_20567_),
    .B(_20568_),
    .Y(_20569_));
 sky130_fd_sc_hd__nand2_1 _23505_ (.A(net1828),
    .B(_20569_),
    .Y(_20570_));
 sky130_fd_sc_hd__o21ai_2 _23506_ (.A1(_20566_),
    .A2(net1832),
    .B1(_20570_),
    .Y(_20571_));
 sky130_fd_sc_hd__xor2_1 _23507_ (.A(net1979),
    .B(net1351),
    .X(_03122_));
 sky130_fd_sc_hd__inv_2 _23508_ (.A(_03122_),
    .Y(_03126_));
 sky130_fd_sc_hd__inv_2 _23509_ (.A(net1395),
    .Y(_20572_));
 sky130_fd_sc_hd__inv_1 _23512_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[5] ),
    .Y(_20574_));
 sky130_fd_sc_hd__inv_1 _23513_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[3] ),
    .Y(_20575_));
 sky130_fd_sc_hd__o22ai_1 _23514_ (.A1(net2212),
    .A2(_20574_),
    .B1(net2209),
    .B2(_20575_),
    .Y(_20576_));
 sky130_fd_sc_hd__a221oi_1 _23515_ (.A1(net2898),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[5] ),
    .B1(net2910),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[3] ),
    .C1(_20576_),
    .Y(_20577_));
 sky130_fd_sc_hd__nand2_1 _23516_ (.A(net2895),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[5] ),
    .Y(_20578_));
 sky130_fd_sc_hd__nand2_1 _23517_ (.A(net2914),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[5] ),
    .Y(_20579_));
 sky130_fd_sc_hd__nand3_1 _23518_ (.A(_20577_),
    .B(_20578_),
    .C(_20579_),
    .Y(_20580_));
 sky130_fd_sc_hd__nand2_1 _23519_ (.A(_20580_),
    .B(net1980),
    .Y(_20581_));
 sky130_fd_sc_hd__o21ai_1 _23520_ (.A1(net2847),
    .A2(net1172),
    .B1(_20581_),
    .Y(_03121_));
 sky130_fd_sc_hd__inv_2 _23521_ (.A(_03121_),
    .Y(_03125_));
 sky130_fd_sc_hd__nor2_1 _23522_ (.A(net2824),
    .B(\inst$top.soc.cpu.sink__payload$24[79] ),
    .Y(_20582_));
 sky130_fd_sc_hd__nor2_1 _23523_ (.A(\inst$top.soc.cpu.sink__payload$24[95] ),
    .B(_20413_),
    .Y(_20583_));
 sky130_fd_sc_hd__nand2_1 _23524_ (.A(net1983),
    .B(\inst$top.soc.cpu.sink__payload$24[79] ),
    .Y(_20584_));
 sky130_fd_sc_hd__inv_1 _23525_ (.A(\inst$top.soc.cpu.sink__payload$24[87] ),
    .Y(_20585_));
 sky130_fd_sc_hd__nand2_1 _23526_ (.A(net2823),
    .B(\inst$top.soc.cpu.sink__payload$24[103] ),
    .Y(_20586_));
 sky130_fd_sc_hd__o21ai_0 _23527_ (.A1(net2823),
    .A2(_20585_),
    .B1(_20586_),
    .Y(_20587_));
 sky130_fd_sc_hd__nand2_1 _23528_ (.A(_20412_),
    .B(_20587_),
    .Y(_20588_));
 sky130_fd_sc_hd__o311ai_0 _23529_ (.A1(_20582_),
    .A2(_20583_),
    .A3(_20419_),
    .B1(_20584_),
    .C1(_20588_),
    .Y(_20589_));
 sky130_fd_sc_hd__nor2_1 _23530_ (.A(net2826),
    .B(\inst$top.soc.cpu.sink__payload$24[46] ),
    .Y(_20590_));
 sky130_fd_sc_hd__nor2_1 _23531_ (.A(\inst$top.soc.cpu.multiplier.w_result[5] ),
    .B(net2196),
    .Y(_20591_));
 sky130_fd_sc_hd__nor2_1 _23532_ (.A(_20590_),
    .B(_20591_),
    .Y(_20592_));
 sky130_fd_sc_hd__mux2i_1 _23533_ (.A0(_20589_),
    .A1(_20592_),
    .S(net2202),
    .Y(_20593_));
 sky130_fd_sc_hd__inv_2 _23534_ (.A(_20593_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[5] ));
 sky130_fd_sc_hd__clkinv_1 _23535_ (.A(\inst$top.soc.cpu.sink__payload$12[6] ),
    .Y(_20594_));
 sky130_fd_sc_hd__nand2_1 _23536_ (.A(net2549),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[6] ),
    .Y(_20595_));
 sky130_fd_sc_hd__nand2_1 _23537_ (.A(net2888),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[6] ),
    .Y(_20596_));
 sky130_fd_sc_hd__nand2_1 _23538_ (.A(_20595_),
    .B(_20596_),
    .Y(_20597_));
 sky130_fd_sc_hd__nand2_1 _23539_ (.A(net1829),
    .B(_20597_),
    .Y(_20598_));
 sky130_fd_sc_hd__o21ai_1 _23540_ (.A1(_20594_),
    .A2(net1832),
    .B1(_20598_),
    .Y(_20599_));
 sky130_fd_sc_hd__xor2_1 _23542_ (.A(net1979),
    .B(net1350),
    .X(_03129_));
 sky130_fd_sc_hd__inv_2 _23543_ (.A(_03129_),
    .Y(_03133_));
 sky130_fd_sc_hd__inv_2 _23544_ (.A(net1397),
    .Y(_20601_));
 sky130_fd_sc_hd__inv_1 _23546_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[6] ),
    .Y(_20602_));
 sky130_fd_sc_hd__inv_1 _23547_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[4] ),
    .Y(_20603_));
 sky130_fd_sc_hd__o22ai_1 _23548_ (.A1(net2211),
    .A2(_20602_),
    .B1(net2210),
    .B2(_20603_),
    .Y(_20604_));
 sky130_fd_sc_hd__a221oi_1 _23549_ (.A1(net2897),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[6] ),
    .B1(net2908),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[4] ),
    .C1(_20604_),
    .Y(_20605_));
 sky130_fd_sc_hd__nand2_1 _23550_ (.A(net2912),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[6] ),
    .Y(_20606_));
 sky130_fd_sc_hd__nand2_1 _23552_ (.A(net2893),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[6] ),
    .Y(_20608_));
 sky130_fd_sc_hd__nand3_1 _23553_ (.A(_20605_),
    .B(_20606_),
    .C(_20608_),
    .Y(_20609_));
 sky130_fd_sc_hd__nand2_1 _23554_ (.A(_20609_),
    .B(net1980),
    .Y(_20610_));
 sky130_fd_sc_hd__o21ai_1 _23555_ (.A1(net2848),
    .A2(net1166),
    .B1(_20610_),
    .Y(_03128_));
 sky130_fd_sc_hd__inv_2 _23556_ (.A(_03128_),
    .Y(_03132_));
 sky130_fd_sc_hd__nor2_1 _23557_ (.A(net2823),
    .B(\inst$top.soc.cpu.sink__payload$24[80] ),
    .Y(_20611_));
 sky130_fd_sc_hd__nor2_1 _23558_ (.A(\inst$top.soc.cpu.sink__payload$24[96] ),
    .B(_20413_),
    .Y(_20612_));
 sky130_fd_sc_hd__nand2_1 _23559_ (.A(net1983),
    .B(\inst$top.soc.cpu.sink__payload$24[80] ),
    .Y(_20613_));
 sky130_fd_sc_hd__nand2_1 _23560_ (.A(_20413_),
    .B(\inst$top.soc.cpu.sink__payload$24[88] ),
    .Y(_20614_));
 sky130_fd_sc_hd__nand2_1 _23561_ (.A(net2823),
    .B(\inst$top.soc.cpu.sink__payload$24[104] ),
    .Y(_20615_));
 sky130_fd_sc_hd__nand2_1 _23562_ (.A(_20614_),
    .B(_20615_),
    .Y(_20616_));
 sky130_fd_sc_hd__nand2_1 _23563_ (.A(_20412_),
    .B(_20616_),
    .Y(_20617_));
 sky130_fd_sc_hd__o311ai_0 _23564_ (.A1(_20611_),
    .A2(_20612_),
    .A3(_20419_),
    .B1(_20613_),
    .C1(_20617_),
    .Y(_20618_));
 sky130_fd_sc_hd__nor2_1 _23565_ (.A(net2827),
    .B(\inst$top.soc.cpu.sink__payload$24[47] ),
    .Y(_20619_));
 sky130_fd_sc_hd__nor2_1 _23566_ (.A(\inst$top.soc.cpu.multiplier.w_result[6] ),
    .B(net2200),
    .Y(_20620_));
 sky130_fd_sc_hd__nor2_1 _23567_ (.A(_20619_),
    .B(_20620_),
    .Y(_20621_));
 sky130_fd_sc_hd__mux2i_1 _23568_ (.A0(_20618_),
    .A1(_20621_),
    .S(net2207),
    .Y(_20622_));
 sky130_fd_sc_hd__inv_2 _23569_ (.A(_20622_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[6] ));
 sky130_fd_sc_hd__inv_1 _23570_ (.A(\inst$top.soc.cpu.sink__payload$12[7] ),
    .Y(_20623_));
 sky130_fd_sc_hd__nand2_1 _23571_ (.A(net2549),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[7] ),
    .Y(_20624_));
 sky130_fd_sc_hd__nand2_1 _23572_ (.A(net2886),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[7] ),
    .Y(_20625_));
 sky130_fd_sc_hd__nand2_1 _23573_ (.A(_20624_),
    .B(_20625_),
    .Y(_20626_));
 sky130_fd_sc_hd__nand2_1 _23574_ (.A(net1828),
    .B(_20626_),
    .Y(_20627_));
 sky130_fd_sc_hd__o21ai_1 _23575_ (.A1(_20623_),
    .A2(net1832),
    .B1(_20627_),
    .Y(_20628_));
 sky130_fd_sc_hd__xor2_1 _23577_ (.A(net1977),
    .B(net1345),
    .X(_03136_));
 sky130_fd_sc_hd__inv_2 _23578_ (.A(_03136_),
    .Y(_03140_));
 sky130_fd_sc_hd__clkinv_1 _23579_ (.A(net1398),
    .Y(_20630_));
 sky130_fd_sc_hd__inv_1 _23581_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mtip.x_data ),
    .Y(_20631_));
 sky130_fd_sc_hd__inv_1 _23584_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[7] ),
    .Y(_20634_));
 sky130_fd_sc_hd__inv_1 _23585_ (.A(\inst$top.soc.cpu.exception.csr_bank.mstatus_x_select ),
    .Y(_20635_));
 sky130_fd_sc_hd__inv_1 _23586_ (.A(\inst$top.soc.cpu.exception.csr_bank.mstatus.mpie.x_data ),
    .Y(_20636_));
 sky130_fd_sc_hd__o22ai_1 _23587_ (.A1(net2211),
    .A2(_20634_),
    .B1(_20635_),
    .B2(_20636_),
    .Y(_20637_));
 sky130_fd_sc_hd__a221oi_1 _23588_ (.A1(net2892),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[5] ),
    .B1(\inst$top.soc.cpu.exception.csr_bank.mie_x_select ),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mie.mtie.x_data ),
    .C1(_20637_),
    .Y(_20638_));
 sky130_fd_sc_hd__nand2_1 _23589_ (.A(net2897),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[7] ),
    .Y(_20639_));
 sky130_fd_sc_hd__nand2_1 _23590_ (.A(net2912),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[7] ),
    .Y(_20640_));
 sky130_fd_sc_hd__nand2_1 _23591_ (.A(net2908),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[5] ),
    .Y(_20641_));
 sky130_fd_sc_hd__nand4_1 _23592_ (.A(_20638_),
    .B(_20639_),
    .C(_20640_),
    .D(_20641_),
    .Y(_20642_));
 sky130_fd_sc_hd__a21oi_1 _23593_ (.A1(net2893),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[7] ),
    .B1(_20642_),
    .Y(_20643_));
 sky130_fd_sc_hd__o21ai_0 _23594_ (.A1(_20509_),
    .A2(_20631_),
    .B1(_20643_),
    .Y(_20644_));
 sky130_fd_sc_hd__nand2_1 _23596_ (.A(_20644_),
    .B(net1981),
    .Y(_20646_));
 sky130_fd_sc_hd__o21ai_1 _23597_ (.A1(net2845),
    .A2(net3043),
    .B1(_20646_),
    .Y(_03135_));
 sky130_fd_sc_hd__inv_2 _23598_ (.A(_03135_),
    .Y(_03139_));
 sky130_fd_sc_hd__nor2_1 _23600_ (.A(\inst$top.soc.cpu.multiplier.w_result[7] ),
    .B(net2196),
    .Y(_20648_));
 sky130_fd_sc_hd__o21ai_0 _23602_ (.A1(net2825),
    .A2(\inst$top.soc.cpu.sink__payload$24[48] ),
    .B1(net2201),
    .Y(_20650_));
 sky130_fd_sc_hd__inv_1 _23603_ (.A(\inst$top.soc.cpu.sink__payload$24[81] ),
    .Y(_20651_));
 sky130_fd_sc_hd__nor2_1 _23604_ (.A(\inst$top.soc.cpu.sink__payload$24[39] ),
    .B(_20417_),
    .Y(_20652_));
 sky130_fd_sc_hd__inv_1 _23605_ (.A(_20652_),
    .Y(_20653_));
 sky130_fd_sc_hd__nand2_1 _23606_ (.A(_20413_),
    .B(_20651_),
    .Y(_20654_));
 sky130_fd_sc_hd__o21ai_0 _23607_ (.A1(\inst$top.soc.cpu.sink__payload$24[97] ),
    .A2(_20413_),
    .B1(_20654_),
    .Y(_20655_));
 sky130_fd_sc_hd__inv_1 _23608_ (.A(\inst$top.soc.cpu.sink__payload$24[89] ),
    .Y(_20656_));
 sky130_fd_sc_hd__nand2_1 _23609_ (.A(net2822),
    .B(\inst$top.soc.cpu.sink__payload$24[105] ),
    .Y(_20657_));
 sky130_fd_sc_hd__o21ai_0 _23610_ (.A1(net2822),
    .A2(_20656_),
    .B1(_20657_),
    .Y(_20658_));
 sky130_fd_sc_hd__nand2_1 _23611_ (.A(_20655_),
    .B(_20409_),
    .Y(_20659_));
 sky130_fd_sc_hd__o211ai_1 _23612_ (.A1(_20409_),
    .A2(_20658_),
    .B1(_20410_),
    .C1(_20659_),
    .Y(_20660_));
 sky130_fd_sc_hd__o221ai_1 _23613_ (.A1(_20651_),
    .A2(_20447_),
    .B1(_20653_),
    .B2(_20655_),
    .C1(_20660_),
    .Y(_20661_));
 sky130_fd_sc_hd__nand2_1 _23614_ (.A(_20661_),
    .B(\inst$top.soc.cpu.d.sink__payload$16.load ),
    .Y(_20662_));
 sky130_fd_sc_hd__o21a_1 _23615_ (.A1(_20648_),
    .A2(_20650_),
    .B1(_20662_),
    .X(_20663_));
 sky130_fd_sc_hd__inv_2 _23616_ (.A(_20663_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[7] ));
 sky130_fd_sc_hd__inv_1 _23617_ (.A(\inst$top.soc.cpu.sink__payload$12[8] ),
    .Y(_20664_));
 sky130_fd_sc_hd__nand2_1 _23619_ (.A(net2549),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[8] ),
    .Y(_20666_));
 sky130_fd_sc_hd__nand2_1 _23620_ (.A(net2888),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[8] ),
    .Y(_20667_));
 sky130_fd_sc_hd__nand2_1 _23621_ (.A(_20666_),
    .B(_20667_),
    .Y(_20668_));
 sky130_fd_sc_hd__nand2_1 _23622_ (.A(net1829),
    .B(_20668_),
    .Y(_20669_));
 sky130_fd_sc_hd__o21ai_1 _23623_ (.A1(_20664_),
    .A2(net1832),
    .B1(_20669_),
    .Y(_20670_));
 sky130_fd_sc_hd__xor2_1 _23625_ (.A(net1979),
    .B(net1341),
    .X(_03143_));
 sky130_fd_sc_hd__inv_2 _23626_ (.A(_03143_),
    .Y(_03147_));
 sky130_fd_sc_hd__inv_1 _23628_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[6] ),
    .Y(_20672_));
 sky130_fd_sc_hd__nand2_1 _23629_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa_x_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[8] ),
    .Y(_20673_));
 sky130_fd_sc_hd__o21ai_0 _23630_ (.A1(net2208),
    .A2(_20672_),
    .B1(_20673_),
    .Y(_20674_));
 sky130_fd_sc_hd__a221oi_1 _23631_ (.A1(net2898),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[8] ),
    .B1(net2910),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[6] ),
    .C1(_20674_),
    .Y(_20675_));
 sky130_fd_sc_hd__nand2_1 _23632_ (.A(net2895),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[8] ),
    .Y(_20676_));
 sky130_fd_sc_hd__nand2_1 _23633_ (.A(net2914),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[8] ),
    .Y(_20677_));
 sky130_fd_sc_hd__nand3_1 _23634_ (.A(_20675_),
    .B(_20676_),
    .C(_20677_),
    .Y(_20678_));
 sky130_fd_sc_hd__nand2_1 _23635_ (.A(_20678_),
    .B(net1981),
    .Y(_20679_));
 sky130_fd_sc_hd__o21ai_1 _23636_ (.A1(net2847),
    .A2(net1399),
    .B1(_20679_),
    .Y(_03142_));
 sky130_fd_sc_hd__inv_2 _23637_ (.A(_03142_),
    .Y(_03146_));
 sky130_fd_sc_hd__nor2_1 _23638_ (.A(\inst$top.soc.cpu.multiplier.w_result[8] ),
    .B(net2198),
    .Y(_20680_));
 sky130_fd_sc_hd__o21ai_0 _23640_ (.A1(net2827),
    .A2(\inst$top.soc.cpu.sink__payload$24[49] ),
    .B1(net2206),
    .Y(_20682_));
 sky130_fd_sc_hd__nor2_1 _23641_ (.A(\inst$top.soc.cpu.sink__payload$24[40] ),
    .B(_20660_),
    .Y(_20683_));
 sky130_fd_sc_hd__a221oi_1 _23642_ (.A1(\inst$top.soc.cpu.sink__payload$24[82] ),
    .A2(net1983),
    .B1(_20408_),
    .B2(_20652_),
    .C1(net1160),
    .Y(_20684_));
 sky130_fd_sc_hd__o22ai_1 _23643_ (.A1(_20680_),
    .A2(_20682_),
    .B1(net2206),
    .B2(_20684_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[8] ));
 sky130_fd_sc_hd__inv_1 _23644_ (.A(\inst$top.soc.cpu.sink__payload$12[9] ),
    .Y(_20685_));
 sky130_fd_sc_hd__nand2_1 _23645_ (.A(net2549),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[9] ),
    .Y(_20686_));
 sky130_fd_sc_hd__nand2_1 _23646_ (.A(net2888),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[9] ),
    .Y(_20687_));
 sky130_fd_sc_hd__nand2_1 _23647_ (.A(_20686_),
    .B(_20687_),
    .Y(_20688_));
 sky130_fd_sc_hd__nand2_1 _23648_ (.A(net1829),
    .B(_20688_),
    .Y(_20689_));
 sky130_fd_sc_hd__o21ai_1 _23649_ (.A1(_20685_),
    .A2(net1832),
    .B1(_20689_),
    .Y(_20690_));
 sky130_fd_sc_hd__xor2_1 _23651_ (.A(net1978),
    .B(net1336),
    .X(_03150_));
 sky130_fd_sc_hd__inv_2 _23652_ (.A(_03150_),
    .Y(_03154_));
 sky130_fd_sc_hd__inv_1 _23653_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[9] ),
    .Y(_20692_));
 sky130_fd_sc_hd__nand2_1 _23654_ (.A(net2898),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[9] ),
    .Y(_20693_));
 sky130_fd_sc_hd__nand2_1 _23655_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec_x_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[7] ),
    .Y(_20694_));
 sky130_fd_sc_hd__nand2_1 _23656_ (.A(net2910),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[7] ),
    .Y(_20695_));
 sky130_fd_sc_hd__o2111ai_1 _23657_ (.A1(net2212),
    .A2(_20692_),
    .B1(_20693_),
    .C1(_20694_),
    .D1(_20695_),
    .Y(_20696_));
 sky130_fd_sc_hd__a221oi_1 _23658_ (.A1(net2914),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[9] ),
    .B1(net2895),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[9] ),
    .C1(_20696_),
    .Y(_20697_));
 sky130_fd_sc_hd__nor2_1 _23659_ (.A(_20480_),
    .B(_20697_),
    .Y(_20698_));
 sky130_fd_sc_hd__inv_1 _23660_ (.A(_20698_),
    .Y(_20699_));
 sky130_fd_sc_hd__o21ai_1 _23661_ (.A1(net2846),
    .A2(_20067_),
    .B1(_20699_),
    .Y(_03149_));
 sky130_fd_sc_hd__inv_2 _23662_ (.A(_03149_),
    .Y(_03153_));
 sky130_fd_sc_hd__nor2_1 _23663_ (.A(\inst$top.soc.cpu.multiplier.w_result[9] ),
    .B(net2198),
    .Y(_20700_));
 sky130_fd_sc_hd__o21ai_0 _23665_ (.A1(net2827),
    .A2(\inst$top.soc.cpu.sink__payload$24[50] ),
    .B1(net2206),
    .Y(_20702_));
 sky130_fd_sc_hd__a221oi_1 _23667_ (.A1(\inst$top.soc.cpu.sink__payload$24[83] ),
    .A2(net1982),
    .B1(_20652_),
    .B2(_20444_),
    .C1(net1161),
    .Y(_20704_));
 sky130_fd_sc_hd__o22ai_1 _23668_ (.A1(_20700_),
    .A2(_20702_),
    .B1(net2206),
    .B2(_20704_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[9] ));
 sky130_fd_sc_hd__clkinv_1 _23669_ (.A(\inst$top.soc.cpu.sink__payload$12[10] ),
    .Y(_20705_));
 sky130_fd_sc_hd__nand2_1 _23670_ (.A(net2547),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[10] ),
    .Y(_20706_));
 sky130_fd_sc_hd__nand2_1 _23671_ (.A(net2887),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[10] ),
    .Y(_20707_));
 sky130_fd_sc_hd__nand2_1 _23672_ (.A(_20706_),
    .B(_20707_),
    .Y(_20708_));
 sky130_fd_sc_hd__nand2_1 _23673_ (.A(_19881_),
    .B(_20708_),
    .Y(_20709_));
 sky130_fd_sc_hd__o21ai_0 _23674_ (.A1(_20705_),
    .A2(net1832),
    .B1(_20709_),
    .Y(_20710_));
 sky130_fd_sc_hd__xor2_1 _23676_ (.A(net1979),
    .B(net1331),
    .X(_03157_));
 sky130_fd_sc_hd__inv_2 _23677_ (.A(_03157_),
    .Y(_03161_));
 sky130_fd_sc_hd__inv_1 _23679_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[10] ),
    .Y(_20713_));
 sky130_fd_sc_hd__inv_1 _23680_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[8] ),
    .Y(_20714_));
 sky130_fd_sc_hd__o22ai_1 _23681_ (.A1(net2212),
    .A2(_20713_),
    .B1(net2208),
    .B2(_20714_),
    .Y(_20715_));
 sky130_fd_sc_hd__a21oi_1 _23682_ (.A1(net2898),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[10] ),
    .B1(_20715_),
    .Y(_20716_));
 sky130_fd_sc_hd__nand2_1 _23683_ (.A(net2910),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[8] ),
    .Y(_20717_));
 sky130_fd_sc_hd__nand2_1 _23684_ (.A(_20716_),
    .B(_20717_),
    .Y(_20718_));
 sky130_fd_sc_hd__a221oi_1 _23685_ (.A1(net2914),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[10] ),
    .B1(net2895),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[10] ),
    .C1(_20718_),
    .Y(_20719_));
 sky130_fd_sc_hd__nor2_1 _23686_ (.A(_20480_),
    .B(_20719_),
    .Y(_20720_));
 sky130_fd_sc_hd__inv_1 _23687_ (.A(_20720_),
    .Y(_20721_));
 sky130_fd_sc_hd__o21ai_1 _23688_ (.A1(net2847),
    .A2(_20061_),
    .B1(_20721_),
    .Y(_03156_));
 sky130_fd_sc_hd__inv_2 _23689_ (.A(_03156_),
    .Y(_03160_));
 sky130_fd_sc_hd__nor2_1 _23690_ (.A(\inst$top.soc.cpu.multiplier.w_result[10] ),
    .B(net2196),
    .Y(_20722_));
 sky130_fd_sc_hd__o21ai_0 _23691_ (.A1(net2825),
    .A2(\inst$top.soc.cpu.sink__payload$24[51] ),
    .B1(net2203),
    .Y(_20723_));
 sky130_fd_sc_hd__a221oi_1 _23693_ (.A1(\inst$top.soc.cpu.sink__payload$24[84] ),
    .A2(net1982),
    .B1(_20652_),
    .B2(_20490_),
    .C1(net1161),
    .Y(_20725_));
 sky130_fd_sc_hd__o22ai_1 _23694_ (.A1(_20722_),
    .A2(_20723_),
    .B1(net2203),
    .B2(_20725_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[10] ));
 sky130_fd_sc_hd__clkinv_1 _23695_ (.A(\inst$top.soc.cpu.sink__payload$12[11] ),
    .Y(_20726_));
 sky130_fd_sc_hd__nand2_1 _23696_ (.A(net2550),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[11] ),
    .Y(_20727_));
 sky130_fd_sc_hd__nand2_1 _23697_ (.A(net2887),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[11] ),
    .Y(_20728_));
 sky130_fd_sc_hd__nand2_1 _23698_ (.A(_20727_),
    .B(_20728_),
    .Y(_20729_));
 sky130_fd_sc_hd__nand2_1 _23699_ (.A(net1828),
    .B(_20729_),
    .Y(_20730_));
 sky130_fd_sc_hd__o21ai_0 _23700_ (.A1(_20726_),
    .A2(net1831),
    .B1(_20730_),
    .Y(_20731_));
 sky130_fd_sc_hd__xor2_1 _23702_ (.A(net1979),
    .B(net1327),
    .X(_03164_));
 sky130_fd_sc_hd__inv_2 _23703_ (.A(_03164_),
    .Y(_03168_));
 sky130_fd_sc_hd__nand2_1 _23704_ (.A(_19976_),
    .B(_20050_),
    .Y(_20733_));
 sky130_fd_sc_hd__o21ai_4 _23705_ (.A1(net1827),
    .A2(_20053_),
    .B1(_20733_),
    .Y(_20734_));
 sky130_fd_sc_hd__inv_1 _23707_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.meip.x_data ),
    .Y(_20735_));
 sky130_fd_sc_hd__nand2_1 _23708_ (.A(net2896),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[11] ),
    .Y(_20736_));
 sky130_fd_sc_hd__inv_1 _23709_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[9] ),
    .Y(_20737_));
 sky130_fd_sc_hd__nand2_1 _23710_ (.A(net2908),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[9] ),
    .Y(_20738_));
 sky130_fd_sc_hd__nand2_1 _23711_ (.A(net2897),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[11] ),
    .Y(_20739_));
 sky130_fd_sc_hd__inv_1 _23712_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[11] ),
    .Y(_20740_));
 sky130_fd_sc_hd__nand2_1 _23713_ (.A(\inst$top.soc.cpu.exception.csr_bank.mstatus_x_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.mstatus.mpp.x_data[0] ),
    .Y(_20741_));
 sky130_fd_sc_hd__o21ai_0 _23714_ (.A1(net2211),
    .A2(_20740_),
    .B1(_20741_),
    .Y(_20742_));
 sky130_fd_sc_hd__a21oi_1 _23715_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mie_x_select ),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mie.meie.x_data ),
    .B1(_20742_),
    .Y(_20743_));
 sky130_fd_sc_hd__o2111ai_1 _23716_ (.A1(net2210),
    .A2(_20737_),
    .B1(_20738_),
    .C1(_20739_),
    .D1(_20743_),
    .Y(_20744_));
 sky130_fd_sc_hd__a21oi_1 _23717_ (.A1(net2912),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[11] ),
    .B1(_20744_),
    .Y(_20745_));
 sky130_fd_sc_hd__o211ai_1 _23718_ (.A1(_20509_),
    .A2(_20735_),
    .B1(_20736_),
    .C1(_20745_),
    .Y(_20746_));
 sky130_fd_sc_hd__nand2_1 _23719_ (.A(_20746_),
    .B(net1981),
    .Y(_20747_));
 sky130_fd_sc_hd__o21ai_1 _23720_ (.A1(net2847),
    .A2(_20734_),
    .B1(_20747_),
    .Y(_03163_));
 sky130_fd_sc_hd__inv_2 _23721_ (.A(_03163_),
    .Y(_03167_));
 sky130_fd_sc_hd__nor2_1 _23722_ (.A(\inst$top.soc.cpu.multiplier.w_result[11] ),
    .B(net2196),
    .Y(_20748_));
 sky130_fd_sc_hd__o21ai_0 _23723_ (.A1(net2825),
    .A2(\inst$top.soc.cpu.sink__payload$24[52] ),
    .B1(net2203),
    .Y(_20749_));
 sky130_fd_sc_hd__a221oi_1 _23724_ (.A1(\inst$top.soc.cpu.sink__payload$24[85] ),
    .A2(net1982),
    .B1(_20652_),
    .B2(_20529_),
    .C1(net1161),
    .Y(_20750_));
 sky130_fd_sc_hd__o22ai_1 _23725_ (.A1(_20748_),
    .A2(_20749_),
    .B1(net2203),
    .B2(_20750_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[11] ));
 sky130_fd_sc_hd__inv_1 _23726_ (.A(\inst$top.soc.cpu.sink__payload$12[12] ),
    .Y(_20751_));
 sky130_fd_sc_hd__nand2_1 _23727_ (.A(net2548),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[12] ),
    .Y(_20752_));
 sky130_fd_sc_hd__nand2_1 _23728_ (.A(net2888),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[12] ),
    .Y(_20753_));
 sky130_fd_sc_hd__nand2_1 _23729_ (.A(_20752_),
    .B(_20753_),
    .Y(_20754_));
 sky130_fd_sc_hd__nand2_1 _23730_ (.A(net1829),
    .B(_20754_),
    .Y(_20755_));
 sky130_fd_sc_hd__o21ai_1 _23731_ (.A1(_20751_),
    .A2(net1831),
    .B1(_20755_),
    .Y(_20756_));
 sky130_fd_sc_hd__xor2_1 _23733_ (.A(net1978),
    .B(net1322),
    .X(_03171_));
 sky130_fd_sc_hd__inv_2 _23734_ (.A(_03171_),
    .Y(_03175_));
 sky130_fd_sc_hd__nand2_1 _23735_ (.A(net1827),
    .B(_20043_),
    .Y(_20758_));
 sky130_fd_sc_hd__o21ai_4 _23736_ (.A1(net1827),
    .A2(_20046_),
    .B1(_20758_),
    .Y(_20759_));
 sky130_fd_sc_hd__inv_1 _23738_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[10] ),
    .Y(_20760_));
 sky130_fd_sc_hd__nand2_1 _23739_ (.A(net2895),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[12] ),
    .Y(_20761_));
 sky130_fd_sc_hd__nand2_1 _23740_ (.A(\inst$top.soc.cpu.exception.csr_bank.mstatus_x_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.mstatus.mpp.x_data[1] ),
    .Y(_20762_));
 sky130_fd_sc_hd__a22o_1 _23741_ (.A1(\inst$top.soc.cpu.exception.csr_bank.misa_x_select ),
    .A2(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[12] ),
    .B1(net2914),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[12] ),
    .X(_20763_));
 sky130_fd_sc_hd__a221oi_1 _23742_ (.A1(net2898),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[12] ),
    .B1(net2910),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[10] ),
    .C1(_20763_),
    .Y(_20764_));
 sky130_fd_sc_hd__o2111ai_1 _23743_ (.A1(net2209),
    .A2(_20760_),
    .B1(_20761_),
    .C1(_20762_),
    .D1(_20764_),
    .Y(_20765_));
 sky130_fd_sc_hd__nand2_1 _23744_ (.A(_20765_),
    .B(net1980),
    .Y(_20766_));
 sky130_fd_sc_hd__o21ai_1 _23745_ (.A1(net2846),
    .A2(_20759_),
    .B1(_20766_),
    .Y(_03170_));
 sky130_fd_sc_hd__inv_2 _23746_ (.A(_03170_),
    .Y(_03174_));
 sky130_fd_sc_hd__nor2_1 _23747_ (.A(\inst$top.soc.cpu.multiplier.w_result[12] ),
    .B(net2198),
    .Y(_20767_));
 sky130_fd_sc_hd__o21ai_0 _23748_ (.A1(net2827),
    .A2(\inst$top.soc.cpu.sink__payload$24[53] ),
    .B1(net2206),
    .Y(_20768_));
 sky130_fd_sc_hd__a221oi_1 _23749_ (.A1(\inst$top.soc.cpu.sink__payload$24[86] ),
    .A2(net1982),
    .B1(_20652_),
    .B2(_20558_),
    .C1(net1161),
    .Y(_20769_));
 sky130_fd_sc_hd__o22ai_2 _23750_ (.A1(_20767_),
    .A2(_20768_),
    .B1(net2206),
    .B2(_20769_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[12] ));
 sky130_fd_sc_hd__inv_1 _23752_ (.A(\inst$top.soc.cpu.sink__payload$12[13] ),
    .Y(_20771_));
 sky130_fd_sc_hd__nand2_1 _23753_ (.A(net2547),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[13] ),
    .Y(_20772_));
 sky130_fd_sc_hd__nand2_1 _23754_ (.A(net2889),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[13] ),
    .Y(_20773_));
 sky130_fd_sc_hd__nand2_1 _23755_ (.A(_20772_),
    .B(_20773_),
    .Y(_20774_));
 sky130_fd_sc_hd__nand2_1 _23756_ (.A(net1830),
    .B(_20774_),
    .Y(_20775_));
 sky130_fd_sc_hd__o21ai_0 _23757_ (.A1(_20771_),
    .A2(net1832),
    .B1(_20775_),
    .Y(_20776_));
 sky130_fd_sc_hd__xor2_1 _23759_ (.A(net1978),
    .B(net1317),
    .X(_03178_));
 sky130_fd_sc_hd__inv_2 _23760_ (.A(_03178_),
    .Y(_03182_));
 sky130_fd_sc_hd__inv_1 _23761_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[11] ),
    .Y(_20778_));
 sky130_fd_sc_hd__nand2_1 _23762_ (.A(net2913),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[13] ),
    .Y(_20779_));
 sky130_fd_sc_hd__nand2_1 _23763_ (.A(net2910),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[11] ),
    .Y(_20780_));
 sky130_fd_sc_hd__nand2_1 _23764_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa_x_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[13] ),
    .Y(_20781_));
 sky130_fd_sc_hd__o2111ai_1 _23765_ (.A1(net2208),
    .A2(_20778_),
    .B1(_20779_),
    .C1(_20780_),
    .D1(_20781_),
    .Y(_20782_));
 sky130_fd_sc_hd__a221oi_1 _23766_ (.A1(net2898),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[13] ),
    .B1(net2894),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[13] ),
    .C1(_20782_),
    .Y(_20783_));
 sky130_fd_sc_hd__nor2_1 _23767_ (.A(_20480_),
    .B(_20783_),
    .Y(_20784_));
 sky130_fd_sc_hd__inv_1 _23768_ (.A(_20784_),
    .Y(_20785_));
 sky130_fd_sc_hd__o21ai_1 _23769_ (.A1(net2843),
    .A2(_03017_),
    .B1(_20785_),
    .Y(_03177_));
 sky130_fd_sc_hd__inv_2 _23770_ (.A(_03177_),
    .Y(_03181_));
 sky130_fd_sc_hd__nor2_1 _23771_ (.A(\inst$top.soc.cpu.multiplier.w_result[13] ),
    .B(net2196),
    .Y(_20786_));
 sky130_fd_sc_hd__o21ai_0 _23772_ (.A1(net2826),
    .A2(\inst$top.soc.cpu.sink__payload$24[54] ),
    .B1(net2204),
    .Y(_20787_));
 sky130_fd_sc_hd__a221oi_1 _23773_ (.A1(\inst$top.soc.cpu.sink__payload$24[87] ),
    .A2(net1983),
    .B1(_20652_),
    .B2(_20587_),
    .C1(net1160),
    .Y(_20788_));
 sky130_fd_sc_hd__o22ai_2 _23774_ (.A1(_20786_),
    .A2(_20787_),
    .B1(net2204),
    .B2(_20788_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[13] ));
 sky130_fd_sc_hd__clkinv_1 _23775_ (.A(\inst$top.soc.cpu.sink__payload$12[14] ),
    .Y(_20789_));
 sky130_fd_sc_hd__nand2_1 _23776_ (.A(net2546),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[14] ),
    .Y(_20790_));
 sky130_fd_sc_hd__nand2_1 _23777_ (.A(net2888),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[14] ),
    .Y(_20791_));
 sky130_fd_sc_hd__nand2_1 _23778_ (.A(_20790_),
    .B(_20791_),
    .Y(_20792_));
 sky130_fd_sc_hd__nand2_1 _23779_ (.A(net1830),
    .B(_20792_),
    .Y(_20793_));
 sky130_fd_sc_hd__o21ai_0 _23780_ (.A1(_20789_),
    .A2(net1832),
    .B1(_20793_),
    .Y(_20794_));
 sky130_fd_sc_hd__xor2_1 _23782_ (.A(net1977),
    .B(net1312),
    .X(_03185_));
 sky130_fd_sc_hd__inv_2 _23783_ (.A(_03185_),
    .Y(_03189_));
 sky130_fd_sc_hd__inv_1 _23784_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[12] ),
    .Y(_20796_));
 sky130_fd_sc_hd__nand2_1 _23785_ (.A(net2914),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[14] ),
    .Y(_20797_));
 sky130_fd_sc_hd__nand2_1 _23786_ (.A(net2910),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[12] ),
    .Y(_20798_));
 sky130_fd_sc_hd__nand2_1 _23787_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa_x_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[14] ),
    .Y(_20799_));
 sky130_fd_sc_hd__o2111ai_1 _23788_ (.A1(net2208),
    .A2(_20796_),
    .B1(_20797_),
    .C1(_20798_),
    .D1(_20799_),
    .Y(_20800_));
 sky130_fd_sc_hd__a221oi_1 _23789_ (.A1(net2898),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[14] ),
    .B1(net2895),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[14] ),
    .C1(_20800_),
    .Y(_20801_));
 sky130_fd_sc_hd__nor2_1 _23790_ (.A(_20480_),
    .B(_20801_),
    .Y(_20802_));
 sky130_fd_sc_hd__inv_1 _23791_ (.A(_20802_),
    .Y(_20803_));
 sky130_fd_sc_hd__o21ai_1 _23792_ (.A1(net2845),
    .A2(_03011_),
    .B1(_20803_),
    .Y(_03184_));
 sky130_fd_sc_hd__inv_2 _23793_ (.A(_03184_),
    .Y(_03188_));
 sky130_fd_sc_hd__nor2_1 _23794_ (.A(\inst$top.soc.cpu.multiplier.w_result[14] ),
    .B(net2200),
    .Y(_20804_));
 sky130_fd_sc_hd__o21ai_0 _23795_ (.A1(net2827),
    .A2(\inst$top.soc.cpu.sink__payload$24[55] ),
    .B1(net2207),
    .Y(_20805_));
 sky130_fd_sc_hd__a221oi_1 _23796_ (.A1(\inst$top.soc.cpu.sink__payload$24[88] ),
    .A2(net1983),
    .B1(_20652_),
    .B2(_20616_),
    .C1(net1160),
    .Y(_20806_));
 sky130_fd_sc_hd__o22ai_2 _23797_ (.A1(_20804_),
    .A2(_20805_),
    .B1(net2202),
    .B2(_20806_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[14] ));
 sky130_fd_sc_hd__inv_1 _23798_ (.A(\inst$top.soc.cpu.sink__payload$12[15] ),
    .Y(_20807_));
 sky130_fd_sc_hd__nand2_1 _23799_ (.A(net2546),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[15] ),
    .Y(_20808_));
 sky130_fd_sc_hd__nand2_1 _23800_ (.A(net2886),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[15] ),
    .Y(_20809_));
 sky130_fd_sc_hd__nand2_1 _23801_ (.A(_20808_),
    .B(_20809_),
    .Y(_20810_));
 sky130_fd_sc_hd__nand2_1 _23802_ (.A(net1828),
    .B(_20810_),
    .Y(_20811_));
 sky130_fd_sc_hd__o21ai_1 _23803_ (.A1(_20807_),
    .A2(net1832),
    .B1(_20811_),
    .Y(_20812_));
 sky130_fd_sc_hd__xor2_1 _23805_ (.A(net1978),
    .B(net1308),
    .X(_03192_));
 sky130_fd_sc_hd__inv_2 _23806_ (.A(_03192_),
    .Y(_03196_));
 sky130_fd_sc_hd__inv_1 _23810_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[15] ),
    .Y(_20816_));
 sky130_fd_sc_hd__inv_1 _23811_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[13] ),
    .Y(_20817_));
 sky130_fd_sc_hd__o22ai_1 _23812_ (.A1(net2212),
    .A2(_20816_),
    .B1(net2208),
    .B2(_20817_),
    .Y(_20818_));
 sky130_fd_sc_hd__a221oi_1 _23813_ (.A1(net2898),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[15] ),
    .B1(net2910),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[13] ),
    .C1(_20818_),
    .Y(_20819_));
 sky130_fd_sc_hd__nand2_1 _23814_ (.A(net2895),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[15] ),
    .Y(_20820_));
 sky130_fd_sc_hd__nand2_1 _23816_ (.A(net2914),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[15] ),
    .Y(_20822_));
 sky130_fd_sc_hd__nand3_1 _23817_ (.A(_20819_),
    .B(_20820_),
    .C(_20822_),
    .Y(_20823_));
 sky130_fd_sc_hd__nand2_1 _23818_ (.A(_20823_),
    .B(_20481_),
    .Y(_20824_));
 sky130_fd_sc_hd__o21ai_1 _23819_ (.A1(net2846),
    .A2(net1713),
    .B1(_20824_),
    .Y(_03191_));
 sky130_fd_sc_hd__inv_2 _23820_ (.A(_03191_),
    .Y(_03195_));
 sky130_fd_sc_hd__nor2_1 _23821_ (.A(\inst$top.soc.cpu.multiplier.w_result[15] ),
    .B(net2196),
    .Y(_05592_));
 sky130_fd_sc_hd__o21ai_0 _23822_ (.A1(net2825),
    .A2(\inst$top.soc.cpu.sink__payload$24[56] ),
    .B1(net2203),
    .Y(_05593_));
 sky130_fd_sc_hd__nand2_1 _23823_ (.A(_20658_),
    .B(_20652_),
    .Y(_05594_));
 sky130_fd_sc_hd__o21ai_0 _23824_ (.A1(_20656_),
    .A2(_20447_),
    .B1(_05594_),
    .Y(_05595_));
 sky130_fd_sc_hd__o21ai_0 _23825_ (.A1(_05595_),
    .A2(net1161),
    .B1(\inst$top.soc.cpu.d.sink__payload$16.load ),
    .Y(_05596_));
 sky130_fd_sc_hd__o21a_1 _23826_ (.A1(_05592_),
    .A2(_05593_),
    .B1(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__inv_2 _23827_ (.A(_05597_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[15] ));
 sky130_fd_sc_hd__inv_1 _23828_ (.A(\inst$top.soc.cpu.sink__payload$12[16] ),
    .Y(_05598_));
 sky130_fd_sc_hd__nand2_1 _23829_ (.A(net2547),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[16] ),
    .Y(_05599_));
 sky130_fd_sc_hd__nand2_1 _23830_ (.A(net2887),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[16] ),
    .Y(_05600_));
 sky130_fd_sc_hd__nand2_1 _23831_ (.A(_05599_),
    .B(_05600_),
    .Y(_05601_));
 sky130_fd_sc_hd__nand2_1 _23832_ (.A(net1830),
    .B(_05601_),
    .Y(_05602_));
 sky130_fd_sc_hd__o21ai_0 _23833_ (.A1(_05598_),
    .A2(net1831),
    .B1(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__xor2_1 _23835_ (.A(_20498_),
    .B(net1303),
    .X(_03199_));
 sky130_fd_sc_hd__inv_2 _23836_ (.A(_03199_),
    .Y(_03203_));
 sky130_fd_sc_hd__inv_1 _23838_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[14] ),
    .Y(_05605_));
 sky130_fd_sc_hd__nand2_1 _23839_ (.A(net2894),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[16] ),
    .Y(_05606_));
 sky130_fd_sc_hd__o21ai_0 _23840_ (.A1(net2208),
    .A2(_05605_),
    .B1(_05606_),
    .Y(_05607_));
 sky130_fd_sc_hd__inv_1 _23841_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[0] ),
    .Y(_05608_));
 sky130_fd_sc_hd__nand2_1 _23842_ (.A(net2912),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[16] ),
    .Y(_05609_));
 sky130_fd_sc_hd__nand2_1 _23843_ (.A(net2911),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[14] ),
    .Y(_05610_));
 sky130_fd_sc_hd__inv_1 _23844_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[16] ),
    .Y(_05611_));
 sky130_fd_sc_hd__nand2_1 _23845_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie_x_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[0] ),
    .Y(_05612_));
 sky130_fd_sc_hd__o21ai_0 _23846_ (.A1(net2213),
    .A2(_05611_),
    .B1(_05612_),
    .Y(_05613_));
 sky130_fd_sc_hd__a21oi_1 _23847_ (.A1(net2897),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[16] ),
    .B1(_05613_),
    .Y(_05614_));
 sky130_fd_sc_hd__o2111ai_1 _23848_ (.A1(_20509_),
    .A2(_05608_),
    .B1(_05609_),
    .C1(_05610_),
    .D1(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__o21ai_0 _23849_ (.A1(_05607_),
    .A2(_05615_),
    .B1(net1980),
    .Y(_05616_));
 sky130_fd_sc_hd__o21ai_1 _23850_ (.A1(net2848),
    .A2(net1716),
    .B1(net3045),
    .Y(_03198_));
 sky130_fd_sc_hd__inv_2 _23851_ (.A(_03198_),
    .Y(_03202_));
 sky130_fd_sc_hd__nor2_1 _23852_ (.A(\inst$top.soc.cpu.multiplier.w_result[16] ),
    .B(net2198),
    .Y(_05617_));
 sky130_fd_sc_hd__o21ai_0 _23853_ (.A1(net2826),
    .A2(\inst$top.soc.cpu.sink__payload$24[57] ),
    .B1(net2204),
    .Y(_05618_));
 sky130_fd_sc_hd__nor2_1 _23854_ (.A(\inst$top.soc.cpu.sink__payload$24[40] ),
    .B(_05594_),
    .Y(_05619_));
 sky130_fd_sc_hd__a211oi_1 _23856_ (.A1(\inst$top.soc.cpu.sink__payload$24[90] ),
    .A2(net1984),
    .B1(net1680),
    .C1(net1160),
    .Y(_05621_));
 sky130_fd_sc_hd__o22ai_4 _23857_ (.A1(_05617_),
    .A2(_05618_),
    .B1(net2204),
    .B2(_05621_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[16] ));
 sky130_fd_sc_hd__inv_1 _23858_ (.A(\inst$top.soc.cpu.sink__payload$12[17] ),
    .Y(_05622_));
 sky130_fd_sc_hd__nand2_1 _23859_ (.A(net2550),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[17] ),
    .Y(_05623_));
 sky130_fd_sc_hd__nand2_1 _23860_ (.A(net2889),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[17] ),
    .Y(_05624_));
 sky130_fd_sc_hd__nand2_1 _23861_ (.A(_05623_),
    .B(_05624_),
    .Y(_05625_));
 sky130_fd_sc_hd__nand2_1 _23862_ (.A(net1830),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__o21ai_0 _23863_ (.A1(_05622_),
    .A2(net1831),
    .B1(_05626_),
    .Y(_05627_));
 sky130_fd_sc_hd__xor2_1 _23865_ (.A(net1978),
    .B(net1299),
    .X(_03206_));
 sky130_fd_sc_hd__inv_2 _23866_ (.A(_03206_),
    .Y(_03210_));
 sky130_fd_sc_hd__inv_1 _23868_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[17] ),
    .Y(_05629_));
 sky130_fd_sc_hd__inv_1 _23869_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie_x_select ),
    .Y(_05630_));
 sky130_fd_sc_hd__inv_1 _23870_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[1] ),
    .Y(_05631_));
 sky130_fd_sc_hd__nand2_1 _23871_ (.A(net2892),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[15] ),
    .Y(_05632_));
 sky130_fd_sc_hd__o221ai_1 _23872_ (.A1(net2213),
    .A2(_05629_),
    .B1(net2194),
    .B2(_05631_),
    .C1(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__a221oi_1 _23873_ (.A1(net2899),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[17] ),
    .B1(net2909),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[15] ),
    .C1(_05633_),
    .Y(_05634_));
 sky130_fd_sc_hd__nand2_1 _23874_ (.A(net2913),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[17] ),
    .Y(_05635_));
 sky130_fd_sc_hd__nand2_1 _23875_ (.A(net2894),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[17] ),
    .Y(_05636_));
 sky130_fd_sc_hd__nand2_1 _23877_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip_x_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[1] ),
    .Y(_05638_));
 sky130_fd_sc_hd__a41oi_1 _23878_ (.A1(_05634_),
    .A2(_05635_),
    .A3(_05636_),
    .A4(_05638_),
    .B1(_20480_),
    .Y(_05639_));
 sky130_fd_sc_hd__inv_1 _23879_ (.A(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__o21ai_1 _23880_ (.A1(net2843),
    .A2(net1720),
    .B1(_05640_),
    .Y(_03205_));
 sky130_fd_sc_hd__inv_2 _23881_ (.A(_03205_),
    .Y(_03209_));
 sky130_fd_sc_hd__nor2_1 _23882_ (.A(\inst$top.soc.cpu.multiplier.w_result[17] ),
    .B(net2198),
    .Y(_05641_));
 sky130_fd_sc_hd__o21ai_0 _23883_ (.A1(net2828),
    .A2(\inst$top.soc.cpu.sink__payload$24[58] ),
    .B1(net2205),
    .Y(_05642_));
 sky130_fd_sc_hd__a211oi_1 _23884_ (.A1(\inst$top.soc.cpu.sink__payload$24[91] ),
    .A2(net1984),
    .B1(net1680),
    .C1(net1160),
    .Y(_05643_));
 sky130_fd_sc_hd__o22ai_4 _23885_ (.A1(_05641_),
    .A2(_05642_),
    .B1(net2205),
    .B2(_05643_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[17] ));
 sky130_fd_sc_hd__inv_1 _23886_ (.A(\inst$top.soc.cpu.sink__payload$12[18] ),
    .Y(_05644_));
 sky130_fd_sc_hd__inv_1 _23887_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[18] ),
    .Y(_05645_));
 sky130_fd_sc_hd__nand2_1 _23888_ (.A(net2546),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[18] ),
    .Y(_05646_));
 sky130_fd_sc_hd__o21ai_0 _23889_ (.A1(net2546),
    .A2(_05645_),
    .B1(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__nand2_1 _23890_ (.A(_05647_),
    .B(net1828),
    .Y(_05648_));
 sky130_fd_sc_hd__o21ai_0 _23891_ (.A1(_05644_),
    .A2(net1831),
    .B1(_05648_),
    .Y(_05649_));
 sky130_fd_sc_hd__xor2_1 _23893_ (.A(net1979),
    .B(net1295),
    .X(_03213_));
 sky130_fd_sc_hd__inv_2 _23894_ (.A(_03213_),
    .Y(_03217_));
 sky130_fd_sc_hd__inv_1 _23895_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[18] ),
    .Y(_05651_));
 sky130_fd_sc_hd__inv_1 _23896_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[2] ),
    .Y(_05652_));
 sky130_fd_sc_hd__o22ai_1 _23897_ (.A1(net2212),
    .A2(_05651_),
    .B1(net2194),
    .B2(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__a21oi_1 _23898_ (.A1(net2892),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[16] ),
    .B1(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__nand2_1 _23899_ (.A(net2909),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[16] ),
    .Y(_05655_));
 sky130_fd_sc_hd__nand2_1 _23900_ (.A(net2899),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[18] ),
    .Y(_05656_));
 sky130_fd_sc_hd__nand3_1 _23901_ (.A(_05654_),
    .B(_05655_),
    .C(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__a21oi_1 _23902_ (.A1(net2913),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[18] ),
    .B1(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__nand2_1 _23903_ (.A(net2905),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[2] ),
    .Y(_05659_));
 sky130_fd_sc_hd__nand2_1 _23904_ (.A(net2894),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[18] ),
    .Y(_05660_));
 sky130_fd_sc_hd__a31o_2 _23905_ (.A1(_05658_),
    .A2(_05659_),
    .A3(_05660_),
    .B1(_20480_),
    .X(_05661_));
 sky130_fd_sc_hd__o21ai_1 _23906_ (.A1(net2848),
    .A2(net1722),
    .B1(_05661_),
    .Y(_03212_));
 sky130_fd_sc_hd__inv_2 _23907_ (.A(_03212_),
    .Y(_03216_));
 sky130_fd_sc_hd__a211oi_1 _23908_ (.A1(\inst$top.soc.cpu.sink__payload$24[92] ),
    .A2(net1982),
    .B1(net1681),
    .C1(net1161),
    .Y(_05662_));
 sky130_fd_sc_hd__nor2_1 _23909_ (.A(net2826),
    .B(\inst$top.soc.cpu.sink__payload$24[59] ),
    .Y(_05663_));
 sky130_fd_sc_hd__nor2_1 _23910_ (.A(\inst$top.soc.cpu.d.sink__payload$16.load ),
    .B(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__o21ai_0 _23911_ (.A1(net2197),
    .A2(\inst$top.soc.cpu.multiplier.w_result[18] ),
    .B1(_05664_),
    .Y(_05665_));
 sky130_fd_sc_hd__o21ai_1 _23912_ (.A1(net2202),
    .A2(_05662_),
    .B1(_05665_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[18] ));
 sky130_fd_sc_hd__inv_1 _23913_ (.A(\inst$top.soc.cpu.sink__payload$12[19] ),
    .Y(_05666_));
 sky130_fd_sc_hd__inv_1 _23914_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[19] ),
    .Y(_05667_));
 sky130_fd_sc_hd__nand2_1 _23915_ (.A(net2547),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[19] ),
    .Y(_05668_));
 sky130_fd_sc_hd__o21ai_0 _23916_ (.A1(net2547),
    .A2(_05667_),
    .B1(_05668_),
    .Y(_05669_));
 sky130_fd_sc_hd__nand2_1 _23917_ (.A(_05669_),
    .B(net1830),
    .Y(_05670_));
 sky130_fd_sc_hd__o21ai_4 _23918_ (.A1(_05666_),
    .A2(net1831),
    .B1(_05670_),
    .Y(_05671_));
 sky130_fd_sc_hd__xor2_1 _23920_ (.A(net1977),
    .B(net1289),
    .X(_03220_));
 sky130_fd_sc_hd__inv_2 _23921_ (.A(_03220_),
    .Y(_03224_));
 sky130_fd_sc_hd__inv_1 _23923_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[3] ),
    .Y(_05674_));
 sky130_fd_sc_hd__nand2_1 _23924_ (.A(net2905),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[3] ),
    .Y(_05675_));
 sky130_fd_sc_hd__nand2_1 _23925_ (.A(net2909),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[17] ),
    .Y(_05676_));
 sky130_fd_sc_hd__nand2_1 _23926_ (.A(net2894),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[19] ),
    .Y(_05677_));
 sky130_fd_sc_hd__o2111ai_1 _23927_ (.A1(net2194),
    .A2(_05674_),
    .B1(_05675_),
    .C1(_05676_),
    .D1(_05677_),
    .Y(_05678_));
 sky130_fd_sc_hd__inv_1 _23928_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[19] ),
    .Y(_05679_));
 sky130_fd_sc_hd__nand2_1 _23929_ (.A(net2913),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[19] ),
    .Y(_05680_));
 sky130_fd_sc_hd__nand2_1 _23930_ (.A(net2899),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[19] ),
    .Y(_05681_));
 sky130_fd_sc_hd__nand2_1 _23931_ (.A(net2892),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[17] ),
    .Y(_05682_));
 sky130_fd_sc_hd__o2111ai_1 _23932_ (.A1(net2212),
    .A2(_05679_),
    .B1(_05680_),
    .C1(_05681_),
    .D1(_05682_),
    .Y(_05683_));
 sky130_fd_sc_hd__o21ai_0 _23933_ (.A1(_05678_),
    .A2(_05683_),
    .B1(net1980),
    .Y(_05684_));
 sky130_fd_sc_hd__o21ai_1 _23934_ (.A1(net2845),
    .A2(_02983_),
    .B1(_05684_),
    .Y(_03219_));
 sky130_fd_sc_hd__inv_2 _23935_ (.A(_03219_),
    .Y(_03223_));
 sky130_fd_sc_hd__nor2_1 _23936_ (.A(\inst$top.soc.cpu.multiplier.w_result[19] ),
    .B(net2198),
    .Y(_05685_));
 sky130_fd_sc_hd__o21ai_0 _23937_ (.A1(net2827),
    .A2(\inst$top.soc.cpu.sink__payload$24[60] ),
    .B1(net2206),
    .Y(_05686_));
 sky130_fd_sc_hd__a211oi_1 _23938_ (.A1(\inst$top.soc.cpu.sink__payload$24[93] ),
    .A2(net1984),
    .B1(net1681),
    .C1(net1162),
    .Y(_05687_));
 sky130_fd_sc_hd__o22ai_2 _23939_ (.A1(_05685_),
    .A2(_05686_),
    .B1(net2206),
    .B2(_05687_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[19] ));
 sky130_fd_sc_hd__inv_1 _23940_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[20] ),
    .Y(_05688_));
 sky130_fd_sc_hd__nand2_1 _23941_ (.A(net2548),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[20] ),
    .Y(_05689_));
 sky130_fd_sc_hd__o21ai_0 _23942_ (.A1(net2548),
    .A2(_05688_),
    .B1(_05689_),
    .Y(_05690_));
 sky130_fd_sc_hd__nand2_1 _23943_ (.A(_05690_),
    .B(net1829),
    .Y(_05691_));
 sky130_fd_sc_hd__nand2_1 _23944_ (.A(_19871_),
    .B(\inst$top.soc.cpu.sink__payload$12[20] ),
    .Y(_05692_));
 sky130_fd_sc_hd__nand2_2 _23945_ (.A(_05691_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__xor2_1 _23946_ (.A(net1977),
    .B(net1286),
    .X(_03227_));
 sky130_fd_sc_hd__inv_2 _23947_ (.A(_03227_),
    .Y(_03231_));
 sky130_fd_sc_hd__inv_1 _23949_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[18] ),
    .Y(_05695_));
 sky130_fd_sc_hd__inv_1 _23950_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[4] ),
    .Y(_05696_));
 sky130_fd_sc_hd__o22ai_1 _23951_ (.A1(net2210),
    .A2(_05695_),
    .B1(_20509_),
    .B2(_05696_),
    .Y(_05697_));
 sky130_fd_sc_hd__inv_1 _23952_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[20] ),
    .Y(_05698_));
 sky130_fd_sc_hd__inv_1 _23953_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[4] ),
    .Y(_05699_));
 sky130_fd_sc_hd__o22ai_1 _23954_ (.A1(net2211),
    .A2(_05698_),
    .B1(net2195),
    .B2(_05699_),
    .Y(_05700_));
 sky130_fd_sc_hd__a21oi_1 _23955_ (.A1(net2900),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[20] ),
    .B1(_05700_),
    .Y(_05701_));
 sky130_fd_sc_hd__nand2_1 _23956_ (.A(net2915),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[20] ),
    .Y(_05702_));
 sky130_fd_sc_hd__nand2_1 _23957_ (.A(net2909),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[18] ),
    .Y(_05703_));
 sky130_fd_sc_hd__nand2_1 _23958_ (.A(net2896),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[20] ),
    .Y(_05704_));
 sky130_fd_sc_hd__nand4_1 _23959_ (.A(_05701_),
    .B(_05702_),
    .C(_05703_),
    .D(_05704_),
    .Y(_05705_));
 sky130_fd_sc_hd__o21ai_1 _23960_ (.A1(_05697_),
    .A2(_05705_),
    .B1(net1980),
    .Y(_05706_));
 sky130_fd_sc_hd__o21ai_1 _23961_ (.A1(net2843),
    .A2(_20003_),
    .B1(_05706_),
    .Y(_03226_));
 sky130_fd_sc_hd__inv_2 _23962_ (.A(_03226_),
    .Y(_03230_));
 sky130_fd_sc_hd__nor2_1 _23963_ (.A(\inst$top.soc.cpu.multiplier.w_result[20] ),
    .B(net2199),
    .Y(_05707_));
 sky130_fd_sc_hd__o21ai_0 _23964_ (.A1(net2828),
    .A2(\inst$top.soc.cpu.sink__payload$24[61] ),
    .B1(net2205),
    .Y(_05708_));
 sky130_fd_sc_hd__a211oi_1 _23965_ (.A1(\inst$top.soc.cpu.sink__payload$24[94] ),
    .A2(net1983),
    .B1(net1680),
    .C1(net1160),
    .Y(_05709_));
 sky130_fd_sc_hd__o22ai_1 _23966_ (.A1(_05707_),
    .A2(_05708_),
    .B1(net2207),
    .B2(_05709_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[20] ));
 sky130_fd_sc_hd__nand2_1 _23967_ (.A(net2548),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[21] ),
    .Y(_05710_));
 sky130_fd_sc_hd__nand2_1 _23968_ (.A(net2889),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[21] ),
    .Y(_05711_));
 sky130_fd_sc_hd__nand2_1 _23969_ (.A(_05710_),
    .B(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__nand2_1 _23970_ (.A(net1829),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__nand2_1 _23971_ (.A(_19871_),
    .B(\inst$top.soc.cpu.sink__payload$12[21] ),
    .Y(_05714_));
 sky130_fd_sc_hd__nand2_1 _23972_ (.A(_05713_),
    .B(_05714_),
    .Y(_05715_));
 sky130_fd_sc_hd__xor2_1 _23973_ (.A(net1979),
    .B(net1281),
    .X(_03234_));
 sky130_fd_sc_hd__inv_2 _23974_ (.A(_03234_),
    .Y(_03238_));
 sky130_fd_sc_hd__inv_1 _23976_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[5] ),
    .Y(_05716_));
 sky130_fd_sc_hd__nand2_1 _23977_ (.A(net2913),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[21] ),
    .Y(_05717_));
 sky130_fd_sc_hd__nand2_1 _23978_ (.A(net2894),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[21] ),
    .Y(_05718_));
 sky130_fd_sc_hd__inv_1 _23979_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[21] ),
    .Y(_05719_));
 sky130_fd_sc_hd__inv_1 _23980_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[5] ),
    .Y(_05720_));
 sky130_fd_sc_hd__nand2_1 _23981_ (.A(net2892),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[19] ),
    .Y(_05721_));
 sky130_fd_sc_hd__o221ai_1 _23982_ (.A1(net2212),
    .A2(_05719_),
    .B1(net2194),
    .B2(_05720_),
    .C1(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__a221oi_1 _23983_ (.A1(net2900),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[21] ),
    .B1(net2909),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[19] ),
    .C1(_05722_),
    .Y(_05723_));
 sky130_fd_sc_hd__o2111ai_1 _23984_ (.A1(_20509_),
    .A2(_05716_),
    .B1(_05717_),
    .C1(_05718_),
    .D1(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__nand2_1 _23985_ (.A(_05724_),
    .B(net1980),
    .Y(_05725_));
 sky130_fd_sc_hd__o21ai_1 _23986_ (.A1(net2848),
    .A2(net1437),
    .B1(_05725_),
    .Y(_03233_));
 sky130_fd_sc_hd__inv_2 _23987_ (.A(_03233_),
    .Y(_03237_));
 sky130_fd_sc_hd__nor2_1 _23988_ (.A(\inst$top.soc.cpu.multiplier.w_result[21] ),
    .B(net2199),
    .Y(_05726_));
 sky130_fd_sc_hd__o21ai_0 _23989_ (.A1(net2828),
    .A2(\inst$top.soc.cpu.sink__payload$24[62] ),
    .B1(net2205),
    .Y(_05727_));
 sky130_fd_sc_hd__a211oi_1 _23990_ (.A1(\inst$top.soc.cpu.sink__payload$24[95] ),
    .A2(net1983),
    .B1(net1680),
    .C1(net1162),
    .Y(_05728_));
 sky130_fd_sc_hd__o22ai_2 _23991_ (.A1(_05726_),
    .A2(_05727_),
    .B1(net2205),
    .B2(_05728_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[21] ));
 sky130_fd_sc_hd__inv_1 _23992_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[22] ),
    .Y(_05729_));
 sky130_fd_sc_hd__nand2_1 _23993_ (.A(net2548),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[22] ),
    .Y(_05730_));
 sky130_fd_sc_hd__o21ai_1 _23994_ (.A1(net2548),
    .A2(_05729_),
    .B1(_05730_),
    .Y(_05731_));
 sky130_fd_sc_hd__a22oi_2 _23995_ (.A1(\inst$top.soc.cpu.sink__payload$12[22] ),
    .A2(_19871_),
    .B1(_05731_),
    .B2(net1828),
    .Y(_05732_));
 sky130_fd_sc_hd__xor2_1 _23997_ (.A(_20373_),
    .B(net1678),
    .X(_03241_));
 sky130_fd_sc_hd__inv_2 _23998_ (.A(_03241_),
    .Y(_03245_));
 sky130_fd_sc_hd__inv_1 _23999_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[20] ),
    .Y(_05734_));
 sky130_fd_sc_hd__inv_1 _24000_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[6] ),
    .Y(_05735_));
 sky130_fd_sc_hd__o22ai_1 _24001_ (.A1(net2208),
    .A2(_05734_),
    .B1(_20509_),
    .B2(_05735_),
    .Y(_05736_));
 sky130_fd_sc_hd__inv_1 _24002_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[22] ),
    .Y(_05737_));
 sky130_fd_sc_hd__inv_1 _24003_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[6] ),
    .Y(_05738_));
 sky130_fd_sc_hd__o22ai_1 _24004_ (.A1(net2212),
    .A2(_05737_),
    .B1(net2195),
    .B2(_05738_),
    .Y(_05739_));
 sky130_fd_sc_hd__a21oi_1 _24005_ (.A1(net2899),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[22] ),
    .B1(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__nand2_1 _24006_ (.A(net2914),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[22] ),
    .Y(_05741_));
 sky130_fd_sc_hd__nand2_1 _24007_ (.A(net2894),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[22] ),
    .Y(_05742_));
 sky130_fd_sc_hd__nand2_1 _24008_ (.A(net2910),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[20] ),
    .Y(_05743_));
 sky130_fd_sc_hd__nand4_1 _24009_ (.A(_05740_),
    .B(_05741_),
    .C(_05742_),
    .D(_05743_),
    .Y(_05744_));
 sky130_fd_sc_hd__o21ai_2 _24010_ (.A1(_05736_),
    .A2(_05744_),
    .B1(net1981),
    .Y(_05745_));
 sky130_fd_sc_hd__o21ai_1 _24011_ (.A1(net2849),
    .A2(net1211),
    .B1(_05745_),
    .Y(_03240_));
 sky130_fd_sc_hd__inv_2 _24012_ (.A(_03240_),
    .Y(_03244_));
 sky130_fd_sc_hd__nor2_1 _24013_ (.A(\inst$top.soc.cpu.multiplier.w_result[22] ),
    .B(net2199),
    .Y(_05746_));
 sky130_fd_sc_hd__o21ai_0 _24014_ (.A1(net2828),
    .A2(\inst$top.soc.cpu.sink__payload$24[63] ),
    .B1(net2207),
    .Y(_05747_));
 sky130_fd_sc_hd__a211oi_1 _24015_ (.A1(\inst$top.soc.cpu.sink__payload$24[96] ),
    .A2(net1984),
    .B1(net1680),
    .C1(net1160),
    .Y(_05748_));
 sky130_fd_sc_hd__o22ai_1 _24016_ (.A1(_05746_),
    .A2(_05747_),
    .B1(net2205),
    .B2(_05748_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[22] ));
 sky130_fd_sc_hd__inv_1 _24017_ (.A(\inst$top.soc.cpu.sink__payload$12[23] ),
    .Y(_05749_));
 sky130_fd_sc_hd__inv_1 _24018_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[23] ),
    .Y(_05750_));
 sky130_fd_sc_hd__nand2_1 _24019_ (.A(net2548),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[23] ),
    .Y(_05751_));
 sky130_fd_sc_hd__o21ai_0 _24020_ (.A1(net2548),
    .A2(_05750_),
    .B1(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__nand2_1 _24021_ (.A(_05752_),
    .B(net1829),
    .Y(_05753_));
 sky130_fd_sc_hd__o21ai_1 _24022_ (.A1(_05749_),
    .A2(net1831),
    .B1(_05753_),
    .Y(_05754_));
 sky130_fd_sc_hd__xor2_1 _24023_ (.A(net1977),
    .B(net1276),
    .X(_03248_));
 sky130_fd_sc_hd__inv_2 _24024_ (.A(_03248_),
    .Y(_03252_));
 sky130_fd_sc_hd__inv_1 _24025_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[7] ),
    .Y(_05755_));
 sky130_fd_sc_hd__nand2_1 _24026_ (.A(net2895),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[23] ),
    .Y(_05756_));
 sky130_fd_sc_hd__nand2_1 _24027_ (.A(net2914),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[23] ),
    .Y(_05757_));
 sky130_fd_sc_hd__inv_1 _24028_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[23] ),
    .Y(_05758_));
 sky130_fd_sc_hd__inv_1 _24029_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[7] ),
    .Y(_05759_));
 sky130_fd_sc_hd__nand2_1 _24030_ (.A(net2892),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[21] ),
    .Y(_05760_));
 sky130_fd_sc_hd__o221ai_1 _24031_ (.A1(net2212),
    .A2(_05758_),
    .B1(net2195),
    .B2(_05759_),
    .C1(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__a221oi_1 _24032_ (.A1(net2899),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[23] ),
    .B1(net2911),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[21] ),
    .C1(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__o2111ai_1 _24033_ (.A1(_20509_),
    .A2(_05755_),
    .B1(_05756_),
    .C1(_05757_),
    .D1(_05762_),
    .Y(_05763_));
 sky130_fd_sc_hd__nand2_1 _24034_ (.A(_05763_),
    .B(net1981),
    .Y(_05764_));
 sky130_fd_sc_hd__o21ai_1 _24035_ (.A1(net2843),
    .A2(net1213),
    .B1(_05764_),
    .Y(_03247_));
 sky130_fd_sc_hd__inv_2 _24036_ (.A(_03247_),
    .Y(_03251_));
 sky130_fd_sc_hd__nor2_1 _24037_ (.A(\inst$top.soc.cpu.multiplier.w_result[23] ),
    .B(net2198),
    .Y(_05765_));
 sky130_fd_sc_hd__o21ai_0 _24038_ (.A1(net2827),
    .A2(\inst$top.soc.cpu.sink__payload$24[64] ),
    .B1(net2206),
    .Y(_05766_));
 sky130_fd_sc_hd__a211oi_1 _24039_ (.A1(\inst$top.soc.cpu.sink__payload$24[97] ),
    .A2(net1984),
    .B1(net1680),
    .C1(net1160),
    .Y(_05767_));
 sky130_fd_sc_hd__o22ai_1 _24040_ (.A1(_05765_),
    .A2(_05766_),
    .B1(net2206),
    .B2(_05767_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[23] ));
 sky130_fd_sc_hd__inv_1 _24041_ (.A(\inst$top.soc.cpu.sink__payload$12[24] ),
    .Y(_05768_));
 sky130_fd_sc_hd__nand2_1 _24042_ (.A(net2548),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[24] ),
    .Y(_05769_));
 sky130_fd_sc_hd__nand2_1 _24043_ (.A(net2888),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[24] ),
    .Y(_05770_));
 sky130_fd_sc_hd__nand2_1 _24044_ (.A(_05769_),
    .B(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__nand2_1 _24045_ (.A(net1829),
    .B(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__o21ai_4 _24046_ (.A1(_05768_),
    .A2(net1831),
    .B1(_05772_),
    .Y(_05773_));
 sky130_fd_sc_hd__xor2_1 _24047_ (.A(net1977),
    .B(net1272),
    .X(_03255_));
 sky130_fd_sc_hd__inv_2 _24048_ (.A(_03255_),
    .Y(_03259_));
 sky130_fd_sc_hd__inv_1 _24051_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[24] ),
    .Y(_05775_));
 sky130_fd_sc_hd__inv_1 _24052_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[8] ),
    .Y(_05776_));
 sky130_fd_sc_hd__o22ai_1 _24053_ (.A1(net2212),
    .A2(_05775_),
    .B1(net2194),
    .B2(_05776_),
    .Y(_05777_));
 sky130_fd_sc_hd__a21oi_1 _24054_ (.A1(net2892),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[22] ),
    .B1(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hd__nand2_1 _24055_ (.A(net2909),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[22] ),
    .Y(_05779_));
 sky130_fd_sc_hd__nand2_1 _24056_ (.A(net2899),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[24] ),
    .Y(_05780_));
 sky130_fd_sc_hd__nand3_1 _24057_ (.A(_05778_),
    .B(_05779_),
    .C(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__a21oi_1 _24058_ (.A1(net2913),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[24] ),
    .B1(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__nand2_1 _24059_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip_x_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[8] ),
    .Y(_05783_));
 sky130_fd_sc_hd__nand2_1 _24060_ (.A(net2894),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[24] ),
    .Y(_05784_));
 sky130_fd_sc_hd__a31o_2 _24061_ (.A1(_05782_),
    .A2(_05783_),
    .A3(_05784_),
    .B1(_20480_),
    .X(_05785_));
 sky130_fd_sc_hd__o21ai_1 _24062_ (.A1(net2844),
    .A2(net1450),
    .B1(_05785_),
    .Y(_03254_));
 sky130_fd_sc_hd__inv_2 _24063_ (.A(_03254_),
    .Y(_03258_));
 sky130_fd_sc_hd__nor2_1 _24064_ (.A(\inst$top.soc.cpu.multiplier.w_result[24] ),
    .B(net2199),
    .Y(_05786_));
 sky130_fd_sc_hd__o21ai_0 _24065_ (.A1(net2828),
    .A2(\inst$top.soc.cpu.sink__payload$24[65] ),
    .B1(net2205),
    .Y(_05787_));
 sky130_fd_sc_hd__a211oi_2 _24066_ (.A1(\inst$top.soc.cpu.sink__payload$24[98] ),
    .A2(net1983),
    .B1(net1680),
    .C1(net1160),
    .Y(_05788_));
 sky130_fd_sc_hd__o22ai_1 _24067_ (.A1(_05786_),
    .A2(_05787_),
    .B1(net2205),
    .B2(_05788_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[24] ));
 sky130_fd_sc_hd__inv_1 _24068_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[25] ),
    .Y(_05789_));
 sky130_fd_sc_hd__nand2_1 _24069_ (.A(net2548),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[25] ),
    .Y(_05790_));
 sky130_fd_sc_hd__o21ai_0 _24070_ (.A1(net2547),
    .A2(_05789_),
    .B1(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hd__a22oi_2 _24071_ (.A1(\inst$top.soc.cpu.sink__payload$12[25] ),
    .A2(_19871_),
    .B1(_05791_),
    .B2(net1828),
    .Y(_05792_));
 sky130_fd_sc_hd__xor2_1 _24073_ (.A(_20373_),
    .B(net1674),
    .X(_03262_));
 sky130_fd_sc_hd__inv_2 _24074_ (.A(_03262_),
    .Y(_03266_));
 sky130_fd_sc_hd__inv_2 _24075_ (.A(net1725),
    .Y(_05794_));
 sky130_fd_sc_hd__inv_1 _24077_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[25] ),
    .Y(_05795_));
 sky130_fd_sc_hd__inv_1 _24078_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[9] ),
    .Y(_05796_));
 sky130_fd_sc_hd__o22ai_1 _24079_ (.A1(net2213),
    .A2(_05795_),
    .B1(net2195),
    .B2(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__a221oi_1 _24080_ (.A1(net2892),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[23] ),
    .B1(net2900),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[25] ),
    .C1(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__nand2_1 _24081_ (.A(net2908),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[23] ),
    .Y(_05799_));
 sky130_fd_sc_hd__nand2_1 _24082_ (.A(net2912),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[25] ),
    .Y(_05800_));
 sky130_fd_sc_hd__nand3_1 _24083_ (.A(_05798_),
    .B(_05799_),
    .C(_05800_),
    .Y(_05801_));
 sky130_fd_sc_hd__a221oi_1 _24084_ (.A1(net2893),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[25] ),
    .B1(net2905),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[9] ),
    .C1(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__nor2_2 _24085_ (.A(_20480_),
    .B(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__inv_1 _24086_ (.A(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__o21ai_1 _24087_ (.A1(net2844),
    .A2(net1268),
    .B1(_05804_),
    .Y(_03261_));
 sky130_fd_sc_hd__inv_2 _24088_ (.A(_03261_),
    .Y(_03265_));
 sky130_fd_sc_hd__nor2_1 _24089_ (.A(\inst$top.soc.cpu.multiplier.w_result[25] ),
    .B(net2198),
    .Y(_05805_));
 sky130_fd_sc_hd__o21ai_0 _24090_ (.A1(net2825),
    .A2(\inst$top.soc.cpu.sink__payload$24[66] ),
    .B1(net2203),
    .Y(_05806_));
 sky130_fd_sc_hd__a211oi_1 _24091_ (.A1(\inst$top.soc.cpu.sink__payload$24[99] ),
    .A2(net1985),
    .B1(net1681),
    .C1(net1161),
    .Y(_05807_));
 sky130_fd_sc_hd__o22ai_1 _24092_ (.A1(_05805_),
    .A2(_05806_),
    .B1(net2203),
    .B2(_05807_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[25] ));
 sky130_fd_sc_hd__nand2_1 _24093_ (.A(net2549),
    .B(\inst$top.soc.cpu.gprf.mem_rp1__data[26] ),
    .Y(_05808_));
 sky130_fd_sc_hd__nand2_1 _24094_ (.A(net2886),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[26] ),
    .Y(_05809_));
 sky130_fd_sc_hd__nand2_1 _24095_ (.A(_05808_),
    .B(_05809_),
    .Y(_05810_));
 sky130_fd_sc_hd__a22oi_2 _24096_ (.A1(\inst$top.soc.cpu.sink__payload$12[26] ),
    .A2(_19871_),
    .B1(net1828),
    .B2(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__xor2_1 _24098_ (.A(_20373_),
    .B(net1670),
    .X(_03269_));
 sky130_fd_sc_hd__inv_2 _24099_ (.A(_03269_),
    .Y(_03273_));
 sky130_fd_sc_hd__inv_2 _24100_ (.A(net1729),
    .Y(_05813_));
 sky130_fd_sc_hd__inv_1 _24102_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[24] ),
    .Y(_05814_));
 sky130_fd_sc_hd__inv_1 _24103_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[10] ),
    .Y(_05815_));
 sky130_fd_sc_hd__o22ai_1 _24104_ (.A1(net2209),
    .A2(_05814_),
    .B1(net2194),
    .B2(_05815_),
    .Y(_05816_));
 sky130_fd_sc_hd__a221oi_1 _24105_ (.A1(net2899),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[26] ),
    .B1(net2909),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[24] ),
    .C1(_05816_),
    .Y(_05817_));
 sky130_fd_sc_hd__nand2_1 _24106_ (.A(net2905),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[10] ),
    .Y(_05818_));
 sky130_fd_sc_hd__nand2_1 _24107_ (.A(net2915),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[26] ),
    .Y(_05819_));
 sky130_fd_sc_hd__nand2_1 _24108_ (.A(net2895),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[26] ),
    .Y(_05820_));
 sky130_fd_sc_hd__nand4_1 _24109_ (.A(_05817_),
    .B(_05818_),
    .C(_05819_),
    .D(_05820_),
    .Y(_05821_));
 sky130_fd_sc_hd__nand2_1 _24110_ (.A(_05821_),
    .B(net1981),
    .Y(_05822_));
 sky130_fd_sc_hd__o21ai_1 _24111_ (.A1(net2849),
    .A2(net1265),
    .B1(_05822_),
    .Y(_03268_));
 sky130_fd_sc_hd__inv_2 _24112_ (.A(_03268_),
    .Y(_03272_));
 sky130_fd_sc_hd__nor2_1 _24113_ (.A(\inst$top.soc.cpu.multiplier.w_result[26] ),
    .B(net2200),
    .Y(_05823_));
 sky130_fd_sc_hd__o21ai_0 _24114_ (.A1(net2825),
    .A2(\inst$top.soc.cpu.sink__payload$24[67] ),
    .B1(net2201),
    .Y(_05824_));
 sky130_fd_sc_hd__a211oi_1 _24115_ (.A1(\inst$top.soc.cpu.sink__payload$24[100] ),
    .A2(net1982),
    .B1(net1681),
    .C1(net1161),
    .Y(_05825_));
 sky130_fd_sc_hd__o22ai_4 _24116_ (.A1(_05823_),
    .A2(_05824_),
    .B1(net2201),
    .B2(_05825_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[26] ));
 sky130_fd_sc_hd__xor2_1 _24117_ (.A(net1977),
    .B(net1453),
    .X(_03276_));
 sky130_fd_sc_hd__inv_2 _24118_ (.A(_03276_),
    .Y(_03280_));
 sky130_fd_sc_hd__inv_2 _24119_ (.A(net1732),
    .Y(_05826_));
 sky130_fd_sc_hd__inv_1 _24121_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[25] ),
    .Y(_05827_));
 sky130_fd_sc_hd__inv_1 _24122_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[11] ),
    .Y(_05828_));
 sky130_fd_sc_hd__o22ai_1 _24123_ (.A1(net2208),
    .A2(_05827_),
    .B1(net2194),
    .B2(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__a221oi_1 _24124_ (.A1(net2899),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[27] ),
    .B1(net2911),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[25] ),
    .C1(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__nand2_1 _24125_ (.A(net2913),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[27] ),
    .Y(_05831_));
 sky130_fd_sc_hd__nand2_1 _24126_ (.A(net2905),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[11] ),
    .Y(_05832_));
 sky130_fd_sc_hd__nand2_1 _24127_ (.A(net2896),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[27] ),
    .Y(_05833_));
 sky130_fd_sc_hd__nand4_1 _24128_ (.A(_05830_),
    .B(_05831_),
    .C(_05832_),
    .D(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__nand2_1 _24129_ (.A(_05834_),
    .B(net1981),
    .Y(_05835_));
 sky130_fd_sc_hd__o21ai_1 _24130_ (.A1(net2843),
    .A2(net1264),
    .B1(_05835_),
    .Y(_03275_));
 sky130_fd_sc_hd__inv_2 _24131_ (.A(_03275_),
    .Y(_03279_));
 sky130_fd_sc_hd__nor2_1 _24132_ (.A(\inst$top.soc.cpu.multiplier.w_result[27] ),
    .B(net2197),
    .Y(_05836_));
 sky130_fd_sc_hd__o21ai_0 _24133_ (.A1(net2826),
    .A2(\inst$top.soc.cpu.sink__payload$24[68] ),
    .B1(net2202),
    .Y(_05837_));
 sky130_fd_sc_hd__a211oi_1 _24134_ (.A1(\inst$top.soc.cpu.sink__payload$24[101] ),
    .A2(net1985),
    .B1(net1681),
    .C1(net1161),
    .Y(_05838_));
 sky130_fd_sc_hd__o22ai_1 _24135_ (.A1(_05836_),
    .A2(_05837_),
    .B1(net2201),
    .B2(_05838_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[27] ));
 sky130_fd_sc_hd__xor2_1 _24136_ (.A(_20373_),
    .B(net1735),
    .X(_03283_));
 sky130_fd_sc_hd__inv_2 _24137_ (.A(_03283_),
    .Y(_03287_));
 sky130_fd_sc_hd__nand2_1 _24138_ (.A(net2913),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[28] ),
    .Y(_05839_));
 sky130_fd_sc_hd__inv_1 _24139_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[26] ),
    .Y(_05840_));
 sky130_fd_sc_hd__inv_1 _24140_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[12] ),
    .Y(_05841_));
 sky130_fd_sc_hd__nand2_1 _24141_ (.A(net2899),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[28] ),
    .Y(_05842_));
 sky130_fd_sc_hd__o221ai_1 _24142_ (.A1(net2209),
    .A2(_05840_),
    .B1(net2194),
    .B2(_05841_),
    .C1(_05842_),
    .Y(_05843_));
 sky130_fd_sc_hd__a21oi_1 _24143_ (.A1(net2909),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[26] ),
    .B1(_05843_),
    .Y(_05844_));
 sky130_fd_sc_hd__nand2_1 _24144_ (.A(net2905),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[12] ),
    .Y(_05845_));
 sky130_fd_sc_hd__nand2_1 _24145_ (.A(net2894),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[28] ),
    .Y(_05846_));
 sky130_fd_sc_hd__a41o_1 _24146_ (.A1(_05839_),
    .A2(_05844_),
    .A3(_05845_),
    .A4(_05846_),
    .B1(_20480_),
    .X(_05847_));
 sky130_fd_sc_hd__o21ai_1 _24147_ (.A1(net2848),
    .A2(net1217),
    .B1(_05847_),
    .Y(_03282_));
 sky130_fd_sc_hd__inv_2 _24148_ (.A(_03282_),
    .Y(_03286_));
 sky130_fd_sc_hd__nor2_1 _24149_ (.A(\inst$top.soc.cpu.multiplier.w_result[28] ),
    .B(net2199),
    .Y(_05848_));
 sky130_fd_sc_hd__o21ai_0 _24150_ (.A1(net2827),
    .A2(\inst$top.soc.cpu.sink__payload$24[69] ),
    .B1(net2207),
    .Y(_05849_));
 sky130_fd_sc_hd__a211oi_1 _24151_ (.A1(\inst$top.soc.cpu.sink__payload$24[102] ),
    .A2(net1983),
    .B1(net1680),
    .C1(net1162),
    .Y(_05850_));
 sky130_fd_sc_hd__o22ai_4 _24152_ (.A1(_05848_),
    .A2(_05849_),
    .B1(net2207),
    .B2(_05850_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[28] ));
 sky130_fd_sc_hd__xor2_1 _24153_ (.A(net1977),
    .B(net1468),
    .X(_03290_));
 sky130_fd_sc_hd__inv_2 _24154_ (.A(_03290_),
    .Y(_03294_));
 sky130_fd_sc_hd__inv_1 _24155_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[13] ),
    .Y(_05851_));
 sky130_fd_sc_hd__nand2_1 _24156_ (.A(net2896),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[29] ),
    .Y(_05852_));
 sky130_fd_sc_hd__inv_1 _24157_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[27] ),
    .Y(_05853_));
 sky130_fd_sc_hd__inv_1 _24158_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[13] ),
    .Y(_05854_));
 sky130_fd_sc_hd__nand2_1 _24159_ (.A(net2898),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[29] ),
    .Y(_05855_));
 sky130_fd_sc_hd__o221ai_1 _24160_ (.A1(net2208),
    .A2(_05853_),
    .B1(net2194),
    .B2(_05854_),
    .C1(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__a221oi_1 _24161_ (.A1(net2913),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[29] ),
    .B1(net2909),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[27] ),
    .C1(_05856_),
    .Y(_05857_));
 sky130_fd_sc_hd__o211ai_1 _24162_ (.A1(_20509_),
    .A2(_05851_),
    .B1(_05852_),
    .C1(_05857_),
    .Y(_05858_));
 sky130_fd_sc_hd__nand2_1 _24163_ (.A(_05858_),
    .B(net1981),
    .Y(_05859_));
 sky130_fd_sc_hd__o21ai_1 _24164_ (.A1(net2844),
    .A2(net1218),
    .B1(_05859_),
    .Y(_03289_));
 sky130_fd_sc_hd__inv_2 _24165_ (.A(_03289_),
    .Y(_03293_));
 sky130_fd_sc_hd__nor2_1 _24166_ (.A(\inst$top.soc.cpu.multiplier.w_result[29] ),
    .B(net2198),
    .Y(_05860_));
 sky130_fd_sc_hd__o21ai_0 _24167_ (.A1(net2827),
    .A2(\inst$top.soc.cpu.sink__payload$24[70] ),
    .B1(net2205),
    .Y(_05861_));
 sky130_fd_sc_hd__a211oi_1 _24168_ (.A1(\inst$top.soc.cpu.sink__payload$24[103] ),
    .A2(net1984),
    .B1(net1680),
    .C1(net1160),
    .Y(_05862_));
 sky130_fd_sc_hd__o22ai_1 _24169_ (.A1(_05860_),
    .A2(_05861_),
    .B1(net2205),
    .B2(_05862_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[29] ));
 sky130_fd_sc_hd__xor2_1 _24170_ (.A(net1977),
    .B(net1475),
    .X(_03297_));
 sky130_fd_sc_hd__inv_2 _24171_ (.A(_03297_),
    .Y(_03301_));
 sky130_fd_sc_hd__inv_1 _24172_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[14] ),
    .Y(_05863_));
 sky130_fd_sc_hd__nand2_1 _24173_ (.A(net2913),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[30] ),
    .Y(_05864_));
 sky130_fd_sc_hd__o21ai_0 _24174_ (.A1(net2194),
    .A2(_05863_),
    .B1(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__inv_1 _24175_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[28] ),
    .Y(_05866_));
 sky130_fd_sc_hd__nand2_1 _24176_ (.A(net2898),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[30] ),
    .Y(_05867_));
 sky130_fd_sc_hd__o21ai_0 _24177_ (.A1(net2208),
    .A2(_05866_),
    .B1(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__nand2_1 _24178_ (.A(net2894),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[30] ),
    .Y(_05869_));
 sky130_fd_sc_hd__nand2_1 _24179_ (.A(net2909),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[28] ),
    .Y(_05870_));
 sky130_fd_sc_hd__nand2_1 _24180_ (.A(net2905),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[14] ),
    .Y(_05871_));
 sky130_fd_sc_hd__nand2_1 _24181_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa_x_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.misa.mxl.x_data[0] ),
    .Y(_05872_));
 sky130_fd_sc_hd__nand4_1 _24182_ (.A(_05869_),
    .B(_05870_),
    .C(_05871_),
    .D(_05872_),
    .Y(_05873_));
 sky130_fd_sc_hd__o31ai_1 _24183_ (.A1(_05865_),
    .A2(_05868_),
    .A3(_05873_),
    .B1(net1981),
    .Y(_05874_));
 sky130_fd_sc_hd__o21ai_1 _24184_ (.A1(net2845),
    .A2(net1219),
    .B1(_05874_),
    .Y(_03296_));
 sky130_fd_sc_hd__inv_2 _24185_ (.A(_03296_),
    .Y(_03300_));
 sky130_fd_sc_hd__nor2_1 _24186_ (.A(\inst$top.soc.cpu.multiplier.w_result[30] ),
    .B(net2198),
    .Y(_05875_));
 sky130_fd_sc_hd__o21ai_0 _24187_ (.A1(net2826),
    .A2(\inst$top.soc.cpu.sink__payload$24[71] ),
    .B1(net2201),
    .Y(_05876_));
 sky130_fd_sc_hd__a211oi_1 _24188_ (.A1(\inst$top.soc.cpu.sink__payload$24[104] ),
    .A2(net1984),
    .B1(net1680),
    .C1(net1162),
    .Y(_05877_));
 sky130_fd_sc_hd__o22ai_1 _24189_ (.A1(_05875_),
    .A2(_05876_),
    .B1(net2201),
    .B2(_05877_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[30] ));
 sky130_fd_sc_hd__xor2_1 _24191_ (.A(net1977),
    .B(net1482),
    .X(_03304_));
 sky130_fd_sc_hd__inv_2 _24192_ (.A(_03304_),
    .Y(_03308_));
 sky130_fd_sc_hd__inv_1 _24194_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa.mxl.x_data[1] ),
    .Y(_05879_));
 sky130_fd_sc_hd__inv_1 _24195_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[29] ),
    .Y(_05880_));
 sky130_fd_sc_hd__nand2_1 _24196_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie_x_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[15] ),
    .Y(_05881_));
 sky130_fd_sc_hd__o221ai_1 _24197_ (.A1(net2211),
    .A2(_05879_),
    .B1(net2210),
    .B2(_05880_),
    .C1(_05881_),
    .Y(_05882_));
 sky130_fd_sc_hd__a221oi_1 _24198_ (.A1(net2897),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[31] ),
    .B1(net2908),
    .B2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[29] ),
    .C1(_05882_),
    .Y(_05883_));
 sky130_fd_sc_hd__nand2_1 _24199_ (.A(net2893),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[31] ),
    .Y(_05884_));
 sky130_fd_sc_hd__nand2_1 _24200_ (.A(net2912),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[31] ),
    .Y(_05885_));
 sky130_fd_sc_hd__nand3_1 _24201_ (.A(_05883_),
    .B(_05884_),
    .C(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__a21oi_1 _24202_ (.A1(net2905),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[15] ),
    .B1(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__o21ai_0 _24204_ (.A1(_20432_),
    .A2(_05887_),
    .B1(net2845),
    .Y(_05889_));
 sky130_fd_sc_hd__o21ai_1 _24205_ (.A1(net2843),
    .A2(net1480),
    .B1(_05889_),
    .Y(_03307_));
 sky130_fd_sc_hd__nor2_1 _24206_ (.A(\inst$top.soc.cpu.multiplier.w_result[31] ),
    .B(net2197),
    .Y(_05890_));
 sky130_fd_sc_hd__o21ai_0 _24207_ (.A1(net2825),
    .A2(\inst$top.soc.cpu.sink__payload$24[72] ),
    .B1(net2203),
    .Y(_05891_));
 sky130_fd_sc_hd__a211oi_1 _24208_ (.A1(\inst$top.soc.cpu.sink__payload$24[105] ),
    .A2(net1982),
    .B1(net1681),
    .C1(net1161),
    .Y(_05892_));
 sky130_fd_sc_hd__o22ai_1 _24209_ (.A1(_05890_),
    .A2(_05891_),
    .B1(net2203),
    .B2(_05892_),
    .Y(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[31] ));
 sky130_fd_sc_hd__nor2_1 _24210_ (.A(net1691),
    .B(net1166),
    .Y(_03367_));
 sky130_fd_sc_hd__inv_2 _24211_ (.A(net1706),
    .Y(_05893_));
 sky130_fd_sc_hd__nand2_1 _24213_ (.A(net1262),
    .B(net1396),
    .Y(_00173_));
 sky130_fd_sc_hd__inv_2 _24214_ (.A(net1694),
    .Y(_03082_));
 sky130_fd_sc_hd__nand2_1 _24215_ (.A(_03082_),
    .B(net1396),
    .Y(_00183_));
 sky130_fd_sc_hd__inv_2 _24216_ (.A(net1356),
    .Y(_05894_));
 sky130_fd_sc_hd__nor2_1 _24217_ (.A(net1181),
    .B(_05894_),
    .Y(_00177_));
 sky130_fd_sc_hd__inv_2 _24219_ (.A(net1351),
    .Y(_05896_));
 sky130_fd_sc_hd__nor2_1 _24220_ (.A(net1697),
    .B(_05896_),
    .Y(_00176_));
 sky130_fd_sc_hd__inv_1 _24221_ (.A(net1350),
    .Y(_05897_));
 sky130_fd_sc_hd__nor2_1 _24223_ (.A(net1683),
    .B(net1159),
    .Y(_00175_));
 sky130_fd_sc_hd__nor2_1 _24224_ (.A(net1707),
    .B(net1173),
    .Y(_03369_));
 sky130_fd_sc_hd__nor2_1 _24225_ (.A(net1691),
    .B(net1196),
    .Y(_03368_));
 sky130_fd_sc_hd__nor2_1 _24226_ (.A(net1173),
    .B(net1692),
    .Y(_03377_));
 sky130_fd_sc_hd__nor2_1 _24227_ (.A(net1707),
    .B(net1683),
    .Y(_02913_));
 sky130_fd_sc_hd__nor2_1 _24228_ (.A(net1691),
    .B(net1698),
    .Y(_02912_));
 sky130_fd_sc_hd__nor2_1 _24229_ (.A(net1691),
    .B(net1163),
    .Y(_03383_));
 sky130_fd_sc_hd__nor2_1 _24230_ (.A(net1707),
    .B(net1166),
    .Y(_03382_));
 sky130_fd_sc_hd__nor2_1 _24232_ (.A(net1366),
    .B(net1170),
    .Y(_00212_));
 sky130_fd_sc_hd__inv_2 _24233_ (.A(net1362),
    .Y(_05900_));
 sky130_fd_sc_hd__nor2_1 _24234_ (.A(net1196),
    .B(_05900_),
    .Y(_00211_));
 sky130_fd_sc_hd__nor2_1 _24235_ (.A(net1173),
    .B(_05894_),
    .Y(_00210_));
 sky130_fd_sc_hd__nor2_1 _24236_ (.A(net1181),
    .B(_05896_),
    .Y(_00217_));
 sky130_fd_sc_hd__nor2_1 _24237_ (.A(net1697),
    .B(net1159),
    .Y(_00216_));
 sky130_fd_sc_hd__inv_1 _24238_ (.A(net1343),
    .Y(_05901_));
 sky130_fd_sc_hd__nor2_1 _24240_ (.A(net1682),
    .B(net1158),
    .Y(_00215_));
 sky130_fd_sc_hd__nor2_1 _24241_ (.A(net1399),
    .B(net1691),
    .Y(_00227_));
 sky130_fd_sc_hd__nor2_1 _24242_ (.A(net1707),
    .B(net1163),
    .Y(_00226_));
 sky130_fd_sc_hd__nor2_1 _24243_ (.A(net1366),
    .B(net1166),
    .Y(_00225_));
 sky130_fd_sc_hd__nor2_1 _24244_ (.A(net1170),
    .B(_05900_),
    .Y(_00229_));
 sky130_fd_sc_hd__nor2_1 _24245_ (.A(net1173),
    .B(_05896_),
    .Y(_00228_));
 sky130_fd_sc_hd__nor2_1 _24246_ (.A(net1181),
    .B(net1159),
    .Y(_00235_));
 sky130_fd_sc_hd__nor2_1 _24247_ (.A(net1697),
    .B(net1158),
    .Y(_00234_));
 sky130_fd_sc_hd__inv_1 _24248_ (.A(net1339),
    .Y(_05903_));
 sky130_fd_sc_hd__nor2_1 _24250_ (.A(net1682),
    .B(net1157),
    .Y(_00233_));
 sky130_fd_sc_hd__nor2_1 _24253_ (.A(net1691),
    .B(_20067_),
    .Y(_03395_));
 sky130_fd_sc_hd__nor2_1 _24254_ (.A(net1706),
    .B(net1399),
    .Y(_00246_));
 sky130_fd_sc_hd__nor2_1 _24255_ (.A(net1366),
    .B(net1163),
    .Y(_00245_));
 sky130_fd_sc_hd__nor2_1 _24256_ (.A(net1166),
    .B(_05900_),
    .Y(_00244_));
 sky130_fd_sc_hd__nor2_1 _24257_ (.A(net1170),
    .B(_05894_),
    .Y(_00249_));
 sky130_fd_sc_hd__nor2_1 _24258_ (.A(net1196),
    .B(_05896_),
    .Y(_00248_));
 sky130_fd_sc_hd__nor2_1 _24259_ (.A(net1173),
    .B(net1159),
    .Y(_00247_));
 sky130_fd_sc_hd__nor2_1 _24260_ (.A(net1181),
    .B(net1158),
    .Y(_00254_));
 sky130_fd_sc_hd__nor2_1 _24261_ (.A(net1697),
    .B(net1157),
    .Y(_00253_));
 sky130_fd_sc_hd__inv_2 _24262_ (.A(net1334),
    .Y(_05907_));
 sky130_fd_sc_hd__nor2_1 _24263_ (.A(net1682),
    .B(_05907_),
    .Y(_00252_));
 sky130_fd_sc_hd__nor2_1 _24264_ (.A(_20061_),
    .B(net1691),
    .Y(_03404_));
 sky130_fd_sc_hd__nor2_1 _24265_ (.A(net1706),
    .B(_20067_),
    .Y(_03403_));
 sky130_fd_sc_hd__nor2_1 _24266_ (.A(net1399),
    .B(net1366),
    .Y(_00270_));
 sky130_fd_sc_hd__nor2_1 _24267_ (.A(net1163),
    .B(_05900_),
    .Y(_00269_));
 sky130_fd_sc_hd__nor2_1 _24268_ (.A(net1166),
    .B(_05894_),
    .Y(_00268_));
 sky130_fd_sc_hd__nor2_1 _24269_ (.A(net1196),
    .B(net1159),
    .Y(_00272_));
 sky130_fd_sc_hd__nor2_1 _24270_ (.A(net1173),
    .B(net1158),
    .Y(_00271_));
 sky130_fd_sc_hd__nor2_1 _24271_ (.A(net1181),
    .B(net1157),
    .Y(_00278_));
 sky130_fd_sc_hd__nor2_1 _24272_ (.A(net1697),
    .B(_05907_),
    .Y(_00277_));
 sky130_fd_sc_hd__inv_1 _24273_ (.A(net1330),
    .Y(_05908_));
 sky130_fd_sc_hd__nor2_1 _24275_ (.A(net1682),
    .B(net1156),
    .Y(_00276_));
 sky130_fd_sc_hd__inv_2 _24276_ (.A(net1366),
    .Y(_05910_));
 sky130_fd_sc_hd__nand2_1 _24279_ (.A(net1153),
    .B(net1403),
    .Y(_00294_));
 sky130_fd_sc_hd__nor2_1 _24280_ (.A(net1399),
    .B(_05900_),
    .Y(_00300_));
 sky130_fd_sc_hd__nor2_1 _24281_ (.A(net1163),
    .B(_05894_),
    .Y(_00299_));
 sky130_fd_sc_hd__nor2_1 _24282_ (.A(net1166),
    .B(_05896_),
    .Y(_00298_));
 sky130_fd_sc_hd__nor2_1 _24283_ (.A(net1170),
    .B(net1159),
    .Y(_00304_));
 sky130_fd_sc_hd__nor2_1 _24284_ (.A(net1196),
    .B(net1158),
    .Y(_00303_));
 sky130_fd_sc_hd__nor2_1 _24285_ (.A(net1173),
    .B(net1157),
    .Y(_00302_));
 sky130_fd_sc_hd__nor2_1 _24286_ (.A(net1181),
    .B(_05907_),
    .Y(_00309_));
 sky130_fd_sc_hd__nor2_1 _24287_ (.A(net1698),
    .B(net1156),
    .Y(_00308_));
 sky130_fd_sc_hd__clkinv_1 _24288_ (.A(net1327),
    .Y(_05912_));
 sky130_fd_sc_hd__nor2_1 _24290_ (.A(net1682),
    .B(net1152),
    .Y(_00307_));
 sky130_fd_sc_hd__nor2_1 _24291_ (.A(net1318),
    .B(net1691),
    .Y(_03416_));
 sky130_fd_sc_hd__nand2_1 _24294_ (.A(net1361),
    .B(net1403),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2_1 _24297_ (.A(net1357),
    .B(_03045_),
    .Y(_00324_));
 sky130_fd_sc_hd__nor2_1 _24298_ (.A(net1172),
    .B(net1158),
    .Y(_00331_));
 sky130_fd_sc_hd__nor2_1 _24299_ (.A(net1197),
    .B(net1157),
    .Y(_00330_));
 sky130_fd_sc_hd__nor2_1 _24300_ (.A(net1173),
    .B(_05907_),
    .Y(_00329_));
 sky130_fd_sc_hd__nor2_1 _24301_ (.A(net1181),
    .B(net1156),
    .Y(_00336_));
 sky130_fd_sc_hd__nor2_1 _24302_ (.A(net1697),
    .B(net1152),
    .Y(_00335_));
 sky130_fd_sc_hd__clkinv_1 _24303_ (.A(net1322),
    .Y(_05916_));
 sky130_fd_sc_hd__nor2_1 _24305_ (.A(net1682),
    .B(net1150),
    .Y(_00334_));
 sky130_fd_sc_hd__nor2_1 _24306_ (.A(net1692),
    .B(_03017_),
    .Y(_03422_));
 sky130_fd_sc_hd__nor2_1 _24307_ (.A(net1706),
    .B(net1318),
    .Y(_03421_));
 sky130_fd_sc_hd__nand2_1 _24308_ (.A(net1357),
    .B(net1403),
    .Y(_00346_));
 sky130_fd_sc_hd__nor2_1 _24309_ (.A(net1399),
    .B(_05896_),
    .Y(_00352_));
 sky130_fd_sc_hd__nor2_1 _24310_ (.A(net1163),
    .B(net1159),
    .Y(_00351_));
 sky130_fd_sc_hd__nor2_1 _24311_ (.A(net1166),
    .B(net1158),
    .Y(_00350_));
 sky130_fd_sc_hd__nor2_1 _24312_ (.A(net1170),
    .B(net1157),
    .Y(_00363_));
 sky130_fd_sc_hd__nor2_1 _24313_ (.A(net1197),
    .B(_05907_),
    .Y(_00362_));
 sky130_fd_sc_hd__nor2_1 _24314_ (.A(net1173),
    .B(net1156),
    .Y(_00361_));
 sky130_fd_sc_hd__nor2_1 _24317_ (.A(net1182),
    .B(net1152),
    .Y(_00368_));
 sky130_fd_sc_hd__nor2_1 _24318_ (.A(net1697),
    .B(net1150),
    .Y(_00367_));
 sky130_fd_sc_hd__inv_1 _24319_ (.A(net1317),
    .Y(_05920_));
 sky130_fd_sc_hd__nor2_1 _24321_ (.A(net1682),
    .B(net1148),
    .Y(_00366_));
 sky130_fd_sc_hd__nand2_1 _24323_ (.A(net1403),
    .B(net1351),
    .Y(_00383_));
 sky130_fd_sc_hd__nor2_1 _24324_ (.A(net1399),
    .B(_05897_),
    .Y(_00390_));
 sky130_fd_sc_hd__nor2_1 _24326_ (.A(net1166),
    .B(net1157),
    .Y(_00389_));
 sky130_fd_sc_hd__nor2_1 _24327_ (.A(net1170),
    .B(_05907_),
    .Y(_00403_));
 sky130_fd_sc_hd__nor2_1 _24328_ (.A(net1197),
    .B(net1156),
    .Y(_00402_));
 sky130_fd_sc_hd__nor2_1 _24330_ (.A(net1174),
    .B(net1152),
    .Y(_00401_));
 sky130_fd_sc_hd__nor2_1 _24331_ (.A(net1182),
    .B(net1150),
    .Y(_00408_));
 sky130_fd_sc_hd__nor2_1 _24333_ (.A(net1698),
    .B(net1148),
    .Y(_00407_));
 sky130_fd_sc_hd__inv_1 _24336_ (.A(net1312),
    .Y(_05928_));
 sky130_fd_sc_hd__nor2_1 _24338_ (.A(net1683),
    .B(net1145),
    .Y(_00406_));
 sky130_fd_sc_hd__nor2_1 _24339_ (.A(net1693),
    .B(net1713),
    .Y(_03435_));
 sky130_fd_sc_hd__nand2_1 _24341_ (.A(net1262),
    .B(net1424),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _24344_ (.A(net1155),
    .B(net1420),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2_1 _24345_ (.A(net1362),
    .B(net1415),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_1 _24346_ (.A(net1357),
    .B(net1411),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _24347_ (.A(_20062_),
    .B(net1351),
    .Y(_00424_));
 sky130_fd_sc_hd__nand2_1 _24349_ (.A(net1406),
    .B(net1350),
    .Y(_00423_));
 sky130_fd_sc_hd__nand2_1 _24351_ (.A(net1337),
    .B(net1397),
    .Y(_00428_));
 sky130_fd_sc_hd__nor2_1 _24352_ (.A(net1170),
    .B(net1156),
    .Y(_00434_));
 sky130_fd_sc_hd__nor2_1 _24353_ (.A(net1197),
    .B(net1152),
    .Y(_00433_));
 sky130_fd_sc_hd__nor2_1 _24354_ (.A(net1174),
    .B(net1150),
    .Y(_00432_));
 sky130_fd_sc_hd__nor2_1 _24355_ (.A(net1181),
    .B(net1148),
    .Y(_00439_));
 sky130_fd_sc_hd__nor2_1 _24356_ (.A(net1698),
    .B(net1145),
    .Y(_00438_));
 sky130_fd_sc_hd__inv_1 _24357_ (.A(net1308),
    .Y(_05931_));
 sky130_fd_sc_hd__nor2_1 _24359_ (.A(net1683),
    .B(net1143),
    .Y(_00437_));
 sky130_fd_sc_hd__nor2_1 _24360_ (.A(net1693),
    .B(net1716),
    .Y(_03445_));
 sky130_fd_sc_hd__nor2_1 _24362_ (.A(net1707),
    .B(net1713),
    .Y(_03444_));
 sky130_fd_sc_hd__nand2_1 _24363_ (.A(net1153),
    .B(net1424),
    .Y(_00457_));
 sky130_fd_sc_hd__nand2_1 _24364_ (.A(net1362),
    .B(net1420),
    .Y(_00456_));
 sky130_fd_sc_hd__nand2_1 _24365_ (.A(net1357),
    .B(net1415),
    .Y(_00455_));
 sky130_fd_sc_hd__nand2_1 _24367_ (.A(net1355),
    .B(net1411),
    .Y(_00460_));
 sky130_fd_sc_hd__nand2_1 _24369_ (.A(net1203),
    .B(net1350),
    .Y(_00459_));
 sky130_fd_sc_hd__nand2_1 _24371_ (.A(net1406),
    .B(net1346),
    .Y(_00458_));
 sky130_fd_sc_hd__nand2_1 _24373_ (.A(net1331),
    .B(net1397),
    .Y(_00462_));
 sky130_fd_sc_hd__nand2_1 _24375_ (.A(net1317),
    .B(net1394),
    .Y(_00466_));
 sky130_fd_sc_hd__nor2_1 _24376_ (.A(net1183),
    .B(net1145),
    .Y(_00471_));
 sky130_fd_sc_hd__nor2_1 _24377_ (.A(net1698),
    .B(net1143),
    .Y(_00470_));
 sky130_fd_sc_hd__inv_1 _24378_ (.A(net1300),
    .Y(_05935_));
 sky130_fd_sc_hd__nor2_1 _24380_ (.A(net1684),
    .B(net1142),
    .Y(_00469_));
 sky130_fd_sc_hd__inv_2 _24381_ (.A(_00485_),
    .Y(_00482_));
 sky130_fd_sc_hd__nor2_1 _24382_ (.A(net1693),
    .B(net1720),
    .Y(_00488_));
 sky130_fd_sc_hd__nor2_1 _24383_ (.A(net1707),
    .B(net1716),
    .Y(_00487_));
 sky130_fd_sc_hd__nor2_1 _24384_ (.A(net1713),
    .B(net1368),
    .Y(_00486_));
 sky130_fd_sc_hd__nand2_1 _24385_ (.A(net1362),
    .B(net1424),
    .Y(_00491_));
 sky130_fd_sc_hd__nand2_1 _24386_ (.A(net1360),
    .B(net1420),
    .Y(_00490_));
 sky130_fd_sc_hd__nand2_1 _24387_ (.A(net1354),
    .B(net1415),
    .Y(_00489_));
 sky130_fd_sc_hd__nand2_1 _24388_ (.A(net1349),
    .B(net1411),
    .Y(_00494_));
 sky130_fd_sc_hd__nand2_1 _24389_ (.A(net1203),
    .B(net1344),
    .Y(_00493_));
 sky130_fd_sc_hd__nand2_1 _24391_ (.A(net1403),
    .B(net1341),
    .Y(_00492_));
 sky130_fd_sc_hd__nor2_1 _24392_ (.A(net1163),
    .B(net1156),
    .Y(_00497_));
 sky130_fd_sc_hd__nor2_1 _24393_ (.A(net1169),
    .B(net1152),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_1 _24395_ (.A(net1311),
    .B(net1394),
    .Y(_00502_));
 sky130_fd_sc_hd__nor2_1 _24396_ (.A(net1183),
    .B(net1144),
    .Y(_00507_));
 sky130_fd_sc_hd__nor2_1 _24397_ (.A(net1699),
    .B(net1142),
    .Y(_00506_));
 sky130_fd_sc_hd__inv_1 _24398_ (.A(net1299),
    .Y(_05938_));
 sky130_fd_sc_hd__nor2_1 _24400_ (.A(net1684),
    .B(net1139),
    .Y(_00505_));
 sky130_fd_sc_hd__inv_2 _24401_ (.A(_00522_),
    .Y(_00518_));
 sky130_fd_sc_hd__nor2_1 _24402_ (.A(net1693),
    .B(net1722),
    .Y(_03466_));
 sky130_fd_sc_hd__nor2_1 _24403_ (.A(net1708),
    .B(net1721),
    .Y(_00525_));
 sky130_fd_sc_hd__nor2_1 _24404_ (.A(net1368),
    .B(net1716),
    .Y(_00524_));
 sky130_fd_sc_hd__nor2_1 _24405_ (.A(net1712),
    .B(_05900_),
    .Y(_00523_));
 sky130_fd_sc_hd__nand2_1 _24406_ (.A(net1360),
    .B(net1424),
    .Y(_00528_));
 sky130_fd_sc_hd__nand2_1 _24407_ (.A(net1354),
    .B(net1420),
    .Y(_00527_));
 sky130_fd_sc_hd__nand2_1 _24408_ (.A(net1349),
    .B(net1415),
    .Y(_00526_));
 sky130_fd_sc_hd__nor2_1 _24409_ (.A(net1163),
    .B(net1152),
    .Y(_00538_));
 sky130_fd_sc_hd__nor2_1 _24410_ (.A(net1169),
    .B(net1150),
    .Y(_00537_));
 sky130_fd_sc_hd__nand2_1 _24412_ (.A(net1307),
    .B(net1394),
    .Y(_00544_));
 sky130_fd_sc_hd__nor2_1 _24413_ (.A(net1183),
    .B(net1142),
    .Y(_00549_));
 sky130_fd_sc_hd__nor2_1 _24414_ (.A(net1699),
    .B(net1139),
    .Y(_00548_));
 sky130_fd_sc_hd__inv_1 _24415_ (.A(net1295),
    .Y(_05940_));
 sky130_fd_sc_hd__nor2_1 _24417_ (.A(net1684),
    .B(net1137),
    .Y(_00547_));
 sky130_fd_sc_hd__inv_2 _24418_ (.A(_00565_),
    .Y(_00561_));
 sky130_fd_sc_hd__nor2_1 _24419_ (.A(net1695),
    .B(_02983_),
    .Y(_03478_));
 sky130_fd_sc_hd__nor2_1 _24420_ (.A(net1708),
    .B(net1722),
    .Y(_03477_));
 sky130_fd_sc_hd__nand2_1 _24421_ (.A(net1360),
    .B(net1425),
    .Y(_00566_));
 sky130_fd_sc_hd__nand2_1 _24422_ (.A(net1354),
    .B(net1423),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _24423_ (.A(net1349),
    .B(net1419),
    .Y(_00572_));
 sky130_fd_sc_hd__nand2_1 _24424_ (.A(net1344),
    .B(net1415),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _24426_ (.A(net1340),
    .B(net1411),
    .Y(_00576_));
 sky130_fd_sc_hd__nand2_1 _24428_ (.A(net1203),
    .B(net1335),
    .Y(_00575_));
 sky130_fd_sc_hd__nand2_1 _24429_ (.A(net1403),
    .B(net1330),
    .Y(_00574_));
 sky130_fd_sc_hd__nor2_1 _24432_ (.A(_20630_),
    .B(net1150),
    .Y(_00580_));
 sky130_fd_sc_hd__nor2_1 _24433_ (.A(net1169),
    .B(net1149),
    .Y(_00579_));
 sky130_fd_sc_hd__nand2_1 _24435_ (.A(net1302),
    .B(net1394),
    .Y(_00587_));
 sky130_fd_sc_hd__nor2_1 _24436_ (.A(net1183),
    .B(_05938_),
    .Y(_00592_));
 sky130_fd_sc_hd__nor2_1 _24437_ (.A(net1699),
    .B(net1138),
    .Y(_00591_));
 sky130_fd_sc_hd__clkinv_1 _24438_ (.A(net1287),
    .Y(_05945_));
 sky130_fd_sc_hd__nor2_1 _24440_ (.A(net1684),
    .B(net3042),
    .Y(_00590_));
 sky130_fd_sc_hd__inv_2 _24441_ (.A(_00610_),
    .Y(_00607_));
 sky130_fd_sc_hd__inv_2 _24442_ (.A(_20003_),
    .Y(_05947_));
 sky130_fd_sc_hd__nand2_1 _24444_ (.A(net1134),
    .B(_03082_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand2_1 _24446_ (.A(net1263),
    .B(net1434),
    .Y(_00612_));
 sky130_fd_sc_hd__nand2_1 _24447_ (.A(net1431),
    .B(net1155),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _24448_ (.A(net1428),
    .B(net1365),
    .Y(_00617_));
 sky130_fd_sc_hd__nand2_1 _24449_ (.A(net1427),
    .B(net1360),
    .Y(_00616_));
 sky130_fd_sc_hd__nand2_1 _24450_ (.A(net1425),
    .B(net1354),
    .Y(_00615_));
 sky130_fd_sc_hd__nand2_1 _24451_ (.A(net1349),
    .B(net1423),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _24452_ (.A(net1344),
    .B(net1419),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _24453_ (.A(net1340),
    .B(net1414),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _24455_ (.A(net1405),
    .B(net1326),
    .Y(_00625_));
 sky130_fd_sc_hd__nor2_1 _24456_ (.A(net1165),
    .B(net1149),
    .Y(_00631_));
 sky130_fd_sc_hd__nor2_1 _24457_ (.A(net1169),
    .B(net1147),
    .Y(_00630_));
 sky130_fd_sc_hd__nand2_1 _24459_ (.A(net1296),
    .B(net1393),
    .Y(_00637_));
 sky130_fd_sc_hd__nor2_1 _24460_ (.A(net1183),
    .B(_05940_),
    .Y(_00642_));
 sky130_fd_sc_hd__nor2_1 _24461_ (.A(net1699),
    .B(net3042),
    .Y(_00641_));
 sky130_fd_sc_hd__inv_2 _24462_ (.A(net1286),
    .Y(_05948_));
 sky130_fd_sc_hd__nor2_1 _24464_ (.A(net1684),
    .B(net1131),
    .Y(_00640_));
 sky130_fd_sc_hd__inv_2 _24465_ (.A(_00660_),
    .Y(_00657_));
 sky130_fd_sc_hd__nor2_1 _24466_ (.A(net1695),
    .B(net1439),
    .Y(_03498_));
 sky130_fd_sc_hd__nand2_1 _24467_ (.A(net1134),
    .B(net1263),
    .Y(_00663_));
 sky130_fd_sc_hd__nand2_1 _24468_ (.A(net1154),
    .B(net1434),
    .Y(_00662_));
 sky130_fd_sc_hd__nand2_1 _24469_ (.A(net1431),
    .B(net1364),
    .Y(_00661_));
 sky130_fd_sc_hd__nand2_1 _24470_ (.A(net1428),
    .B(net1359),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_1 _24471_ (.A(net1427),
    .B(net1354),
    .Y(_00666_));
 sky130_fd_sc_hd__nand2_1 _24472_ (.A(net1425),
    .B(net1349),
    .Y(_00665_));
 sky130_fd_sc_hd__nand2_1 _24473_ (.A(net1344),
    .B(net1423),
    .Y(_00671_));
 sky130_fd_sc_hd__nand2_1 _24474_ (.A(net1340),
    .B(net1419),
    .Y(_00670_));
 sky130_fd_sc_hd__nand2_1 _24475_ (.A(net1335),
    .B(net1414),
    .Y(_00669_));
 sky130_fd_sc_hd__nand2_1 _24476_ (.A(net1330),
    .B(net1410),
    .Y(_00674_));
 sky130_fd_sc_hd__nand2_1 _24477_ (.A(net1206),
    .B(net1326),
    .Y(_00673_));
 sky130_fd_sc_hd__nand2_1 _24479_ (.A(net1405),
    .B(net1321),
    .Y(_00672_));
 sky130_fd_sc_hd__nor2_1 _24480_ (.A(net1165),
    .B(net1147),
    .Y(_00679_));
 sky130_fd_sc_hd__nor2_1 _24481_ (.A(net1167),
    .B(_05931_),
    .Y(_00678_));
 sky130_fd_sc_hd__nand2_1 _24483_ (.A(net1292),
    .B(net1393),
    .Y(_00685_));
 sky130_fd_sc_hd__nor2_1 _24484_ (.A(net1190),
    .B(net3042),
    .Y(_00690_));
 sky130_fd_sc_hd__nor2_1 _24485_ (.A(net1705),
    .B(net1129),
    .Y(_00689_));
 sky130_fd_sc_hd__inv_2 _24486_ (.A(net1280),
    .Y(_05950_));
 sky130_fd_sc_hd__nor2_1 _24488_ (.A(net1689),
    .B(net1126),
    .Y(_00688_));
 sky130_fd_sc_hd__inv_2 _24489_ (.A(_00708_),
    .Y(_00705_));
 sky130_fd_sc_hd__nor2_1 _24490_ (.A(net1695),
    .B(_19992_),
    .Y(_03510_));
 sky130_fd_sc_hd__nor2_1 _24491_ (.A(_20124_),
    .B(net1439),
    .Y(_03509_));
 sky130_fd_sc_hd__nand2_1 _24493_ (.A(net1154),
    .B(net1133),
    .Y(_00711_));
 sky130_fd_sc_hd__nand2_1 _24494_ (.A(net1363),
    .B(net1433),
    .Y(_00710_));
 sky130_fd_sc_hd__nand2_1 _24495_ (.A(net1430),
    .B(net1358),
    .Y(_00709_));
 sky130_fd_sc_hd__nand2_1 _24496_ (.A(_20019_),
    .B(net1353),
    .Y(_00715_));
 sky130_fd_sc_hd__nand2_1 _24497_ (.A(_20024_),
    .B(net1348),
    .Y(_00714_));
 sky130_fd_sc_hd__nand2_1 _24499_ (.A(net1426),
    .B(net1344),
    .Y(_00713_));
 sky130_fd_sc_hd__nand2_1 _24500_ (.A(net1340),
    .B(net1423),
    .Y(_00719_));
 sky130_fd_sc_hd__nand2_1 _24501_ (.A(net1335),
    .B(net1419),
    .Y(_00718_));
 sky130_fd_sc_hd__nand2_1 _24502_ (.A(net1330),
    .B(net1414),
    .Y(_00717_));
 sky130_fd_sc_hd__nand2_1 _24504_ (.A(net1405),
    .B(net1316),
    .Y(_00720_));
 sky130_fd_sc_hd__nor2_1 _24505_ (.A(net1165),
    .B(net1144),
    .Y(_00729_));
 sky130_fd_sc_hd__nor2_1 _24506_ (.A(net1167),
    .B(_05935_),
    .Y(_00728_));
 sky130_fd_sc_hd__nand2_1 _24508_ (.A(net1288),
    .B(net1393),
    .Y(_00735_));
 sky130_fd_sc_hd__nor2_1 _24509_ (.A(net1129),
    .B(net1190),
    .Y(_00740_));
 sky130_fd_sc_hd__nor2_1 _24510_ (.A(net1705),
    .B(net1126),
    .Y(_00739_));
 sky130_fd_sc_hd__nor2_1 _24512_ (.A(net1686),
    .B(net1677),
    .Y(_00738_));
 sky130_fd_sc_hd__inv_2 _24513_ (.A(_00756_),
    .Y(_00753_));
 sky130_fd_sc_hd__nand2_1 _24514_ (.A(net1133),
    .B(net1363),
    .Y(_00764_));
 sky130_fd_sc_hd__nand2_1 _24515_ (.A(net1358),
    .B(net1433),
    .Y(_00763_));
 sky130_fd_sc_hd__nand2_1 _24516_ (.A(net1430),
    .B(net1353),
    .Y(_00762_));
 sky130_fd_sc_hd__nand2_1 _24517_ (.A(_20019_),
    .B(net1348),
    .Y(_00771_));
 sky130_fd_sc_hd__nand2_1 _24518_ (.A(_20024_),
    .B(net1342),
    .Y(_00770_));
 sky130_fd_sc_hd__nand2_1 _24519_ (.A(net1426),
    .B(net1339),
    .Y(_00769_));
 sky130_fd_sc_hd__nand2_1 _24522_ (.A(net1334),
    .B(net1423),
    .Y(_00774_));
 sky130_fd_sc_hd__nand2_1 _24524_ (.A(net1330),
    .B(net1419),
    .Y(_00773_));
 sky130_fd_sc_hd__nand2_1 _24526_ (.A(net1326),
    .B(net1414),
    .Y(_00772_));
 sky130_fd_sc_hd__nand2_1 _24527_ (.A(net1321),
    .B(net1410),
    .Y(_00777_));
 sky130_fd_sc_hd__nand2_1 _24528_ (.A(net1206),
    .B(net1316),
    .Y(_00776_));
 sky130_fd_sc_hd__nand2_1 _24530_ (.A(net1405),
    .B(net1311),
    .Y(_00775_));
 sky130_fd_sc_hd__nor2_1 _24531_ (.A(net1165),
    .B(_05935_),
    .Y(_00783_));
 sky130_fd_sc_hd__nor2_1 _24532_ (.A(net1167),
    .B(_05938_),
    .Y(_00782_));
 sky130_fd_sc_hd__nand2_1 _24535_ (.A(net1283),
    .B(net1393),
    .Y(_00789_));
 sky130_fd_sc_hd__nor2_1 _24536_ (.A(net1126),
    .B(net1190),
    .Y(_00794_));
 sky130_fd_sc_hd__nor2_1 _24537_ (.A(net1700),
    .B(net1677),
    .Y(_00793_));
 sky130_fd_sc_hd__inv_2 _24538_ (.A(net1276),
    .Y(_05962_));
 sky130_fd_sc_hd__nor2_1 _24540_ (.A(net1686),
    .B(net1123),
    .Y(_00792_));
 sky130_fd_sc_hd__inv_2 _24541_ (.A(_00811_),
    .Y(_00808_));
 sky130_fd_sc_hd__nor2_1 _24542_ (.A(net1694),
    .B(net1451),
    .Y(_03537_));
 sky130_fd_sc_hd__nand2_1 _24545_ (.A(net1263),
    .B(net1446),
    .Y(_00814_));
 sky130_fd_sc_hd__nand2_1 _24547_ (.A(net1154),
    .B(net1442),
    .Y(_00813_));
 sky130_fd_sc_hd__nand2_1 _24548_ (.A(net1363),
    .B(net1210),
    .Y(_00812_));
 sky130_fd_sc_hd__nand2_1 _24549_ (.A(net1133),
    .B(net1358),
    .Y(_00817_));
 sky130_fd_sc_hd__nand2_1 _24550_ (.A(net1353),
    .B(net1433),
    .Y(_00816_));
 sky130_fd_sc_hd__nand2_1 _24551_ (.A(net1430),
    .B(net1349),
    .Y(_00815_));
 sky130_fd_sc_hd__nand2_1 _24552_ (.A(_20019_),
    .B(net1342),
    .Y(_00823_));
 sky130_fd_sc_hd__nand2_1 _24553_ (.A(net1427),
    .B(net1339),
    .Y(_00822_));
 sky130_fd_sc_hd__nand2_1 _24554_ (.A(net1425),
    .B(net1333),
    .Y(_00821_));
 sky130_fd_sc_hd__nand2_1 _24555_ (.A(net1316),
    .B(net1410),
    .Y(_00831_));
 sky130_fd_sc_hd__nand2_1 _24556_ (.A(net1206),
    .B(net1311),
    .Y(_00830_));
 sky130_fd_sc_hd__nand2_1 _24559_ (.A(net1405),
    .B(net1307),
    .Y(_00829_));
 sky130_fd_sc_hd__nor2_1 _24560_ (.A(net1165),
    .B(net1140),
    .Y(_00837_));
 sky130_fd_sc_hd__nor2_1 _24561_ (.A(net1167),
    .B(_05940_),
    .Y(_00836_));
 sky130_fd_sc_hd__nand2_1 _24563_ (.A(net1278),
    .B(net1392),
    .Y(_00843_));
 sky130_fd_sc_hd__nor2_1 _24564_ (.A(net1189),
    .B(net1677),
    .Y(_00848_));
 sky130_fd_sc_hd__nor2_1 _24566_ (.A(net1701),
    .B(net1123),
    .Y(_00847_));
 sky130_fd_sc_hd__inv_2 _24567_ (.A(net1270),
    .Y(_05968_));
 sky130_fd_sc_hd__nor2_1 _24569_ (.A(net1689),
    .B(net1121),
    .Y(_00846_));
 sky130_fd_sc_hd__inv_2 _24570_ (.A(_00868_),
    .Y(_00865_));
 sky130_fd_sc_hd__nor2_1 _24571_ (.A(net1694),
    .B(net1269),
    .Y(_03548_));
 sky130_fd_sc_hd__nor2_1 _24572_ (.A(_20124_),
    .B(net1451),
    .Y(_03547_));
 sky130_fd_sc_hd__nand2_1 _24573_ (.A(net1154),
    .B(net1446),
    .Y(_00871_));
 sky130_fd_sc_hd__nand2_1 _24574_ (.A(net1363),
    .B(net1442),
    .Y(_00870_));
 sky130_fd_sc_hd__nand2_1 _24575_ (.A(net1358),
    .B(net1209),
    .Y(_00869_));
 sky130_fd_sc_hd__nand2_1 _24576_ (.A(net1133),
    .B(net1352),
    .Y(_00874_));
 sky130_fd_sc_hd__nand2_1 _24577_ (.A(net1348),
    .B(net1433),
    .Y(_00873_));
 sky130_fd_sc_hd__nand2_1 _24578_ (.A(net1430),
    .B(net1342),
    .Y(_00872_));
 sky130_fd_sc_hd__nand2_1 _24579_ (.A(net1428),
    .B(net1339),
    .Y(_00879_));
 sky130_fd_sc_hd__nand2_1 _24580_ (.A(net1427),
    .B(net1332),
    .Y(_00878_));
 sky130_fd_sc_hd__nand2_1 _24582_ (.A(net1425),
    .B(net1329),
    .Y(_00877_));
 sky130_fd_sc_hd__nand2_1 _24583_ (.A(net1325),
    .B(net1423),
    .Y(_00882_));
 sky130_fd_sc_hd__nand2_1 _24584_ (.A(net1320),
    .B(net1419),
    .Y(_00881_));
 sky130_fd_sc_hd__nand2_1 _24585_ (.A(net1315),
    .B(net1414),
    .Y(_00880_));
 sky130_fd_sc_hd__nand2_1 _24586_ (.A(net1310),
    .B(net1410),
    .Y(_00885_));
 sky130_fd_sc_hd__nand2_1 _24587_ (.A(net1206),
    .B(net1306),
    .Y(_00884_));
 sky130_fd_sc_hd__nand2_1 _24589_ (.A(net1405),
    .B(net1302),
    .Y(_00883_));
 sky130_fd_sc_hd__nor2_1 _24590_ (.A(net1165),
    .B(_05940_),
    .Y(_00894_));
 sky130_fd_sc_hd__nor2_1 _24591_ (.A(net1167),
    .B(net3042),
    .Y(_00893_));
 sky130_fd_sc_hd__inv_1 _24592_ (.A(net1678),
    .Y(_05972_));
 sky130_fd_sc_hd__nand2_1 _24595_ (.A(net1258),
    .B(net1392),
    .Y(_00900_));
 sky130_fd_sc_hd__nor2_1 _24596_ (.A(net1189),
    .B(net1123),
    .Y(_00905_));
 sky130_fd_sc_hd__nor2_1 _24597_ (.A(net1700),
    .B(net1121),
    .Y(_00904_));
 sky130_fd_sc_hd__nor2_1 _24599_ (.A(net1685),
    .B(net1672),
    .Y(_00903_));
 sky130_fd_sc_hd__inv_2 _24600_ (.A(_00924_),
    .Y(_00921_));
 sky130_fd_sc_hd__nor2_1 _24601_ (.A(net1708),
    .B(net1267),
    .Y(_00926_));
 sky130_fd_sc_hd__nor2_1 _24602_ (.A(net1451),
    .B(net1368),
    .Y(_00925_));
 sky130_fd_sc_hd__nand2_1 _24603_ (.A(net1363),
    .B(net1444),
    .Y(_00930_));
 sky130_fd_sc_hd__nand2_1 _24605_ (.A(net1358),
    .B(net1440),
    .Y(_00929_));
 sky130_fd_sc_hd__nand2_1 _24606_ (.A(net1207),
    .B(net1352),
    .Y(_00928_));
 sky130_fd_sc_hd__nand2_1 _24607_ (.A(net1133),
    .B(net1348),
    .Y(_00933_));
 sky130_fd_sc_hd__nand2_1 _24608_ (.A(net1343),
    .B(net1433),
    .Y(_00932_));
 sky130_fd_sc_hd__nand2_1 _24609_ (.A(net1430),
    .B(net1338),
    .Y(_00931_));
 sky130_fd_sc_hd__nand2_1 _24610_ (.A(net1428),
    .B(net1332),
    .Y(_00937_));
 sky130_fd_sc_hd__nand2_1 _24611_ (.A(net1427),
    .B(net1329),
    .Y(_00936_));
 sky130_fd_sc_hd__nand2_1 _24613_ (.A(net1425),
    .B(net1325),
    .Y(_00935_));
 sky130_fd_sc_hd__nand2_1 _24614_ (.A(net1310),
    .B(net1414),
    .Y(_00938_));
 sky130_fd_sc_hd__nand2_1 _24617_ (.A(net1306),
    .B(net1410),
    .Y(_00943_));
 sky130_fd_sc_hd__nand2_1 _24618_ (.A(net1206),
    .B(net1300),
    .Y(_00942_));
 sky130_fd_sc_hd__nand2_1 _24620_ (.A(net1405),
    .B(net1297),
    .Y(_00941_));
 sky130_fd_sc_hd__nor2_1 _24621_ (.A(net1165),
    .B(net1136),
    .Y(_00949_));
 sky130_fd_sc_hd__nor2_1 _24622_ (.A(net1129),
    .B(net1167),
    .Y(_00948_));
 sky130_fd_sc_hd__nand2_1 _24625_ (.A(net1273),
    .B(net1392),
    .Y(_00955_));
 sky130_fd_sc_hd__nor2_1 _24626_ (.A(net1189),
    .B(net1121),
    .Y(_00960_));
 sky130_fd_sc_hd__nor2_1 _24627_ (.A(net1700),
    .B(net1672),
    .Y(_00959_));
 sky130_fd_sc_hd__nor2_1 _24629_ (.A(net1685),
    .B(net1669),
    .Y(_00958_));
 sky130_fd_sc_hd__inv_2 _24630_ (.A(_00978_),
    .Y(_00975_));
 sky130_fd_sc_hd__nor2_1 _24631_ (.A(net1694),
    .B(_05826_),
    .Y(_03573_));
 sky130_fd_sc_hd__nand2_1 _24632_ (.A(net1363),
    .B(net1214),
    .Y(_00979_));
 sky130_fd_sc_hd__nand2_1 _24633_ (.A(net1358),
    .B(net1444),
    .Y(_00986_));
 sky130_fd_sc_hd__nand2_1 _24634_ (.A(net1352),
    .B(net1440),
    .Y(_00985_));
 sky130_fd_sc_hd__nand2_1 _24635_ (.A(net1207),
    .B(net1347),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_1 _24636_ (.A(net1133),
    .B(net1343),
    .Y(_00989_));
 sky130_fd_sc_hd__nand2_1 _24638_ (.A(net1338),
    .B(net1433),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2_1 _24639_ (.A(net1430),
    .B(net1332),
    .Y(_00987_));
 sky130_fd_sc_hd__nor2_1 _24640_ (.A(net1152),
    .B(net1714),
    .Y(_00993_));
 sky130_fd_sc_hd__nor2_1 _24641_ (.A(net1711),
    .B(net1151),
    .Y(_00992_));
 sky130_fd_sc_hd__nand2_1 _24642_ (.A(net1314),
    .B(net1422),
    .Y(_01000_));
 sky130_fd_sc_hd__nand2_1 _24643_ (.A(net1309),
    .B(net1418),
    .Y(_00999_));
 sky130_fd_sc_hd__nand2_1 _24644_ (.A(net1306),
    .B(net1413),
    .Y(_00998_));
 sky130_fd_sc_hd__nand2_1 _24645_ (.A(net1300),
    .B(net1409),
    .Y(_01003_));
 sky130_fd_sc_hd__nand2_1 _24648_ (.A(net1205),
    .B(net1297),
    .Y(_01002_));
 sky130_fd_sc_hd__nand2_1 _24650_ (.A(net1405),
    .B(net1293),
    .Y(_01001_));
 sky130_fd_sc_hd__nor2_1 _24651_ (.A(net1131),
    .B(net1164),
    .Y(_01009_));
 sky130_fd_sc_hd__nor2_1 _24652_ (.A(net1128),
    .B(net1167),
    .Y(_01008_));
 sky130_fd_sc_hd__nand2_1 _24655_ (.A(net1270),
    .B(net1392),
    .Y(_01015_));
 sky130_fd_sc_hd__nor2_1 _24656_ (.A(net1189),
    .B(net1672),
    .Y(_01020_));
 sky130_fd_sc_hd__nor2_1 _24657_ (.A(net1703),
    .B(net1669),
    .Y(_01019_));
 sky130_fd_sc_hd__inv_1 _24658_ (.A(net1453),
    .Y(_05987_));
 sky130_fd_sc_hd__nor2_1 _24661_ (.A(net1688),
    .B(net1117),
    .Y(_01018_));
 sky130_fd_sc_hd__inv_2 _24662_ (.A(_01037_),
    .Y(_01034_));
 sky130_fd_sc_hd__nand2_1 _24663_ (.A(net1154),
    .B(net1727),
    .Y(_01040_));
 sky130_fd_sc_hd__nand2_1 _24665_ (.A(net1363),
    .B(net1723),
    .Y(_01039_));
 sky130_fd_sc_hd__nand2_1 _24666_ (.A(net1358),
    .B(net1214),
    .Y(_01038_));
 sky130_fd_sc_hd__nand2_1 _24667_ (.A(net1352),
    .B(net1444),
    .Y(_01044_));
 sky130_fd_sc_hd__nand2_1 _24668_ (.A(net1347),
    .B(net1440),
    .Y(_01043_));
 sky130_fd_sc_hd__nand2_1 _24669_ (.A(net1207),
    .B(net1343),
    .Y(_01042_));
 sky130_fd_sc_hd__nand2_1 _24670_ (.A(net1132),
    .B(net1338),
    .Y(_01047_));
 sky130_fd_sc_hd__nand2_1 _24671_ (.A(net1332),
    .B(net1432),
    .Y(_01046_));
 sky130_fd_sc_hd__nand2_1 _24672_ (.A(net1429),
    .B(net1328),
    .Y(_01045_));
 sky130_fd_sc_hd__nor2_1 _24673_ (.A(net1151),
    .B(net1714),
    .Y(_01054_));
 sky130_fd_sc_hd__nor2_1 _24674_ (.A(net1711),
    .B(net1149),
    .Y(_01053_));
 sky130_fd_sc_hd__nand2_1 _24675_ (.A(net1300),
    .B(net1413),
    .Y(_01060_));
 sky130_fd_sc_hd__nand2_1 _24677_ (.A(net1406),
    .B(net1287),
    .Y(_01063_));
 sky130_fd_sc_hd__nand2_1 _24678_ (.A(_03045_),
    .B(net1284),
    .Y(_01071_));
 sky130_fd_sc_hd__nor2_1 _24679_ (.A(_20572_),
    .B(net1125),
    .Y(_01075_));
 sky130_fd_sc_hd__nor2_1 _24681_ (.A(net1202),
    .B(net1122),
    .Y(_01074_));
 sky130_fd_sc_hd__nor2_1 _24682_ (.A(net1180),
    .B(net1673),
    .Y(_01073_));
 sky130_fd_sc_hd__nor2_1 _24683_ (.A(net1189),
    .B(net1669),
    .Y(_01080_));
 sky130_fd_sc_hd__nor2_1 _24684_ (.A(net1704),
    .B(net1117),
    .Y(_01079_));
 sky130_fd_sc_hd__nor2_1 _24686_ (.A(net1689),
    .B(net1736),
    .Y(_01078_));
 sky130_fd_sc_hd__inv_2 _24687_ (.A(_01098_),
    .Y(_01095_));
 sky130_fd_sc_hd__nand2_1 _24689_ (.A(net1463),
    .B(_03082_),
    .Y(_01101_));
 sky130_fd_sc_hd__nand2_1 _24691_ (.A(net1263),
    .B(net1455),
    .Y(_01100_));
 sky130_fd_sc_hd__nand2_1 _24693_ (.A(net1154),
    .B(net1731),
    .Y(_01099_));
 sky130_fd_sc_hd__nand2_1 _24694_ (.A(net1363),
    .B(net1727),
    .Y(_01105_));
 sky130_fd_sc_hd__nand2_1 _24695_ (.A(net1358),
    .B(net1723),
    .Y(_01104_));
 sky130_fd_sc_hd__nand2_1 _24696_ (.A(net1214),
    .B(net1352),
    .Y(_01103_));
 sky130_fd_sc_hd__nand2_1 _24697_ (.A(net1347),
    .B(net1444),
    .Y(_01110_));
 sky130_fd_sc_hd__nand2_1 _24698_ (.A(net1343),
    .B(net1440),
    .Y(_01109_));
 sky130_fd_sc_hd__nand2_1 _24699_ (.A(net1207),
    .B(net1338),
    .Y(_01108_));
 sky130_fd_sc_hd__nand2_1 _24700_ (.A(net1132),
    .B(net1332),
    .Y(_01113_));
 sky130_fd_sc_hd__nand2_1 _24701_ (.A(net1328),
    .B(net1432),
    .Y(_01112_));
 sky130_fd_sc_hd__nand2_1 _24703_ (.A(net1429),
    .B(net1324),
    .Y(_01111_));
 sky130_fd_sc_hd__nor2_1 _24704_ (.A(net1149),
    .B(net1714),
    .Y(_01118_));
 sky130_fd_sc_hd__nor2_1 _24705_ (.A(net1711),
    .B(net1147),
    .Y(_01117_));
 sky130_fd_sc_hd__nand2_1 _24706_ (.A(net1306),
    .B(net1421),
    .Y(_01126_));
 sky130_fd_sc_hd__nand2_1 _24707_ (.A(net1301),
    .B(net1417),
    .Y(_01125_));
 sky130_fd_sc_hd__nand2_1 _24708_ (.A(net1297),
    .B(net1412),
    .Y(_01124_));
 sky130_fd_sc_hd__nand2_1 _24709_ (.A(net1404),
    .B(net1284),
    .Y(_01127_));
 sky130_fd_sc_hd__nor2_1 _24710_ (.A(net1400),
    .B(net1128),
    .Y(_01134_));
 sky130_fd_sc_hd__nor2_1 _24711_ (.A(net1164),
    .B(net1679),
    .Y(_01133_));
 sky130_fd_sc_hd__nor2_1 _24713_ (.A(net1168),
    .B(net1125),
    .Y(_01132_));
 sky130_fd_sc_hd__nor2_1 _24714_ (.A(_20572_),
    .B(net1121),
    .Y(_01140_));
 sky130_fd_sc_hd__nor2_1 _24715_ (.A(net1202),
    .B(net1673),
    .Y(_01139_));
 sky130_fd_sc_hd__nor2_1 _24716_ (.A(net1180),
    .B(net1671),
    .Y(_01138_));
 sky130_fd_sc_hd__nor2_1 _24717_ (.A(net1190),
    .B(net1119),
    .Y(_01145_));
 sky130_fd_sc_hd__nor2_1 _24718_ (.A(net1705),
    .B(net1738),
    .Y(_01144_));
 sky130_fd_sc_hd__inv_2 _24719_ (.A(net1467),
    .Y(_05997_));
 sky130_fd_sc_hd__nor2_1 _24721_ (.A(net1690),
    .B(net1116),
    .Y(_01143_));
 sky130_fd_sc_hd__inv_2 _24722_ (.A(_01164_),
    .Y(_01161_));
 sky130_fd_sc_hd__nor2_1 _24723_ (.A(net1694),
    .B(_19919_),
    .Y(_03606_));
 sky130_fd_sc_hd__nand2_1 _24724_ (.A(net1463),
    .B(net1263),
    .Y(_01167_));
 sky130_fd_sc_hd__nand2_1 _24726_ (.A(net1155),
    .B(net1455),
    .Y(_01166_));
 sky130_fd_sc_hd__nand2_1 _24727_ (.A(net1363),
    .B(net1731),
    .Y(_01165_));
 sky130_fd_sc_hd__nand2_1 _24728_ (.A(net1359),
    .B(net1727),
    .Y(_01171_));
 sky130_fd_sc_hd__nand2_1 _24729_ (.A(net1723),
    .B(net1353),
    .Y(_01170_));
 sky130_fd_sc_hd__nand2_1 _24730_ (.A(net1214),
    .B(net1347),
    .Y(_01169_));
 sky130_fd_sc_hd__nand2_1 _24731_ (.A(net1343),
    .B(net1444),
    .Y(_01175_));
 sky130_fd_sc_hd__nand2_1 _24732_ (.A(net1338),
    .B(net1440),
    .Y(_01174_));
 sky130_fd_sc_hd__nand2_1 _24733_ (.A(net1207),
    .B(net1332),
    .Y(_01173_));
 sky130_fd_sc_hd__nand2_1 _24735_ (.A(net1132),
    .B(net1328),
    .Y(_01178_));
 sky130_fd_sc_hd__nand2_1 _24736_ (.A(net1324),
    .B(net1432),
    .Y(_01177_));
 sky130_fd_sc_hd__nand2_1 _24738_ (.A(net1429),
    .B(net1320),
    .Y(_01176_));
 sky130_fd_sc_hd__nand2_1 _24739_ (.A(net1428),
    .B(net1314),
    .Y(_01184_));
 sky130_fd_sc_hd__nand2_1 _24740_ (.A(net1301),
    .B(net1421),
    .Y(_01189_));
 sky130_fd_sc_hd__nand2_1 _24741_ (.A(net1297),
    .B(net1417),
    .Y(_01188_));
 sky130_fd_sc_hd__nand2_1 _24742_ (.A(net1293),
    .B(net1412),
    .Y(_01187_));
 sky130_fd_sc_hd__nand2_1 _24743_ (.A(net1404),
    .B(net1279),
    .Y(_01190_));
 sky130_fd_sc_hd__nor2_1 _24744_ (.A(net1400),
    .B(net1679),
    .Y(_01196_));
 sky130_fd_sc_hd__nor2_1 _24745_ (.A(net1165),
    .B(net1125),
    .Y(_01195_));
 sky130_fd_sc_hd__nor2_1 _24746_ (.A(net1168),
    .B(net1121),
    .Y(_01194_));
 sky130_fd_sc_hd__nor2_1 _24747_ (.A(_20572_),
    .B(net1673),
    .Y(_01203_));
 sky130_fd_sc_hd__nor2_1 _24748_ (.A(net1201),
    .B(net1671),
    .Y(_01202_));
 sky130_fd_sc_hd__nor2_1 _24749_ (.A(net1180),
    .B(net1120),
    .Y(_01201_));
 sky130_fd_sc_hd__nor2_1 _24750_ (.A(net1190),
    .B(net1738),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_1 _24751_ (.A(net1705),
    .B(net1116),
    .Y(_01207_));
 sky130_fd_sc_hd__inv_2 _24752_ (.A(net1476),
    .Y(_06002_));
 sky130_fd_sc_hd__nor2_1 _24754_ (.A(net1690),
    .B(net1112),
    .Y(_01206_));
 sky130_fd_sc_hd__inv_2 _24755_ (.A(_01226_),
    .Y(_01223_));
 sky130_fd_sc_hd__nor2_1 _24756_ (.A(net1740),
    .B(net1694),
    .Y(_03617_));
 sky130_fd_sc_hd__nor2_1 _24757_ (.A(net1708),
    .B(net1220),
    .Y(_03616_));
 sky130_fd_sc_hd__nand2_1 _24759_ (.A(net1154),
    .B(net1463),
    .Y(_01229_));
 sky130_fd_sc_hd__nand2_1 _24760_ (.A(net1363),
    .B(net1455),
    .Y(_01228_));
 sky130_fd_sc_hd__nand2_1 _24761_ (.A(net1359),
    .B(net1731),
    .Y(_01227_));
 sky130_fd_sc_hd__nand2_1 _24762_ (.A(net1727),
    .B(net1352),
    .Y(_01233_));
 sky130_fd_sc_hd__nand2_1 _24763_ (.A(net1723),
    .B(net1348),
    .Y(_01232_));
 sky130_fd_sc_hd__nand2_1 _24764_ (.A(net1214),
    .B(net1343),
    .Y(_01231_));
 sky130_fd_sc_hd__nand2_1 _24765_ (.A(net1338),
    .B(net1444),
    .Y(_01238_));
 sky130_fd_sc_hd__nand2_1 _24766_ (.A(net1332),
    .B(net1440),
    .Y(_01237_));
 sky130_fd_sc_hd__nand2_1 _24767_ (.A(net1207),
    .B(net1329),
    .Y(_01236_));
 sky130_fd_sc_hd__nand2_1 _24768_ (.A(net1132),
    .B(net1325),
    .Y(_01241_));
 sky130_fd_sc_hd__nand2_1 _24769_ (.A(net1319),
    .B(net1432),
    .Y(_01240_));
 sky130_fd_sc_hd__nand2_1 _24770_ (.A(net1429),
    .B(net1314),
    .Y(_01239_));
 sky130_fd_sc_hd__nor2_1 _24771_ (.A(net1144),
    .B(net1714),
    .Y(_01244_));
 sky130_fd_sc_hd__nor2_1 _24772_ (.A(net1711),
    .B(_05935_),
    .Y(_01243_));
 sky130_fd_sc_hd__nand2_1 _24773_ (.A(net1297),
    .B(net1421),
    .Y(_01251_));
 sky130_fd_sc_hd__nand2_1 _24774_ (.A(net1293),
    .B(net1417),
    .Y(_01250_));
 sky130_fd_sc_hd__nand2_1 _24775_ (.A(net1287),
    .B(net1412),
    .Y(_01249_));
 sky130_fd_sc_hd__nand2_1 _24776_ (.A(net1259),
    .B(net1404),
    .Y(_01252_));
 sky130_fd_sc_hd__nor2_1 _24777_ (.A(net1400),
    .B(net1123),
    .Y(_01259_));
 sky130_fd_sc_hd__nor2_1 _24778_ (.A(net1165),
    .B(net1121),
    .Y(_01258_));
 sky130_fd_sc_hd__nor2_1 _24779_ (.A(net1168),
    .B(net1673),
    .Y(_01257_));
 sky130_fd_sc_hd__nor2_1 _24780_ (.A(net1171),
    .B(net1671),
    .Y(_01266_));
 sky130_fd_sc_hd__nor2_1 _24781_ (.A(net1201),
    .B(net1120),
    .Y(_01265_));
 sky130_fd_sc_hd__nor2_1 _24782_ (.A(net1180),
    .B(net1738),
    .Y(_01264_));
 sky130_fd_sc_hd__nor2_1 _24783_ (.A(net1190),
    .B(net1116),
    .Y(_01271_));
 sky130_fd_sc_hd__nor2_1 _24784_ (.A(net1705),
    .B(net1112),
    .Y(_01270_));
 sky130_fd_sc_hd__nor2_1 _24785_ (.A(net1690),
    .B(net1223),
    .Y(_01269_));
 sky130_fd_sc_hd__inv_2 _24786_ (.A(_01285_),
    .Y(_01282_));
 sky130_fd_sc_hd__nand2_1 _24787_ (.A(net1480),
    .B(\inst$top.soc.cpu.multiplier.x_src2_signed ),
    .Y(_06005_));
 sky130_fd_sc_hd__nor2_2 _24788_ (.A(net1693),
    .B(_06005_),
    .Y(_03629_));
 sky130_fd_sc_hd__nand2_1 _24791_ (.A(net1154),
    .B(net1471),
    .Y(_01288_));
 sky130_fd_sc_hd__nand2_1 _24792_ (.A(net1364),
    .B(net1462),
    .Y(_01287_));
 sky130_fd_sc_hd__nand2_1 _24793_ (.A(net1359),
    .B(net1454),
    .Y(_01286_));
 sky130_fd_sc_hd__nand2_1 _24794_ (.A(net1731),
    .B(net1352),
    .Y(_01293_));
 sky130_fd_sc_hd__nand2_1 _24795_ (.A(net1727),
    .B(net1347),
    .Y(_01292_));
 sky130_fd_sc_hd__nand2_1 _24796_ (.A(net1723),
    .B(net1342),
    .Y(_01291_));
 sky130_fd_sc_hd__nand2_1 _24797_ (.A(net1214),
    .B(net1339),
    .Y(_01297_));
 sky130_fd_sc_hd__nand2_1 _24799_ (.A(net1333),
    .B(net1444),
    .Y(_01296_));
 sky130_fd_sc_hd__nand2_1 _24800_ (.A(net1328),
    .B(net1440),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2_1 _24801_ (.A(net1207),
    .B(net1325),
    .Y(_01300_));
 sky130_fd_sc_hd__nand2_1 _24802_ (.A(net1132),
    .B(net1320),
    .Y(_01299_));
 sky130_fd_sc_hd__nand2_1 _24803_ (.A(net1314),
    .B(net1432),
    .Y(_01298_));
 sky130_fd_sc_hd__nand2_1 _24804_ (.A(net1429),
    .B(net1310),
    .Y(_01302_));
 sky130_fd_sc_hd__nand2_1 _24805_ (.A(net1425),
    .B(net1298),
    .Y(_01307_));
 sky130_fd_sc_hd__nand2_1 _24806_ (.A(net1293),
    .B(net1421),
    .Y(_01306_));
 sky130_fd_sc_hd__nand2_1 _24807_ (.A(net1287),
    .B(net1417),
    .Y(_01305_));
 sky130_fd_sc_hd__nand2_1 _24808_ (.A(net1259),
    .B(net1204),
    .Y(_01308_));
 sky130_fd_sc_hd__nor2_1 _24809_ (.A(net1709),
    .B(net1123),
    .Y(_01314_));
 sky130_fd_sc_hd__nor2_1 _24812_ (.A(net1400),
    .B(net1121),
    .Y(_01313_));
 sky130_fd_sc_hd__nor2_1 _24813_ (.A(net1164),
    .B(net1673),
    .Y(_01312_));
 sky130_fd_sc_hd__nor2_1 _24814_ (.A(net1168),
    .B(net1669),
    .Y(_01321_));
 sky130_fd_sc_hd__nor2_1 _24815_ (.A(net1171),
    .B(net1117),
    .Y(_01320_));
 sky130_fd_sc_hd__nor2_1 _24816_ (.A(net1201),
    .B(net1736),
    .Y(_01319_));
 sky130_fd_sc_hd__nor2_1 _24817_ (.A(net1180),
    .B(net1115),
    .Y(_01326_));
 sky130_fd_sc_hd__nor2_1 _24818_ (.A(net1190),
    .B(net1112),
    .Y(_01325_));
 sky130_fd_sc_hd__nor2_1 _24819_ (.A(net1705),
    .B(net1223),
    .Y(_01324_));
 sky130_fd_sc_hd__nand2_1 _24820_ (.A(net1482),
    .B(\inst$top.soc.cpu.multiplier.x_src1_signed ),
    .Y(_06011_));
 sky130_fd_sc_hd__nor2_1 _24823_ (.A(net1690),
    .B(net1108),
    .Y(_01341_));
 sky130_fd_sc_hd__inv_2 _24824_ (.A(_01350_),
    .Y(_01347_));
 sky130_fd_sc_hd__inv_2 _24825_ (.A(_06005_),
    .Y(_06014_));
 sky130_fd_sc_hd__nand2_1 _24827_ (.A(net1047),
    .B(net1708),
    .Y(_01353_));
 sky130_fd_sc_hd__nand2_1 _24829_ (.A(net1154),
    .B(net1479),
    .Y(_01352_));
 sky130_fd_sc_hd__nand2_1 _24830_ (.A(net1364),
    .B(net1471),
    .Y(_01351_));
 sky130_fd_sc_hd__a21oi_1 _24831_ (.A1(net1046),
    .A2(net1694),
    .B1(_03630_),
    .Y(_01357_));
 sky130_fd_sc_hd__nand2_1 _24832_ (.A(net1359),
    .B(net1462),
    .Y(_01356_));
 sky130_fd_sc_hd__nand2_1 _24833_ (.A(net1353),
    .B(net1454),
    .Y(_01355_));
 sky130_fd_sc_hd__nand2_1 _24834_ (.A(net1732),
    .B(net1347),
    .Y(_01354_));
 sky130_fd_sc_hd__nand2_1 _24835_ (.A(net1727),
    .B(net1342),
    .Y(_01360_));
 sky130_fd_sc_hd__nand2_1 _24836_ (.A(net1723),
    .B(net1339),
    .Y(_01359_));
 sky130_fd_sc_hd__nand2_1 _24837_ (.A(net1214),
    .B(net1333),
    .Y(_01358_));
 sky130_fd_sc_hd__nand2_1 _24838_ (.A(net1328),
    .B(net1444),
    .Y(_01363_));
 sky130_fd_sc_hd__nand2_1 _24840_ (.A(net1324),
    .B(net1440),
    .Y(_01362_));
 sky130_fd_sc_hd__nand2_1 _24841_ (.A(net1207),
    .B(net1319),
    .Y(_01361_));
 sky130_fd_sc_hd__nand2_1 _24842_ (.A(net1132),
    .B(net1315),
    .Y(_01366_));
 sky130_fd_sc_hd__nand2_1 _24843_ (.A(net1309),
    .B(net1432),
    .Y(_01365_));
 sky130_fd_sc_hd__nand2_1 _24844_ (.A(net1429),
    .B(net1306),
    .Y(_01364_));
 sky130_fd_sc_hd__nor2_1 _24845_ (.A(net1140),
    .B(net1714),
    .Y(_01368_));
 sky130_fd_sc_hd__nor2_1 _24846_ (.A(net1710),
    .B(net1138),
    .Y(_01367_));
 sky130_fd_sc_hd__nand2_1 _24847_ (.A(net1287),
    .B(net1421),
    .Y(_01375_));
 sky130_fd_sc_hd__nand2_1 _24848_ (.A(net1284),
    .B(net1417),
    .Y(_01374_));
 sky130_fd_sc_hd__nand2_1 _24849_ (.A(net1412),
    .B(net1279),
    .Y(_01373_));
 sky130_fd_sc_hd__nand2_1 _24850_ (.A(net1404),
    .B(net1271),
    .Y(_01376_));
 sky130_fd_sc_hd__nor2_1 _24851_ (.A(net1401),
    .B(net1672),
    .Y(_01382_));
 sky130_fd_sc_hd__nor2_1 _24852_ (.A(net1164),
    .B(net1669),
    .Y(_01381_));
 sky130_fd_sc_hd__nor2_1 _24853_ (.A(net1168),
    .B(net1117),
    .Y(_01380_));
 sky130_fd_sc_hd__nor2_1 _24854_ (.A(net1171),
    .B(net1736),
    .Y(_01389_));
 sky130_fd_sc_hd__nor2_1 _24855_ (.A(net1201),
    .B(net1115),
    .Y(_01388_));
 sky130_fd_sc_hd__nor2_1 _24856_ (.A(net1180),
    .B(net1112),
    .Y(_01387_));
 sky130_fd_sc_hd__nand2_1 _24858_ (.A(net1483),
    .B(net1388),
    .Y(_01393_));
 sky130_fd_sc_hd__nor2_1 _24859_ (.A(net1705),
    .B(net1108),
    .Y(_01450_));
 sky130_fd_sc_hd__nand2_1 _24860_ (.A(net1046),
    .B(net1368),
    .Y(_01412_));
 sky130_fd_sc_hd__nand2_1 _24861_ (.A(net1364),
    .B(net1479),
    .Y(_01411_));
 sky130_fd_sc_hd__nand2_1 _24862_ (.A(net1358),
    .B(net1471),
    .Y(_01410_));
 sky130_fd_sc_hd__nand2_1 _24863_ (.A(net1462),
    .B(net1352),
    .Y(_01415_));
 sky130_fd_sc_hd__nand2_1 _24864_ (.A(net1347),
    .B(net1454),
    .Y(_01414_));
 sky130_fd_sc_hd__nand2_1 _24865_ (.A(net1732),
    .B(net1342),
    .Y(_01413_));
 sky130_fd_sc_hd__nand2_1 _24866_ (.A(net1727),
    .B(net1339),
    .Y(_01418_));
 sky130_fd_sc_hd__nand2_1 _24867_ (.A(net1723),
    .B(net1333),
    .Y(_01417_));
 sky130_fd_sc_hd__nand2_1 _24868_ (.A(net1214),
    .B(net1329),
    .Y(_01416_));
 sky130_fd_sc_hd__nand2_1 _24869_ (.A(net1324),
    .B(net1444),
    .Y(_01421_));
 sky130_fd_sc_hd__nand2_1 _24870_ (.A(net1319),
    .B(net1440),
    .Y(_01420_));
 sky130_fd_sc_hd__nand2_1 _24871_ (.A(net1207),
    .B(net1315),
    .Y(_01419_));
 sky130_fd_sc_hd__nand2_1 _24872_ (.A(net1132),
    .B(net1309),
    .Y(_01424_));
 sky130_fd_sc_hd__nand2_1 _24873_ (.A(net1305),
    .B(net1432),
    .Y(_01423_));
 sky130_fd_sc_hd__nand2_1 _24874_ (.A(net1429),
    .B(net1301),
    .Y(_01422_));
 sky130_fd_sc_hd__nand2_1 _24875_ (.A(net1425),
    .B(net1291),
    .Y(_01425_));
 sky130_fd_sc_hd__nand2_1 _24876_ (.A(net1284),
    .B(net1422),
    .Y(_01432_));
 sky130_fd_sc_hd__nand2_1 _24877_ (.A(net1418),
    .B(net1279),
    .Y(_01431_));
 sky130_fd_sc_hd__nand2_1 _24878_ (.A(net1259),
    .B(net1413),
    .Y(_01430_));
 sky130_fd_sc_hd__inv_2 _24879_ (.A(net1674),
    .Y(_06018_));
 sky130_fd_sc_hd__nand2_1 _24881_ (.A(net1257),
    .B(net1404),
    .Y(_01433_));
 sky130_fd_sc_hd__nor2_1 _24882_ (.A(net1401),
    .B(net1669),
    .Y(_01439_));
 sky130_fd_sc_hd__nor2_1 _24883_ (.A(net1164),
    .B(net1117),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_1 _24884_ (.A(net1168),
    .B(net1736),
    .Y(_01437_));
 sky130_fd_sc_hd__nor2_1 _24885_ (.A(net1171),
    .B(net1115),
    .Y(_01446_));
 sky130_fd_sc_hd__nor2_1 _24886_ (.A(net1201),
    .B(net1111),
    .Y(_01445_));
 sky130_fd_sc_hd__nor2_1 _24887_ (.A(net1180),
    .B(net1223),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_1 _24889_ (.A(net1190),
    .B(net1109),
    .Y(_01449_));
 sky130_fd_sc_hd__inv_2 _24890_ (.A(_01468_),
    .Y(_01465_));
 sky130_fd_sc_hd__nand2_1 _24891_ (.A(net1046),
    .B(_05900_),
    .Y(_01471_));
 sky130_fd_sc_hd__nand2_1 _24892_ (.A(net1358),
    .B(net1479),
    .Y(_01470_));
 sky130_fd_sc_hd__nand2_1 _24894_ (.A(net1472),
    .B(net1352),
    .Y(_01469_));
 sky130_fd_sc_hd__nand2_1 _24895_ (.A(net1462),
    .B(net1347),
    .Y(_01474_));
 sky130_fd_sc_hd__nand2_1 _24896_ (.A(net1342),
    .B(net1454),
    .Y(_01473_));
 sky130_fd_sc_hd__nand2_1 _24897_ (.A(net1731),
    .B(net1338),
    .Y(_01472_));
 sky130_fd_sc_hd__nand2_1 _24898_ (.A(net1727),
    .B(net1333),
    .Y(_01477_));
 sky130_fd_sc_hd__nand2_1 _24899_ (.A(net1723),
    .B(net1328),
    .Y(_01476_));
 sky130_fd_sc_hd__nand2_1 _24900_ (.A(net1214),
    .B(net1324),
    .Y(_01475_));
 sky130_fd_sc_hd__nand2_1 _24901_ (.A(net1319),
    .B(net1445),
    .Y(_01480_));
 sky130_fd_sc_hd__nand2_1 _24902_ (.A(net1314),
    .B(net1441),
    .Y(_01479_));
 sky130_fd_sc_hd__nand2_1 _24904_ (.A(net1208),
    .B(net1309),
    .Y(_01478_));
 sky130_fd_sc_hd__nand2_1 _24905_ (.A(net1135),
    .B(net1306),
    .Y(_01483_));
 sky130_fd_sc_hd__nand2_1 _24906_ (.A(net1301),
    .B(net1436),
    .Y(_01482_));
 sky130_fd_sc_hd__nand2_1 _24907_ (.A(_20014_),
    .B(net1298),
    .Y(_01481_));
 sky130_fd_sc_hd__nor2_1 _24909_ (.A(net1715),
    .B(_05945_),
    .Y(_01485_));
 sky130_fd_sc_hd__nor2_1 _24911_ (.A(net1711),
    .B(net1131),
    .Y(_01484_));
 sky130_fd_sc_hd__nand2_1 _24912_ (.A(net1421),
    .B(net1279),
    .Y(_01492_));
 sky130_fd_sc_hd__nand2_1 _24913_ (.A(net1259),
    .B(net1418),
    .Y(_01491_));
 sky130_fd_sc_hd__nand2_1 _24914_ (.A(net1274),
    .B(net1413),
    .Y(_01490_));
 sky130_fd_sc_hd__inv_1 _24915_ (.A(net1670),
    .Y(_06023_));
 sky130_fd_sc_hd__nand2_1 _24918_ (.A(net1254),
    .B(net1404),
    .Y(_01493_));
 sky130_fd_sc_hd__nor2_1 _24919_ (.A(net1400),
    .B(net1117),
    .Y(_01499_));
 sky130_fd_sc_hd__nor2_1 _24920_ (.A(net1164),
    .B(net1736),
    .Y(_01498_));
 sky130_fd_sc_hd__nor2_1 _24921_ (.A(net1168),
    .B(net1115),
    .Y(_01497_));
 sky130_fd_sc_hd__nor2_1 _24922_ (.A(net1171),
    .B(net1111),
    .Y(_01506_));
 sky130_fd_sc_hd__nor2_1 _24923_ (.A(net1201),
    .B(net1221),
    .Y(_01505_));
 sky130_fd_sc_hd__nor2_1 _24924_ (.A(net1180),
    .B(net1108),
    .Y(_01504_));
 sky130_fd_sc_hd__inv_2 _24925_ (.A(_01524_),
    .Y(_01521_));
 sky130_fd_sc_hd__nand2_1 _24926_ (.A(net1045),
    .B(_05894_),
    .Y(_01527_));
 sky130_fd_sc_hd__nand2_1 _24927_ (.A(net1478),
    .B(net1352),
    .Y(_01526_));
 sky130_fd_sc_hd__nand2_1 _24928_ (.A(net1471),
    .B(net1347),
    .Y(_01525_));
 sky130_fd_sc_hd__nand2_1 _24929_ (.A(net1462),
    .B(net1342),
    .Y(_01530_));
 sky130_fd_sc_hd__nand2_1 _24930_ (.A(net1339),
    .B(net1454),
    .Y(_01529_));
 sky130_fd_sc_hd__nand2_1 _24931_ (.A(net1731),
    .B(net1333),
    .Y(_01528_));
 sky130_fd_sc_hd__nand2_1 _24932_ (.A(net1727),
    .B(net1328),
    .Y(_01533_));
 sky130_fd_sc_hd__nand2_1 _24933_ (.A(net1723),
    .B(net1324),
    .Y(_01532_));
 sky130_fd_sc_hd__nand2_1 _24934_ (.A(net1215),
    .B(net1319),
    .Y(_01531_));
 sky130_fd_sc_hd__nand2_1 _24935_ (.A(net1314),
    .B(net1445),
    .Y(_01536_));
 sky130_fd_sc_hd__nand2_1 _24936_ (.A(net1309),
    .B(net1441),
    .Y(_01535_));
 sky130_fd_sc_hd__nand2_1 _24937_ (.A(net1208),
    .B(net1306),
    .Y(_01534_));
 sky130_fd_sc_hd__nor2_1 _24938_ (.A(net1131),
    .B(net1714),
    .Y(_01544_));
 sky130_fd_sc_hd__nor2_1 _24939_ (.A(net1711),
    .B(net1128),
    .Y(_01543_));
 sky130_fd_sc_hd__nand2_1 _24940_ (.A(net1259),
    .B(net1422),
    .Y(_01552_));
 sky130_fd_sc_hd__nand2_1 _24941_ (.A(net1274),
    .B(net1418),
    .Y(_01551_));
 sky130_fd_sc_hd__nand2_1 _24942_ (.A(net1271),
    .B(net1412),
    .Y(_01550_));
 sky130_fd_sc_hd__nand2_1 _24943_ (.A(net1405),
    .B(_19952_),
    .Y(_01553_));
 sky130_fd_sc_hd__nor2_1 _24944_ (.A(net1400),
    .B(net1736),
    .Y(_01559_));
 sky130_fd_sc_hd__nor2_1 _24945_ (.A(net1164),
    .B(net1115),
    .Y(_01558_));
 sky130_fd_sc_hd__nor2_1 _24946_ (.A(net1167),
    .B(net1111),
    .Y(_01557_));
 sky130_fd_sc_hd__nor2_1 _24947_ (.A(net1201),
    .B(net1108),
    .Y(_01564_));
 sky130_fd_sc_hd__inv_2 _24948_ (.A(_01564_),
    .Y(_01621_));
 sky130_fd_sc_hd__inv_2 _24949_ (.A(_01582_),
    .Y(_01579_));
 sky130_fd_sc_hd__nand2_1 _24950_ (.A(net1045),
    .B(_05896_),
    .Y(_01585_));
 sky130_fd_sc_hd__nand2_1 _24951_ (.A(net1478),
    .B(net1347),
    .Y(_01584_));
 sky130_fd_sc_hd__nand2_1 _24952_ (.A(net1471),
    .B(net1342),
    .Y(_01583_));
 sky130_fd_sc_hd__nand2_1 _24953_ (.A(net1462),
    .B(net1338),
    .Y(_01588_));
 sky130_fd_sc_hd__nand2_1 _24955_ (.A(net1333),
    .B(net1455),
    .Y(_01587_));
 sky130_fd_sc_hd__nand2_1 _24956_ (.A(net1731),
    .B(net1328),
    .Y(_01586_));
 sky130_fd_sc_hd__nand2_1 _24957_ (.A(net1728),
    .B(net1324),
    .Y(_01591_));
 sky130_fd_sc_hd__nand2_1 _24958_ (.A(net1724),
    .B(net1319),
    .Y(_01590_));
 sky130_fd_sc_hd__nand2_1 _24959_ (.A(net1215),
    .B(net1314),
    .Y(_01589_));
 sky130_fd_sc_hd__nand2_1 _24960_ (.A(net1309),
    .B(net1445),
    .Y(_01594_));
 sky130_fd_sc_hd__nand2_1 _24961_ (.A(net1305),
    .B(net1441),
    .Y(_01593_));
 sky130_fd_sc_hd__nand2_1 _24962_ (.A(net1208),
    .B(net1301),
    .Y(_01592_));
 sky130_fd_sc_hd__nand2_1 _24963_ (.A(net1135),
    .B(net1298),
    .Y(_01597_));
 sky130_fd_sc_hd__nand2_1 _24964_ (.A(net1293),
    .B(net1432),
    .Y(_01596_));
 sky130_fd_sc_hd__nand2_1 _24965_ (.A(net1429),
    .B(net1291),
    .Y(_01595_));
 sky130_fd_sc_hd__nor2_1 _24966_ (.A(net1128),
    .B(net1715),
    .Y(_01599_));
 sky130_fd_sc_hd__nor2_1 _24967_ (.A(net1710),
    .B(net1679),
    .Y(_01598_));
 sky130_fd_sc_hd__nand2_1 _24968_ (.A(net1274),
    .B(net1422),
    .Y(_01608_));
 sky130_fd_sc_hd__nand2_1 _24969_ (.A(net1270),
    .B(net1417),
    .Y(_01607_));
 sky130_fd_sc_hd__nand2_1 _24970_ (.A(net1257),
    .B(net1412),
    .Y(_01606_));
 sky130_fd_sc_hd__nand2_1 _24971_ (.A(net1461),
    .B(net1404),
    .Y(_01609_));
 sky130_fd_sc_hd__nor2_1 _24972_ (.A(net1400),
    .B(net1115),
    .Y(_01615_));
 sky130_fd_sc_hd__nor2_1 _24973_ (.A(net1164),
    .B(net1111),
    .Y(_01614_));
 sky130_fd_sc_hd__nor2_1 _24974_ (.A(net1167),
    .B(net1221),
    .Y(_01613_));
 sky130_fd_sc_hd__inv_2 _24975_ (.A(_01636_),
    .Y(_01633_));
 sky130_fd_sc_hd__nand2_1 _24976_ (.A(net1045),
    .B(net1159),
    .Y(_01639_));
 sky130_fd_sc_hd__nand2_1 _24977_ (.A(net1478),
    .B(net1342),
    .Y(_01638_));
 sky130_fd_sc_hd__nand2_1 _24978_ (.A(net1471),
    .B(net1338),
    .Y(_01637_));
 sky130_fd_sc_hd__nand2_1 _24979_ (.A(net1463),
    .B(net1332),
    .Y(_01642_));
 sky130_fd_sc_hd__nand2_1 _24980_ (.A(net1328),
    .B(net1454),
    .Y(_01641_));
 sky130_fd_sc_hd__nand2_1 _24981_ (.A(net1731),
    .B(net1324),
    .Y(_01640_));
 sky130_fd_sc_hd__nand2_1 _24982_ (.A(net1728),
    .B(net1319),
    .Y(_01645_));
 sky130_fd_sc_hd__nand2_1 _24983_ (.A(net1724),
    .B(net1314),
    .Y(_01644_));
 sky130_fd_sc_hd__nand2_1 _24984_ (.A(net1215),
    .B(net1309),
    .Y(_01643_));
 sky130_fd_sc_hd__nand2_1 _24985_ (.A(net1305),
    .B(net1445),
    .Y(_01648_));
 sky130_fd_sc_hd__nand2_1 _24986_ (.A(net1300),
    .B(net1441),
    .Y(_01647_));
 sky130_fd_sc_hd__nand2_1 _24987_ (.A(net1208),
    .B(net1297),
    .Y(_01646_));
 sky130_fd_sc_hd__nand2_1 _24988_ (.A(net1429),
    .B(net1284),
    .Y(_01649_));
 sky130_fd_sc_hd__nor2_1 _24989_ (.A(net1715),
    .B(net1677),
    .Y(_01653_));
 sky130_fd_sc_hd__nor2_1 _24990_ (.A(net1710),
    .B(net1123),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_1 _24991_ (.A(net1270),
    .B(net1421),
    .Y(_01661_));
 sky130_fd_sc_hd__nand2_1 _24992_ (.A(net1255),
    .B(net1417),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2_1 _24993_ (.A(net1254),
    .B(net1412),
    .Y(_01659_));
 sky130_fd_sc_hd__nand2_1 _24994_ (.A(net1470),
    .B(net1404),
    .Y(_01662_));
 sky130_fd_sc_hd__nor2_1 _24995_ (.A(net1400),
    .B(net1111),
    .Y(_01668_));
 sky130_fd_sc_hd__nor2_1 _24996_ (.A(net1164),
    .B(net1221),
    .Y(_01667_));
 sky130_fd_sc_hd__nor2_1 _24997_ (.A(net1167),
    .B(net1108),
    .Y(_01666_));
 sky130_fd_sc_hd__inv_2 _24998_ (.A(_01688_),
    .Y(_01685_));
 sky130_fd_sc_hd__nand2_1 _24999_ (.A(net1046),
    .B(_05901_),
    .Y(_01691_));
 sky130_fd_sc_hd__nand2_1 _25000_ (.A(net1478),
    .B(net1338),
    .Y(_01690_));
 sky130_fd_sc_hd__nand2_1 _25001_ (.A(net1471),
    .B(net1332),
    .Y(_01689_));
 sky130_fd_sc_hd__nand2_1 _25002_ (.A(net1462),
    .B(net1328),
    .Y(_01694_));
 sky130_fd_sc_hd__nand2_1 _25003_ (.A(net1324),
    .B(net1454),
    .Y(_01693_));
 sky130_fd_sc_hd__nand2_1 _25004_ (.A(net1731),
    .B(net1319),
    .Y(_01692_));
 sky130_fd_sc_hd__nand2_1 _25005_ (.A(net1728),
    .B(net1314),
    .Y(_01697_));
 sky130_fd_sc_hd__nand2_1 _25006_ (.A(net1724),
    .B(net1309),
    .Y(_01696_));
 sky130_fd_sc_hd__nand2_1 _25007_ (.A(net1215),
    .B(net1305),
    .Y(_01695_));
 sky130_fd_sc_hd__nand2_1 _25008_ (.A(net1300),
    .B(net1445),
    .Y(_01700_));
 sky130_fd_sc_hd__nand2_1 _25009_ (.A(net1297),
    .B(net1441),
    .Y(_01699_));
 sky130_fd_sc_hd__nand2_1 _25010_ (.A(net1208),
    .B(net1294),
    .Y(_01698_));
 sky130_fd_sc_hd__nand2_1 _25011_ (.A(net1132),
    .B(net1290),
    .Y(_01703_));
 sky130_fd_sc_hd__nand2_1 _25012_ (.A(net1432),
    .B(net1284),
    .Y(_01702_));
 sky130_fd_sc_hd__nand2_1 _25013_ (.A(net1429),
    .B(net1278),
    .Y(_01701_));
 sky130_fd_sc_hd__nor2_1 _25014_ (.A(net1715),
    .B(net1123),
    .Y(_01705_));
 sky130_fd_sc_hd__nor2_1 _25015_ (.A(net1710),
    .B(net1121),
    .Y(_01704_));
 sky130_fd_sc_hd__nand2_1 _25016_ (.A(net1255),
    .B(net1421),
    .Y(_01713_));
 sky130_fd_sc_hd__nand2_1 _25017_ (.A(net1254),
    .B(net1417),
    .Y(_01712_));
 sky130_fd_sc_hd__nand2_1 _25018_ (.A(_19952_),
    .B(net1412),
    .Y(_01711_));
 sky130_fd_sc_hd__nand2_1 _25019_ (.A(net1404),
    .B(net1477),
    .Y(_01714_));
 sky130_fd_sc_hd__nand2_1 _25020_ (.A(net1481),
    .B(_03045_),
    .Y(_01719_));
 sky130_fd_sc_hd__nor2_1 _25021_ (.A(net1164),
    .B(net1108),
    .Y(_01769_));
 sky130_fd_sc_hd__inv_2 _25022_ (.A(_01738_),
    .Y(_01735_));
 sky130_fd_sc_hd__nand2_1 _25023_ (.A(net1046),
    .B(_05903_),
    .Y(_01741_));
 sky130_fd_sc_hd__nand2_1 _25024_ (.A(net1478),
    .B(net1332),
    .Y(_01740_));
 sky130_fd_sc_hd__nand2_1 _25025_ (.A(net1471),
    .B(net1329),
    .Y(_01739_));
 sky130_fd_sc_hd__nand2_1 _25026_ (.A(net1462),
    .B(net1324),
    .Y(_01744_));
 sky130_fd_sc_hd__nand2_1 _25027_ (.A(net1319),
    .B(net1454),
    .Y(_01743_));
 sky130_fd_sc_hd__nand2_1 _25028_ (.A(net1731),
    .B(net1314),
    .Y(_01742_));
 sky130_fd_sc_hd__nand2_1 _25029_ (.A(net1728),
    .B(net1309),
    .Y(_01747_));
 sky130_fd_sc_hd__nand2_1 _25030_ (.A(net1724),
    .B(net1305),
    .Y(_01746_));
 sky130_fd_sc_hd__nand2_1 _25031_ (.A(net1215),
    .B(net1301),
    .Y(_01745_));
 sky130_fd_sc_hd__nand2_1 _25032_ (.A(net1297),
    .B(net1445),
    .Y(_01750_));
 sky130_fd_sc_hd__nand2_1 _25033_ (.A(net1293),
    .B(net1441),
    .Y(_01749_));
 sky130_fd_sc_hd__nand2_1 _25034_ (.A(net1208),
    .B(net1287),
    .Y(_01748_));
 sky130_fd_sc_hd__nand2_1 _25036_ (.A(net1259),
    .B(_20014_),
    .Y(_01751_));
 sky130_fd_sc_hd__nor2_1 _25037_ (.A(net1121),
    .B(net1714),
    .Y(_01755_));
 sky130_fd_sc_hd__nor2_1 _25038_ (.A(net1710),
    .B(net1672),
    .Y(_01754_));
 sky130_fd_sc_hd__nand2_1 _25039_ (.A(net1252),
    .B(net1421),
    .Y(_01763_));
 sky130_fd_sc_hd__nand2_1 _25040_ (.A(_19952_),
    .B(net1417),
    .Y(_01762_));
 sky130_fd_sc_hd__nand2_1 _25041_ (.A(net1461),
    .B(net1412),
    .Y(_01761_));
 sky130_fd_sc_hd__nand2_1 _25042_ (.A(net1481),
    .B(net1404),
    .Y(_01764_));
 sky130_fd_sc_hd__nor2_1 _25043_ (.A(net1400),
    .B(net1109),
    .Y(_01768_));
 sky130_fd_sc_hd__inv_2 _25044_ (.A(_01787_),
    .Y(_01784_));
 sky130_fd_sc_hd__nand2_1 _25045_ (.A(net1046),
    .B(_05907_),
    .Y(_01790_));
 sky130_fd_sc_hd__nand2_1 _25046_ (.A(net1478),
    .B(net1329),
    .Y(_01789_));
 sky130_fd_sc_hd__nand2_1 _25047_ (.A(net1471),
    .B(net1325),
    .Y(_01788_));
 sky130_fd_sc_hd__nand2_1 _25048_ (.A(net1462),
    .B(net1319),
    .Y(_01793_));
 sky130_fd_sc_hd__nand2_1 _25049_ (.A(net1315),
    .B(net1454),
    .Y(_01792_));
 sky130_fd_sc_hd__nand2_1 _25050_ (.A(net1732),
    .B(net1310),
    .Y(_01791_));
 sky130_fd_sc_hd__nand2_1 _25051_ (.A(net1728),
    .B(net1305),
    .Y(_01796_));
 sky130_fd_sc_hd__nand2_1 _25052_ (.A(net1724),
    .B(net1300),
    .Y(_01795_));
 sky130_fd_sc_hd__nand2_1 _25053_ (.A(net1214),
    .B(net1297),
    .Y(_01794_));
 sky130_fd_sc_hd__nand2_1 _25054_ (.A(net1293),
    .B(net1444),
    .Y(_01799_));
 sky130_fd_sc_hd__nand2_1 _25055_ (.A(net1287),
    .B(net1440),
    .Y(_01798_));
 sky130_fd_sc_hd__nand2_1 _25056_ (.A(net1207),
    .B(net1284),
    .Y(_01797_));
 sky130_fd_sc_hd__nand2_1 _25057_ (.A(net1132),
    .B(net1278),
    .Y(_01802_));
 sky130_fd_sc_hd__nand2_1 _25059_ (.A(net1259),
    .B(net1436),
    .Y(_01801_));
 sky130_fd_sc_hd__nand2_1 _25060_ (.A(net1430),
    .B(net1274),
    .Y(_01800_));
 sky130_fd_sc_hd__nor2_1 _25061_ (.A(net1714),
    .B(net1672),
    .Y(_01804_));
 sky130_fd_sc_hd__nor2_1 _25062_ (.A(net1710),
    .B(net1669),
    .Y(_01803_));
 sky130_fd_sc_hd__nand2_1 _25063_ (.A(net1452),
    .B(net1421),
    .Y(_01812_));
 sky130_fd_sc_hd__nand2_1 _25064_ (.A(net1459),
    .B(net1417),
    .Y(_01811_));
 sky130_fd_sc_hd__nand2_1 _25065_ (.A(net1466),
    .B(net1413),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_1 _25067_ (.A(net1323),
    .B(net1112),
    .Y(_01815_));
 sky130_fd_sc_hd__nor2_1 _25068_ (.A(net1407),
    .B(net1221),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_1 _25069_ (.A(net1709),
    .B(net1108),
    .Y(_01813_));
 sky130_fd_sc_hd__inv_2 _25070_ (.A(_01835_),
    .Y(_01832_));
 sky130_fd_sc_hd__nand2_1 _25071_ (.A(net1046),
    .B(_05908_),
    .Y(_01838_));
 sky130_fd_sc_hd__nand2_1 _25072_ (.A(net1478),
    .B(net1325),
    .Y(_01837_));
 sky130_fd_sc_hd__nand2_1 _25073_ (.A(net1471),
    .B(net1320),
    .Y(_01836_));
 sky130_fd_sc_hd__nand2_1 _25074_ (.A(net1462),
    .B(net1315),
    .Y(_01841_));
 sky130_fd_sc_hd__nand2_1 _25075_ (.A(net1310),
    .B(net1454),
    .Y(_01840_));
 sky130_fd_sc_hd__nand2_1 _25076_ (.A(net1732),
    .B(net1305),
    .Y(_01839_));
 sky130_fd_sc_hd__nor2_1 _25077_ (.A(net1140),
    .B(net1267),
    .Y(_01843_));
 sky130_fd_sc_hd__nor2_1 _25078_ (.A(net1449),
    .B(net1138),
    .Y(_01842_));
 sky130_fd_sc_hd__nand2_1 _25079_ (.A(net1258),
    .B(net1133),
    .Y(_01855_));
 sky130_fd_sc_hd__nand2_1 _25080_ (.A(net1274),
    .B(net1433),
    .Y(_01854_));
 sky130_fd_sc_hd__nand2_1 _25081_ (.A(net1430),
    .B(net1270),
    .Y(_01853_));
 sky130_fd_sc_hd__nor2_1 _25082_ (.A(net1669),
    .B(net1714),
    .Y(_01858_));
 sky130_fd_sc_hd__nor2_1 _25083_ (.A(net1710),
    .B(net1117),
    .Y(_01857_));
 sky130_fd_sc_hd__nand2_1 _25084_ (.A(net1459),
    .B(net1422),
    .Y(_01866_));
 sky130_fd_sc_hd__nand2_1 _25085_ (.A(net1466),
    .B(net1418),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _25086_ (.A(net1477),
    .B(net1413),
    .Y(_01864_));
 sky130_fd_sc_hd__inv_2 _25087_ (.A(_01888_),
    .Y(_01885_));
 sky130_fd_sc_hd__nand2_1 _25089_ (.A(net1047),
    .B(_05912_),
    .Y(_01891_));
 sky130_fd_sc_hd__nand2_1 _25090_ (.A(net1478),
    .B(net1320),
    .Y(_01890_));
 sky130_fd_sc_hd__nand2_1 _25091_ (.A(net1472),
    .B(net1315),
    .Y(_01889_));
 sky130_fd_sc_hd__nand2_1 _25092_ (.A(net1463),
    .B(net1310),
    .Y(_01894_));
 sky130_fd_sc_hd__nand2_1 _25093_ (.A(net1305),
    .B(net1456),
    .Y(_01893_));
 sky130_fd_sc_hd__nand2_1 _25094_ (.A(net1732),
    .B(net1300),
    .Y(_01892_));
 sky130_fd_sc_hd__nor2_1 _25095_ (.A(net1267),
    .B(net1138),
    .Y(_01896_));
 sky130_fd_sc_hd__nor2_1 _25096_ (.A(net1449),
    .B(_05945_),
    .Y(_01895_));
 sky130_fd_sc_hd__nor2_1 _25097_ (.A(net1126),
    .B(net1211),
    .Y(_01903_));
 sky130_fd_sc_hd__nor2_1 _25098_ (.A(net1438),
    .B(net1677),
    .Y(_01902_));
 sky130_fd_sc_hd__nand2_1 _25099_ (.A(net1255),
    .B(net1430),
    .Y(_01907_));
 sky130_fd_sc_hd__nand2_1 _25100_ (.A(net1428),
    .B(net1252),
    .Y(_01914_));
 sky130_fd_sc_hd__nor2_1 _25101_ (.A(_03017_),
    .B(net1111),
    .Y(_01917_));
 sky130_fd_sc_hd__nor2_1 _25102_ (.A(net1318),
    .B(net1221),
    .Y(_01916_));
 sky130_fd_sc_hd__inv_2 _25103_ (.A(_01941_),
    .Y(_01938_));
 sky130_fd_sc_hd__nand2_1 _25104_ (.A(net1047),
    .B(net1151),
    .Y(_01944_));
 sky130_fd_sc_hd__nand2_1 _25105_ (.A(net1478),
    .B(net1315),
    .Y(_01943_));
 sky130_fd_sc_hd__nand2_1 _25106_ (.A(net1474),
    .B(net1310),
    .Y(_01942_));
 sky130_fd_sc_hd__nand2_1 _25107_ (.A(net1463),
    .B(net1305),
    .Y(_01947_));
 sky130_fd_sc_hd__nand2_1 _25108_ (.A(net1300),
    .B(net1456),
    .Y(_01946_));
 sky130_fd_sc_hd__nand2_1 _25109_ (.A(net1732),
    .B(net1298),
    .Y(_01945_));
 sky130_fd_sc_hd__nor2_1 _25110_ (.A(net1267),
    .B(_05945_),
    .Y(_01949_));
 sky130_fd_sc_hd__nor2_1 _25111_ (.A(net1129),
    .B(net1449),
    .Y(_01948_));
 sky130_fd_sc_hd__nand2_1 _25112_ (.A(net1209),
    .B(net1273),
    .Y(_01955_));
 sky130_fd_sc_hd__nand2_1 _25113_ (.A(net1431),
    .B(net1252),
    .Y(_01959_));
 sky130_fd_sc_hd__nor2_1 _25115_ (.A(net1718),
    .B(net1117),
    .Y(_01965_));
 sky130_fd_sc_hd__nor2_1 _25117_ (.A(net1736),
    .B(net1714),
    .Y(_01964_));
 sky130_fd_sc_hd__nor2_1 _25118_ (.A(net1710),
    .B(net1115),
    .Y(_01963_));
 sky130_fd_sc_hd__nor2_1 _25119_ (.A(_03011_),
    .B(net1111),
    .Y(_01971_));
 sky130_fd_sc_hd__nor2_1 _25120_ (.A(_03017_),
    .B(net1221),
    .Y(_01970_));
 sky130_fd_sc_hd__nor2_1 _25121_ (.A(net1318),
    .B(net1108),
    .Y(_01969_));
 sky130_fd_sc_hd__inv_2 _25122_ (.A(_01989_),
    .Y(_01986_));
 sky130_fd_sc_hd__nand2_1 _25123_ (.A(net1046),
    .B(net1149),
    .Y(_01992_));
 sky130_fd_sc_hd__nand2_1 _25124_ (.A(net1478),
    .B(net1311),
    .Y(_01991_));
 sky130_fd_sc_hd__nand2_1 _25125_ (.A(net1472),
    .B(net1307),
    .Y(_01990_));
 sky130_fd_sc_hd__nand2_1 _25126_ (.A(net1464),
    .B(net1302),
    .Y(_01995_));
 sky130_fd_sc_hd__nand2_1 _25127_ (.A(net1296),
    .B(net1456),
    .Y(_01994_));
 sky130_fd_sc_hd__nand2_1 _25128_ (.A(net1292),
    .B(net1733),
    .Y(_01993_));
 sky130_fd_sc_hd__nor2_1 _25129_ (.A(net1129),
    .B(net1267),
    .Y(_01997_));
 sky130_fd_sc_hd__nor2_1 _25130_ (.A(net1126),
    .B(net1449),
    .Y(_01996_));
 sky130_fd_sc_hd__nand2_1 _25131_ (.A(net1209),
    .B(net1271),
    .Y(_02003_));
 sky130_fd_sc_hd__nand2_1 _25132_ (.A(net1431),
    .B(net1452),
    .Y(_02006_));
 sky130_fd_sc_hd__nor2_1 _25133_ (.A(net1736),
    .B(net1718),
    .Y(_02011_));
 sky130_fd_sc_hd__nor2_1 _25135_ (.A(net1715),
    .B(net1115),
    .Y(_02010_));
 sky130_fd_sc_hd__nor2_1 _25136_ (.A(net1710),
    .B(net1111),
    .Y(_02009_));
 sky130_fd_sc_hd__nand2_1 _25137_ (.A(net1481),
    .B(net1423),
    .Y(_02017_));
 sky130_fd_sc_hd__inv_1 _25138_ (.A(net1106),
    .Y(_06033_));
 sky130_fd_sc_hd__nand2_1 _25139_ (.A(_06033_),
    .B(net1419),
    .Y(_02016_));
 sky130_fd_sc_hd__inv_2 _25140_ (.A(_02036_),
    .Y(_02033_));
 sky130_fd_sc_hd__nand2_1 _25141_ (.A(net1046),
    .B(net1147),
    .Y(_02039_));
 sky130_fd_sc_hd__nand2_1 _25142_ (.A(net1479),
    .B(net1307),
    .Y(_02038_));
 sky130_fd_sc_hd__nand2_1 _25143_ (.A(net1472),
    .B(net1302),
    .Y(_02037_));
 sky130_fd_sc_hd__nand2_1 _25144_ (.A(net1464),
    .B(net1296),
    .Y(_02042_));
 sky130_fd_sc_hd__nand2_1 _25145_ (.A(net1292),
    .B(net1456),
    .Y(_02041_));
 sky130_fd_sc_hd__nand2_1 _25146_ (.A(net1288),
    .B(net1733),
    .Y(_02040_));
 sky130_fd_sc_hd__nor2_1 _25147_ (.A(net1126),
    .B(net1267),
    .Y(_02044_));
 sky130_fd_sc_hd__nor2_1 _25148_ (.A(net1449),
    .B(net1677),
    .Y(_02043_));
 sky130_fd_sc_hd__nand2_1 _25149_ (.A(net1255),
    .B(net1209),
    .Y(_02050_));
 sky130_fd_sc_hd__nand2_1 _25150_ (.A(net1431),
    .B(net1459),
    .Y(_02054_));
 sky130_fd_sc_hd__nor2_1 _25151_ (.A(net1721),
    .B(net1115),
    .Y(_02059_));
 sky130_fd_sc_hd__nor2_1 _25152_ (.A(net1715),
    .B(net1111),
    .Y(_02058_));
 sky130_fd_sc_hd__nor2_1 _25154_ (.A(net1712),
    .B(net1221),
    .Y(_02057_));
 sky130_fd_sc_hd__nand2_1 _25155_ (.A(_06033_),
    .B(net1423),
    .Y(_02064_));
 sky130_fd_sc_hd__inv_2 _25156_ (.A(_02082_),
    .Y(_02079_));
 sky130_fd_sc_hd__nand2_1 _25157_ (.A(net1046),
    .B(net1144),
    .Y(_02085_));
 sky130_fd_sc_hd__nand2_1 _25158_ (.A(net1479),
    .B(net1302),
    .Y(_02084_));
 sky130_fd_sc_hd__nand2_1 _25159_ (.A(net1472),
    .B(net1296),
    .Y(_02083_));
 sky130_fd_sc_hd__nand2_1 _25160_ (.A(net1292),
    .B(net1464),
    .Y(_02088_));
 sky130_fd_sc_hd__nand2_1 _25161_ (.A(net1288),
    .B(net1456),
    .Y(_02087_));
 sky130_fd_sc_hd__nand2_1 _25162_ (.A(net1733),
    .B(net1283),
    .Y(_02086_));
 sky130_fd_sc_hd__nor2_1 _25163_ (.A(net1267),
    .B(net1677),
    .Y(_02090_));
 sky130_fd_sc_hd__nor2_1 _25164_ (.A(net1449),
    .B(net1123),
    .Y(_02089_));
 sky130_fd_sc_hd__nand2_1 _25165_ (.A(net1252),
    .B(net1209),
    .Y(_02096_));
 sky130_fd_sc_hd__nand2_1 _25166_ (.A(net1466),
    .B(net1431),
    .Y(_02099_));
 sky130_fd_sc_hd__nor2_1 _25167_ (.A(net1721),
    .B(net1111),
    .Y(_02104_));
 sky130_fd_sc_hd__nor2_1 _25168_ (.A(net1715),
    .B(net1221),
    .Y(_02103_));
 sky130_fd_sc_hd__nor2_1 _25169_ (.A(net1712),
    .B(net1107),
    .Y(_02102_));
 sky130_fd_sc_hd__inv_2 _25170_ (.A(_02121_),
    .Y(_02118_));
 sky130_fd_sc_hd__nand2_1 _25171_ (.A(net1047),
    .B(_05935_),
    .Y(_02124_));
 sky130_fd_sc_hd__nand2_1 _25172_ (.A(net1479),
    .B(net1296),
    .Y(_02123_));
 sky130_fd_sc_hd__nand2_1 _25173_ (.A(net1292),
    .B(net1472),
    .Y(_02122_));
 sky130_fd_sc_hd__nand2_1 _25174_ (.A(net1288),
    .B(net1464),
    .Y(_02127_));
 sky130_fd_sc_hd__nand2_1 _25175_ (.A(net1283),
    .B(net1456),
    .Y(_02126_));
 sky130_fd_sc_hd__nand2_1 _25176_ (.A(net1733),
    .B(net1278),
    .Y(_02125_));
 sky130_fd_sc_hd__nand2_1 _25177_ (.A(net1258),
    .B(net1730),
    .Y(_02129_));
 sky130_fd_sc_hd__nand2_1 _25178_ (.A(net1209),
    .B(net1452),
    .Y(_02132_));
 sky130_fd_sc_hd__nand2_1 _25179_ (.A(net1431),
    .B(net1477),
    .Y(_02135_));
 sky130_fd_sc_hd__nand2_1 _25180_ (.A(net1481),
    .B(net1428),
    .Y(_02139_));
 sky130_fd_sc_hd__nor2_1 _25181_ (.A(net1715),
    .B(net1107),
    .Y(_02171_));
 sky130_fd_sc_hd__inv_2 _25182_ (.A(_02151_),
    .Y(_02148_));
 sky130_fd_sc_hd__nand2_1 _25183_ (.A(net1047),
    .B(net1140),
    .Y(_02154_));
 sky130_fd_sc_hd__nand2_1 _25184_ (.A(net1292),
    .B(net1479),
    .Y(_02153_));
 sky130_fd_sc_hd__nand2_1 _25185_ (.A(net1288),
    .B(net1472),
    .Y(_02152_));
 sky130_fd_sc_hd__nand2_1 _25186_ (.A(net1464),
    .B(net1283),
    .Y(_02157_));
 sky130_fd_sc_hd__nand2_1 _25187_ (.A(net1456),
    .B(net1278),
    .Y(_02156_));
 sky130_fd_sc_hd__nand2_1 _25188_ (.A(net1258),
    .B(net1733),
    .Y(_02155_));
 sky130_fd_sc_hd__nor2_1 _25189_ (.A(net1122),
    .B(net1267),
    .Y(_02159_));
 sky130_fd_sc_hd__nor2_1 _25190_ (.A(net1449),
    .B(net1672),
    .Y(_02158_));
 sky130_fd_sc_hd__nand2_1 _25191_ (.A(net1459),
    .B(net1209),
    .Y(_02164_));
 sky130_fd_sc_hd__nand2_1 _25192_ (.A(net1481),
    .B(net1431),
    .Y(_02167_));
 sky130_fd_sc_hd__nor2_1 _25193_ (.A(_20018_),
    .B(net1107),
    .Y(_02170_));
 sky130_fd_sc_hd__inv_2 _25194_ (.A(_02184_),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_1 _25195_ (.A(net1045),
    .B(net1138),
    .Y(_02187_));
 sky130_fd_sc_hd__nand2_1 _25196_ (.A(net1288),
    .B(net1479),
    .Y(_02186_));
 sky130_fd_sc_hd__nand2_1 _25197_ (.A(net1472),
    .B(net1283),
    .Y(_02185_));
 sky130_fd_sc_hd__nor2_1 _25198_ (.A(_19946_),
    .B(net3044),
    .Y(_02189_));
 sky130_fd_sc_hd__nor2_1 _25199_ (.A(_05826_),
    .B(net1125),
    .Y(_02188_));
 sky130_fd_sc_hd__nand2_1 _25200_ (.A(net1466),
    .B(net1210),
    .Y(_02198_));
 sky130_fd_sc_hd__nor2_1 _25201_ (.A(net1722),
    .B(net1107),
    .Y(_02237_));
 sky130_fd_sc_hd__inv_2 _25202_ (.A(_02237_),
    .Y(_02201_));
 sky130_fd_sc_hd__inv_2 _25203_ (.A(_02211_),
    .Y(_02208_));
 sky130_fd_sc_hd__nand2_1 _25204_ (.A(net1045),
    .B(net3042),
    .Y(_02214_));
 sky130_fd_sc_hd__nand2_1 _25205_ (.A(net1479),
    .B(net1283),
    .Y(_02213_));
 sky130_fd_sc_hd__nand2_1 _25207_ (.A(net1472),
    .B(net1280),
    .Y(_02212_));
 sky130_fd_sc_hd__nor2_1 _25208_ (.A(_19946_),
    .B(net1125),
    .Y(_02216_));
 sky130_fd_sc_hd__nor2_1 _25209_ (.A(net1122),
    .B(_05826_),
    .Y(_02215_));
 sky130_fd_sc_hd__nor2_1 _25210_ (.A(net1266),
    .B(net1675),
    .Y(_02223_));
 sky130_fd_sc_hd__nor2_1 _25211_ (.A(net1670),
    .B(net1267),
    .Y(_02222_));
 sky130_fd_sc_hd__nor2_1 _25212_ (.A(net1449),
    .B(net1119),
    .Y(_02221_));
 sky130_fd_sc_hd__nor2_1 _25213_ (.A(_19984_),
    .B(net1737),
    .Y(_02230_));
 sky130_fd_sc_hd__nor2_1 _25214_ (.A(net1211),
    .B(net1116),
    .Y(_02229_));
 sky130_fd_sc_hd__nor2_1 _25215_ (.A(net1438),
    .B(net1113),
    .Y(_02228_));
 sky130_fd_sc_hd__nand2_1 _25216_ (.A(net1481),
    .B(net1135),
    .Y(_02234_));
 sky130_fd_sc_hd__nor2_1 _25217_ (.A(_02983_),
    .B(net1107),
    .Y(_02236_));
 sky130_fd_sc_hd__inv_2 _25218_ (.A(_02236_),
    .Y(_02233_));
 sky130_fd_sc_hd__inv_2 _25219_ (.A(_02245_),
    .Y(_02242_));
 sky130_fd_sc_hd__nand2_1 _25220_ (.A(net1045),
    .B(net1130),
    .Y(_02248_));
 sky130_fd_sc_hd__nand2_1 _25221_ (.A(net1480),
    .B(net1280),
    .Y(_02247_));
 sky130_fd_sc_hd__nand2_1 _25222_ (.A(net1261),
    .B(net1473),
    .Y(_02246_));
 sky130_fd_sc_hd__nor2_1 _25223_ (.A(net1217),
    .B(net1122),
    .Y(_02250_));
 sky130_fd_sc_hd__nor2_1 _25224_ (.A(net1264),
    .B(net1675),
    .Y(_02249_));
 sky130_fd_sc_hd__nor2_1 _25225_ (.A(net1267),
    .B(net1119),
    .Y(_02256_));
 sky130_fd_sc_hd__nor2_1 _25226_ (.A(net1449),
    .B(net1737),
    .Y(_02255_));
 sky130_fd_sc_hd__nor2_1 _25227_ (.A(_19984_),
    .B(net1114),
    .Y(_02265_));
 sky130_fd_sc_hd__nor2_1 _25228_ (.A(net1211),
    .B(net1113),
    .Y(_02264_));
 sky130_fd_sc_hd__nor2_1 _25229_ (.A(net1438),
    .B(net1222),
    .Y(_02263_));
 sky130_fd_sc_hd__nor2_1 _25230_ (.A(_20003_),
    .B(net1107),
    .Y(_02268_));
 sky130_fd_sc_hd__inv_2 _25231_ (.A(_02284_),
    .Y(_02281_));
 sky130_fd_sc_hd__nand2_1 _25232_ (.A(net1045),
    .B(net1127),
    .Y(_02287_));
 sky130_fd_sc_hd__nand2_1 _25233_ (.A(net1261),
    .B(net1480),
    .Y(_02286_));
 sky130_fd_sc_hd__nand2_1 _25234_ (.A(net1275),
    .B(net1473),
    .Y(_02285_));
 sky130_fd_sc_hd__nor2_1 _25235_ (.A(net1217),
    .B(net1675),
    .Y(_02289_));
 sky130_fd_sc_hd__nor2_1 _25236_ (.A(net1670),
    .B(net1264),
    .Y(_02288_));
 sky130_fd_sc_hd__nor2_1 _25237_ (.A(net1265),
    .B(net1119),
    .Y(_02296_));
 sky130_fd_sc_hd__nor2_1 _25238_ (.A(net1737),
    .B(net1269),
    .Y(_02295_));
 sky130_fd_sc_hd__nor2_1 _25239_ (.A(net1449),
    .B(net1114),
    .Y(_02294_));
 sky130_fd_sc_hd__nor2_1 _25240_ (.A(net1212),
    .B(net1113),
    .Y(_02304_));
 sky130_fd_sc_hd__nor2_1 _25241_ (.A(net1211),
    .B(net1222),
    .Y(_02303_));
 sky130_fd_sc_hd__nor2_1 _25242_ (.A(net1438),
    .B(net1106),
    .Y(_02302_));
 sky130_fd_sc_hd__inv_2 _25243_ (.A(_02318_),
    .Y(_02315_));
 sky130_fd_sc_hd__nand2_1 _25244_ (.A(net1045),
    .B(net3044),
    .Y(_02321_));
 sky130_fd_sc_hd__nand2_1 _25245_ (.A(net1275),
    .B(net1480),
    .Y(_02320_));
 sky130_fd_sc_hd__nand2_1 _25246_ (.A(net1473),
    .B(net1272),
    .Y(_02319_));
 sky130_fd_sc_hd__nand2_1 _25247_ (.A(net1256),
    .B(net1465),
    .Y(_02323_));
 sky130_fd_sc_hd__nor2_1 _25248_ (.A(net1735),
    .B(net1265),
    .Y(_02327_));
 sky130_fd_sc_hd__nor2_1 _25249_ (.A(net1269),
    .B(net1114),
    .Y(_02326_));
 sky130_fd_sc_hd__nor2_1 _25250_ (.A(net1450),
    .B(net1110),
    .Y(_02325_));
 sky130_fd_sc_hd__nand2_1 _25251_ (.A(net1482),
    .B(net1447),
    .Y(_02334_));
 sky130_fd_sc_hd__nor2_1 _25252_ (.A(net1211),
    .B(net1106),
    .Y(_02366_));
 sky130_fd_sc_hd__inv_2 _25253_ (.A(_02345_),
    .Y(_02342_));
 sky130_fd_sc_hd__nor2_1 _25254_ (.A(net1740),
    .B(net1122),
    .Y(_02347_));
 sky130_fd_sc_hd__nor2_1 _25255_ (.A(net1220),
    .B(net1675),
    .Y(_02346_));
 sky130_fd_sc_hd__nor2_1 _25256_ (.A(net1670),
    .B(_19932_),
    .Y(_02353_));
 sky130_fd_sc_hd__nor2_1 _25257_ (.A(net1217),
    .B(net1118),
    .Y(_02352_));
 sky130_fd_sc_hd__nor2_1 _25258_ (.A(net1735),
    .B(net1264),
    .Y(_02351_));
 sky130_fd_sc_hd__nor2_1 _25259_ (.A(net1265),
    .B(net1114),
    .Y(_02360_));
 sky130_fd_sc_hd__nor2_1 _25260_ (.A(net1269),
    .B(net1110),
    .Y(_02359_));
 sky130_fd_sc_hd__nor2_1 _25261_ (.A(net1450),
    .B(net1222),
    .Y(_02358_));
 sky130_fd_sc_hd__nor2_1 _25262_ (.A(net1213),
    .B(net1107),
    .Y(_02365_));
 sky130_fd_sc_hd__inv_2 _25263_ (.A(_02375_),
    .Y(_02372_));
 sky130_fd_sc_hd__nor2_1 _25264_ (.A(net1272),
    .B(_06005_),
    .Y(_02378_));
 sky130_fd_sc_hd__nor2_1 _25265_ (.A(net1740),
    .B(net1674),
    .Y(_02377_));
 sky130_fd_sc_hd__nor2_1 _25266_ (.A(net1670),
    .B(net1220),
    .Y(_02376_));
 sky130_fd_sc_hd__nor2_1 _25267_ (.A(_19932_),
    .B(net1118),
    .Y(_02382_));
 sky130_fd_sc_hd__nor2_1 _25268_ (.A(net1264),
    .B(net1114),
    .Y(_02381_));
 sky130_fd_sc_hd__nor2_1 _25269_ (.A(net1265),
    .B(net1110),
    .Y(_02391_));
 sky130_fd_sc_hd__nor2_1 _25270_ (.A(net1269),
    .B(net1222),
    .Y(_02390_));
 sky130_fd_sc_hd__nor2_1 _25271_ (.A(net1450),
    .B(net1106),
    .Y(_02389_));
 sky130_fd_sc_hd__inv_2 _25272_ (.A(_02405_),
    .Y(_02402_));
 sky130_fd_sc_hd__nor2_1 _25273_ (.A(_06005_),
    .B(net1256),
    .Y(_02408_));
 sky130_fd_sc_hd__nor2_1 _25274_ (.A(net1739),
    .B(net1670),
    .Y(_02407_));
 sky130_fd_sc_hd__nor2_1 _25275_ (.A(net1220),
    .B(net1118),
    .Y(_02406_));
 sky130_fd_sc_hd__nor2_1 _25276_ (.A(net1735),
    .B(net1218),
    .Y(_02413_));
 sky130_fd_sc_hd__nor2_1 _25277_ (.A(net1217),
    .B(net1114),
    .Y(_02412_));
 sky130_fd_sc_hd__nor2_1 _25278_ (.A(net1264),
    .B(net1110),
    .Y(_02411_));
 sky130_fd_sc_hd__nand2_1 _25279_ (.A(net1482),
    .B(net1729),
    .Y(_02420_));
 sky130_fd_sc_hd__nor2_1 _25280_ (.A(net1269),
    .B(net1106),
    .Y(_02445_));
 sky130_fd_sc_hd__inv_2 _25281_ (.A(_02430_),
    .Y(_02427_));
 sky130_fd_sc_hd__nor2_1 _25282_ (.A(_06005_),
    .B(net1253),
    .Y(_02433_));
 sky130_fd_sc_hd__nor2_1 _25283_ (.A(net1739),
    .B(net1118),
    .Y(_02432_));
 sky130_fd_sc_hd__nor2_1 _25284_ (.A(net1735),
    .B(net1220),
    .Y(_02431_));
 sky130_fd_sc_hd__nor2_1 _25285_ (.A(net1217),
    .B(net1110),
    .Y(_02437_));
 sky130_fd_sc_hd__nor2_1 _25286_ (.A(net1264),
    .B(net1222),
    .Y(_02436_));
 sky130_fd_sc_hd__nor2_1 _25287_ (.A(net1265),
    .B(net1106),
    .Y(_02444_));
 sky130_fd_sc_hd__inv_2 _25288_ (.A(_02455_),
    .Y(_02452_));
 sky130_fd_sc_hd__nor2_1 _25289_ (.A(net1453),
    .B(_06005_),
    .Y(_02458_));
 sky130_fd_sc_hd__nor2_1 _25290_ (.A(net1739),
    .B(net1735),
    .Y(_02457_));
 sky130_fd_sc_hd__nor2_1 _25291_ (.A(net1220),
    .B(net1114),
    .Y(_02456_));
 sky130_fd_sc_hd__nor2_1 _25292_ (.A(net1218),
    .B(net1110),
    .Y(_02463_));
 sky130_fd_sc_hd__nor2_1 _25293_ (.A(net1217),
    .B(net1222),
    .Y(_02462_));
 sky130_fd_sc_hd__nor2_1 _25294_ (.A(net1264),
    .B(net1106),
    .Y(_02461_));
 sky130_fd_sc_hd__inv_2 _25295_ (.A(_02476_),
    .Y(_02473_));
 sky130_fd_sc_hd__nand2_1 _25296_ (.A(net1045),
    .B(net1735),
    .Y(_02478_));
 sky130_fd_sc_hd__nand2_1 _25297_ (.A(net1482),
    .B(net1465),
    .Y(_02482_));
 sky130_fd_sc_hd__nor2_1 _25298_ (.A(net1217),
    .B(net1106),
    .Y(_02497_));
 sky130_fd_sc_hd__inv_2 _25299_ (.A(_02491_),
    .Y(_02488_));
 sky130_fd_sc_hd__nor2_1 _25300_ (.A(_06005_),
    .B(net1467),
    .Y(_02494_));
 sky130_fd_sc_hd__nor2_1 _25301_ (.A(net1739),
    .B(net1110),
    .Y(_02493_));
 sky130_fd_sc_hd__nor2_1 _25302_ (.A(net1220),
    .B(net1222),
    .Y(_02492_));
 sky130_fd_sc_hd__nor2_1 _25303_ (.A(net1218),
    .B(net1106),
    .Y(_02496_));
 sky130_fd_sc_hd__inv_2 _25304_ (.A(_02510_),
    .Y(_02507_));
 sky130_fd_sc_hd__inv_2 _25305_ (.A(_02540_),
    .Y(_02537_));
 sky130_fd_sc_hd__inv_2 _25306_ (.A(_02499_),
    .Y(_02502_));
 sky130_fd_sc_hd__inv_2 _25307_ (.A(_02520_),
    .Y(_02521_));
 sky130_fd_sc_hd__inv_2 _25308_ (.A(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__inv_2 _25309_ (.A(_02176_),
    .Y(_02178_));
 sky130_fd_sc_hd__inv_2 _25310_ (.A(_02175_),
    .Y(_02205_));
 sky130_fd_sc_hd__inv_2 _25311_ (.A(net2578),
    .Y(_02745_));
 sky130_fd_sc_hd__inv_2 _25312_ (.A(net2579),
    .Y(_02744_));
 sky130_fd_sc_hd__inv_1 _25313_ (.A(_20283_),
    .Y(_06036_));
 sky130_fd_sc_hd__nor2_1 _25314_ (.A(_20293_),
    .B(_06036_),
    .Y(_06037_));
 sky130_fd_sc_hd__inv_1 _25315_ (.A(net2597),
    .Y(_06038_));
 sky130_fd_sc_hd__nand2_1 _25316_ (.A(_20298_),
    .B(_20308_),
    .Y(_06039_));
 sky130_fd_sc_hd__inv_1 _25317_ (.A(_06037_),
    .Y(_06040_));
 sky130_fd_sc_hd__nand2_1 _25318_ (.A(_06039_),
    .B(_06040_),
    .Y(_06041_));
 sky130_fd_sc_hd__o2bb2ai_2 _25319_ (.A1_N(\inst$top.soc.cpu.sink__payload$6[42] ),
    .A2_N(_06037_),
    .B1(_06038_),
    .B2(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__inv_1 _25321_ (.A(\inst$top.soc.cpu.sink__payload$6[41] ),
    .Y(_06043_));
 sky130_fd_sc_hd__o22ai_4 _25322_ (.A1(_06043_),
    .A2(_06040_),
    .B1(net2460),
    .B2(_06041_),
    .Y(_06044_));
 sky130_fd_sc_hd__inv_1 _25324_ (.A(\inst$top.soc.cpu.sink__payload$6[57] ),
    .Y(_06045_));
 sky130_fd_sc_hd__nor2_1 _25325_ (.A(_06037_),
    .B(_06039_),
    .Y(_06046_));
 sky130_fd_sc_hd__nor2_1 _25326_ (.A(_06045_),
    .B(_06046_),
    .Y(\inst$top.soc.cpu.csrf.d_addr[5] ));
 sky130_fd_sc_hd__inv_1 _25327_ (.A(\inst$top.soc.cpu.sink__payload$6[43] ),
    .Y(_06047_));
 sky130_fd_sc_hd__o22ai_2 _25328_ (.A1(_06047_),
    .A2(_06040_),
    .B1(net2450),
    .B2(_06041_),
    .Y(\inst$top.soc.cpu.csrf.d_addr[4] ));
 sky130_fd_sc_hd__inv_1 _25329_ (.A(\inst$top.soc.cpu.sink__payload$6[58] ),
    .Y(_06048_));
 sky130_fd_sc_hd__nor2_2 _25330_ (.A(_06048_),
    .B(_06046_),
    .Y(\inst$top.soc.cpu.csrf.d_addr[6] ));
 sky130_fd_sc_hd__inv_1 _25331_ (.A(\inst$top.soc.cpu.sink__payload$6[59] ),
    .Y(_06049_));
 sky130_fd_sc_hd__nor2_2 _25332_ (.A(_06049_),
    .B(_06046_),
    .Y(\inst$top.soc.cpu.csrf.d_addr[7] ));
 sky130_fd_sc_hd__inv_1 _25333_ (.A(\inst$top.soc.cpu.sink__payload$6[60] ),
    .Y(_06050_));
 sky130_fd_sc_hd__nor2_1 _25334_ (.A(_06050_),
    .B(_06046_),
    .Y(\inst$top.soc.cpu.csrf.d_addr[8] ));
 sky130_fd_sc_hd__inv_1 _25335_ (.A(\inst$top.soc.cpu.sink__payload$6[62] ),
    .Y(_06051_));
 sky130_fd_sc_hd__nor2_1 _25336_ (.A(_06051_),
    .B(_06046_),
    .Y(\inst$top.soc.cpu.csrf.d_addr[10] ));
 sky130_fd_sc_hd__inv_1 _25337_ (.A(\inst$top.soc.cpu.sink__payload$6[61] ),
    .Y(_06052_));
 sky130_fd_sc_hd__nor2_1 _25338_ (.A(_06052_),
    .B(_06046_),
    .Y(\inst$top.soc.cpu.csrf.d_addr[9] ));
 sky130_fd_sc_hd__nor2_1 _25341_ (.A(\inst$top.soc.cpu.gprf.mem[15][0] ),
    .B(net2461),
    .Y(_06055_));
 sky130_fd_sc_hd__o21ai_0 _25347_ (.A1(net2653),
    .A2(\inst$top.soc.cpu.gprf.mem[14][0] ),
    .B1(net2616),
    .Y(_06061_));
 sky130_fd_sc_hd__nor2_1 _25350_ (.A(net2639),
    .B(net2484),
    .Y(_06064_));
 sky130_fd_sc_hd__a221oi_1 _25355_ (.A1(net2506),
    .A2(\inst$top.soc.cpu.gprf.mem[12][0] ),
    .B1(net1945),
    .B2(\inst$top.soc.cpu.gprf.mem[13][0] ),
    .C1(net2451),
    .Y(_06069_));
 sky130_fd_sc_hd__o21ai_0 _25356_ (.A1(_06055_),
    .A2(_06061_),
    .B1(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__nor2_1 _25359_ (.A(\inst$top.soc.cpu.gprf.mem[11][0] ),
    .B(net2462),
    .Y(_06073_));
 sky130_fd_sc_hd__o21ai_0 _25364_ (.A1(net2653),
    .A2(\inst$top.soc.cpu.gprf.mem[10][0] ),
    .B1(net2617),
    .Y(_06078_));
 sky130_fd_sc_hd__a221oi_1 _25370_ (.A1(net2507),
    .A2(\inst$top.soc.cpu.gprf.mem[8][0] ),
    .B1(net1945),
    .B2(\inst$top.soc.cpu.gprf.mem[9][0] ),
    .C1(net2607),
    .Y(_06084_));
 sky130_fd_sc_hd__o21ai_0 _25371_ (.A1(_06073_),
    .A2(_06078_),
    .B1(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__nand3_1 _25374_ (.A(_06070_),
    .B(_06085_),
    .C(net2600),
    .Y(_06088_));
 sky130_fd_sc_hd__nor2_1 _25376_ (.A(\inst$top.soc.cpu.gprf.mem[7][0] ),
    .B(net2463),
    .Y(_06090_));
 sky130_fd_sc_hd__o21ai_0 _25379_ (.A1(net2686),
    .A2(\inst$top.soc.cpu.gprf.mem[6][0] ),
    .B1(net2618),
    .Y(_06093_));
 sky130_fd_sc_hd__a22oi_1 _25385_ (.A1(net2508),
    .A2(\inst$top.soc.cpu.gprf.mem[4][0] ),
    .B1(net1947),
    .B2(\inst$top.soc.cpu.gprf.mem[5][0] ),
    .Y(_06099_));
 sky130_fd_sc_hd__o21ai_0 _25386_ (.A1(_06090_),
    .A2(_06093_),
    .B1(_06099_),
    .Y(_06100_));
 sky130_fd_sc_hd__nor2_1 _25387_ (.A(net2601),
    .B(net2454),
    .Y(_06101_));
 sky130_fd_sc_hd__nand2_1 _25390_ (.A(_06100_),
    .B(net1942),
    .Y(_06104_));
 sky130_fd_sc_hd__nor2_1 _25393_ (.A(\inst$top.soc.cpu.gprf.mem[3][0] ),
    .B(net2463),
    .Y(_06107_));
 sky130_fd_sc_hd__o21ai_0 _25396_ (.A1(net2686),
    .A2(\inst$top.soc.cpu.gprf.mem[2][0] ),
    .B1(net2618),
    .Y(_06110_));
 sky130_fd_sc_hd__a22oi_1 _25399_ (.A1(net2505),
    .A2(\inst$top.soc.cpu.gprf.mem[0][0] ),
    .B1(net1944),
    .B2(\inst$top.soc.cpu.gprf.mem[1][0] ),
    .Y(_06113_));
 sky130_fd_sc_hd__o21ai_0 _25400_ (.A1(_06107_),
    .A2(_06110_),
    .B1(_06113_),
    .Y(_06114_));
 sky130_fd_sc_hd__a21oi_1 _25404_ (.A1(_06114_),
    .A2(net2496),
    .B1(net2591),
    .Y(_06118_));
 sky130_fd_sc_hd__nor2_1 _25407_ (.A(\inst$top.soc.cpu.gprf.mem[19][0] ),
    .B(net2462),
    .Y(_06121_));
 sky130_fd_sc_hd__o21ai_0 _25410_ (.A1(net2655),
    .A2(\inst$top.soc.cpu.gprf.mem[18][0] ),
    .B1(net2617),
    .Y(_06124_));
 sky130_fd_sc_hd__a22oi_1 _25413_ (.A1(net2507),
    .A2(\inst$top.soc.cpu.gprf.mem[16][0] ),
    .B1(net1946),
    .B2(\inst$top.soc.cpu.gprf.mem[17][0] ),
    .Y(_06127_));
 sky130_fd_sc_hd__o21ai_0 _25414_ (.A1(_06121_),
    .A2(_06124_),
    .B1(_06127_),
    .Y(_06128_));
 sky130_fd_sc_hd__nor2_1 _25415_ (.A(\inst$top.soc.cpu.gprf.mem[23][0] ),
    .B(net2462),
    .Y(_06129_));
 sky130_fd_sc_hd__o21ai_0 _25416_ (.A1(net2655),
    .A2(\inst$top.soc.cpu.gprf.mem[22][0] ),
    .B1(net2617),
    .Y(_06130_));
 sky130_fd_sc_hd__a22oi_1 _25417_ (.A1(net2506),
    .A2(\inst$top.soc.cpu.gprf.mem[20][0] ),
    .B1(net1946),
    .B2(\inst$top.soc.cpu.gprf.mem[21][0] ),
    .Y(_06131_));
 sky130_fd_sc_hd__o21ai_0 _25418_ (.A1(_06129_),
    .A2(_06130_),
    .B1(_06131_),
    .Y(_06132_));
 sky130_fd_sc_hd__nor2_1 _25422_ (.A(net2655),
    .B(\inst$top.soc.cpu.gprf.mem[26][0] ),
    .Y(_06136_));
 sky130_fd_sc_hd__nor2_1 _25423_ (.A(_20261_),
    .B(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__o21ai_0 _25424_ (.A1(net2464),
    .A2(\inst$top.soc.cpu.gprf.mem[27][0] ),
    .B1(_06137_),
    .Y(_06138_));
 sky130_fd_sc_hd__a221oi_1 _25425_ (.A1(net2508),
    .A2(\inst$top.soc.cpu.gprf.mem[24][0] ),
    .B1(net1947),
    .B2(\inst$top.soc.cpu.gprf.mem[25][0] ),
    .C1(net2607),
    .Y(_06139_));
 sky130_fd_sc_hd__nor2_1 _25426_ (.A(\inst$top.soc.cpu.gprf.mem[31][0] ),
    .B(net2463),
    .Y(_06140_));
 sky130_fd_sc_hd__o21ai_0 _25427_ (.A1(net2655),
    .A2(\inst$top.soc.cpu.gprf.mem[30][0] ),
    .B1(net2617),
    .Y(_06141_));
 sky130_fd_sc_hd__nand2_1 _25428_ (.A(net2508),
    .B(\inst$top.soc.cpu.gprf.mem[28][0] ),
    .Y(_06142_));
 sky130_fd_sc_hd__nand2_1 _25429_ (.A(net1947),
    .B(\inst$top.soc.cpu.gprf.mem[29][0] ),
    .Y(_06143_));
 sky130_fd_sc_hd__o211ai_1 _25430_ (.A1(_06140_),
    .A2(_06141_),
    .B1(_06142_),
    .C1(_06143_),
    .Y(_06144_));
 sky130_fd_sc_hd__o21ai_0 _25431_ (.A1(net2452),
    .A2(_06144_),
    .B1(net2597),
    .Y(_06145_));
 sky130_fd_sc_hd__a21oi_1 _25432_ (.A1(_06138_),
    .A2(_06139_),
    .B1(_06145_),
    .Y(_06146_));
 sky130_fd_sc_hd__a221oi_1 _25433_ (.A1(net2496),
    .A2(_06128_),
    .B1(_06132_),
    .B2(net1943),
    .C1(_06146_),
    .Y(_06147_));
 sky130_fd_sc_hd__a32oi_1 _25436_ (.A1(_06088_),
    .A2(_06104_),
    .A3(_06118_),
    .B1(_06147_),
    .B2(net2591),
    .Y(_00000_));
 sky130_fd_sc_hd__nor2_1 _25437_ (.A(\inst$top.soc.cpu.gprf.mem[15][1] ),
    .B(net2461),
    .Y(_06150_));
 sky130_fd_sc_hd__o21ai_0 _25438_ (.A1(net2653),
    .A2(\inst$top.soc.cpu.gprf.mem[14][1] ),
    .B1(net2616),
    .Y(_06151_));
 sky130_fd_sc_hd__a221oi_1 _25439_ (.A1(net2506),
    .A2(\inst$top.soc.cpu.gprf.mem[12][1] ),
    .B1(net1945),
    .B2(\inst$top.soc.cpu.gprf.mem[13][1] ),
    .C1(net2451),
    .Y(_06152_));
 sky130_fd_sc_hd__o21ai_0 _25440_ (.A1(_06150_),
    .A2(_06151_),
    .B1(_06152_),
    .Y(_06153_));
 sky130_fd_sc_hd__nor2_1 _25441_ (.A(\inst$top.soc.cpu.gprf.mem[11][1] ),
    .B(net2461),
    .Y(_06154_));
 sky130_fd_sc_hd__o21ai_0 _25442_ (.A1(net2653),
    .A2(\inst$top.soc.cpu.gprf.mem[10][1] ),
    .B1(net2616),
    .Y(_06155_));
 sky130_fd_sc_hd__a221oi_1 _25443_ (.A1(net2506),
    .A2(\inst$top.soc.cpu.gprf.mem[8][1] ),
    .B1(net1945),
    .B2(\inst$top.soc.cpu.gprf.mem[9][1] ),
    .C1(net2607),
    .Y(_06156_));
 sky130_fd_sc_hd__o21ai_0 _25444_ (.A1(_06154_),
    .A2(_06155_),
    .B1(_06156_),
    .Y(_06157_));
 sky130_fd_sc_hd__nand3_1 _25445_ (.A(_06153_),
    .B(_06157_),
    .C(net2600),
    .Y(_06158_));
 sky130_fd_sc_hd__nor2_1 _25446_ (.A(\inst$top.soc.cpu.gprf.mem[7][1] ),
    .B(net2463),
    .Y(_06159_));
 sky130_fd_sc_hd__o21ai_0 _25447_ (.A1(net2652),
    .A2(\inst$top.soc.cpu.gprf.mem[6][1] ),
    .B1(net2618),
    .Y(_06160_));
 sky130_fd_sc_hd__a22oi_1 _25448_ (.A1(net2505),
    .A2(\inst$top.soc.cpu.gprf.mem[4][1] ),
    .B1(net1944),
    .B2(\inst$top.soc.cpu.gprf.mem[5][1] ),
    .Y(_06161_));
 sky130_fd_sc_hd__o21ai_0 _25449_ (.A1(_06159_),
    .A2(_06160_),
    .B1(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__nand2_1 _25450_ (.A(_06162_),
    .B(net1942),
    .Y(_06163_));
 sky130_fd_sc_hd__nor2_1 _25451_ (.A(\inst$top.soc.cpu.gprf.mem[3][1] ),
    .B(net2463),
    .Y(_06164_));
 sky130_fd_sc_hd__o21ai_0 _25452_ (.A1(net2686),
    .A2(\inst$top.soc.cpu.gprf.mem[2][1] ),
    .B1(net2618),
    .Y(_06165_));
 sky130_fd_sc_hd__a22oi_1 _25453_ (.A1(net2505),
    .A2(\inst$top.soc.cpu.gprf.mem[0][1] ),
    .B1(net1944),
    .B2(\inst$top.soc.cpu.gprf.mem[1][1] ),
    .Y(_06166_));
 sky130_fd_sc_hd__o21ai_0 _25454_ (.A1(_06164_),
    .A2(_06165_),
    .B1(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__a21oi_1 _25455_ (.A1(_06167_),
    .A2(net2496),
    .B1(net2591),
    .Y(_06168_));
 sky130_fd_sc_hd__nor2_1 _25457_ (.A(\inst$top.soc.cpu.gprf.mem[19][1] ),
    .B(net2462),
    .Y(_06170_));
 sky130_fd_sc_hd__o21ai_0 _25460_ (.A1(net2653),
    .A2(\inst$top.soc.cpu.gprf.mem[18][1] ),
    .B1(net2617),
    .Y(_06173_));
 sky130_fd_sc_hd__a22oi_1 _25463_ (.A1(net2506),
    .A2(\inst$top.soc.cpu.gprf.mem[16][1] ),
    .B1(net1945),
    .B2(\inst$top.soc.cpu.gprf.mem[17][1] ),
    .Y(_06176_));
 sky130_fd_sc_hd__o21ai_0 _25464_ (.A1(_06170_),
    .A2(_06173_),
    .B1(_06176_),
    .Y(_06177_));
 sky130_fd_sc_hd__nor2_1 _25466_ (.A(\inst$top.soc.cpu.gprf.mem[23][1] ),
    .B(net2462),
    .Y(_06179_));
 sky130_fd_sc_hd__o21ai_0 _25469_ (.A1(net2653),
    .A2(\inst$top.soc.cpu.gprf.mem[22][1] ),
    .B1(net2617),
    .Y(_06182_));
 sky130_fd_sc_hd__a22oi_1 _25472_ (.A1(net2506),
    .A2(\inst$top.soc.cpu.gprf.mem[20][1] ),
    .B1(net1945),
    .B2(\inst$top.soc.cpu.gprf.mem[21][1] ),
    .Y(_06185_));
 sky130_fd_sc_hd__o21ai_0 _25473_ (.A1(_06179_),
    .A2(_06182_),
    .B1(_06185_),
    .Y(_06186_));
 sky130_fd_sc_hd__a221oi_1 _25476_ (.A1(_06177_),
    .A2(net2496),
    .B1(net1943),
    .B2(_06186_),
    .C1(net2450),
    .Y(_06189_));
 sky130_fd_sc_hd__nor2_1 _25478_ (.A(\inst$top.soc.cpu.gprf.mem[31][1] ),
    .B(net2463),
    .Y(_06191_));
 sky130_fd_sc_hd__o21ai_0 _25481_ (.A1(net2652),
    .A2(\inst$top.soc.cpu.gprf.mem[30][1] ),
    .B1(net2616),
    .Y(_06194_));
 sky130_fd_sc_hd__a221oi_1 _25485_ (.A1(net2505),
    .A2(\inst$top.soc.cpu.gprf.mem[28][1] ),
    .B1(net1944),
    .B2(\inst$top.soc.cpu.gprf.mem[29][1] ),
    .C1(net2452),
    .Y(_06198_));
 sky130_fd_sc_hd__o21ai_0 _25486_ (.A1(_06191_),
    .A2(_06194_),
    .B1(_06198_),
    .Y(_06199_));
 sky130_fd_sc_hd__nor2_1 _25488_ (.A(\inst$top.soc.cpu.gprf.mem[27][1] ),
    .B(net2461),
    .Y(_06201_));
 sky130_fd_sc_hd__o21ai_0 _25491_ (.A1(net2652),
    .A2(\inst$top.soc.cpu.gprf.mem[26][1] ),
    .B1(net2616),
    .Y(_06204_));
 sky130_fd_sc_hd__a221oi_1 _25495_ (.A1(net2505),
    .A2(\inst$top.soc.cpu.gprf.mem[24][1] ),
    .B1(net1944),
    .B2(\inst$top.soc.cpu.gprf.mem[25][1] ),
    .C1(net2607),
    .Y(_06208_));
 sky130_fd_sc_hd__o21ai_0 _25496_ (.A1(_06201_),
    .A2(_06204_),
    .B1(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__nand3_1 _25498_ (.A(_06199_),
    .B(_06209_),
    .C(net2606),
    .Y(_06211_));
 sky130_fd_sc_hd__a32oi_1 _25499_ (.A1(_06158_),
    .A2(_06163_),
    .A3(_06168_),
    .B1(_06189_),
    .B2(_06211_),
    .Y(_00011_));
 sky130_fd_sc_hd__nor2_1 _25500_ (.A(\inst$top.soc.cpu.gprf.mem[11][2] ),
    .B(net2461),
    .Y(_06212_));
 sky130_fd_sc_hd__o21ai_0 _25503_ (.A1(net2652),
    .A2(\inst$top.soc.cpu.gprf.mem[10][2] ),
    .B1(net2616),
    .Y(_06215_));
 sky130_fd_sc_hd__a221oi_1 _25506_ (.A1(net2506),
    .A2(\inst$top.soc.cpu.gprf.mem[8][2] ),
    .B1(net1945),
    .B2(\inst$top.soc.cpu.gprf.mem[9][2] ),
    .C1(net2607),
    .Y(_06218_));
 sky130_fd_sc_hd__o21ai_0 _25507_ (.A1(_06212_),
    .A2(_06215_),
    .B1(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__nor2_1 _25508_ (.A(\inst$top.soc.cpu.gprf.mem[15][2] ),
    .B(net2461),
    .Y(_06220_));
 sky130_fd_sc_hd__o21ai_0 _25509_ (.A1(net2652),
    .A2(\inst$top.soc.cpu.gprf.mem[14][2] ),
    .B1(net2616),
    .Y(_06221_));
 sky130_fd_sc_hd__a221oi_1 _25511_ (.A1(net2505),
    .A2(\inst$top.soc.cpu.gprf.mem[12][2] ),
    .B1(net1944),
    .B2(\inst$top.soc.cpu.gprf.mem[13][2] ),
    .C1(net2452),
    .Y(_06223_));
 sky130_fd_sc_hd__o21ai_0 _25512_ (.A1(_06220_),
    .A2(_06221_),
    .B1(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__nand3_1 _25513_ (.A(_06219_),
    .B(_06224_),
    .C(net2606),
    .Y(_06225_));
 sky130_fd_sc_hd__nor2_1 _25515_ (.A(\inst$top.soc.cpu.gprf.mem[7][2] ),
    .B(net2463),
    .Y(_06227_));
 sky130_fd_sc_hd__o21ai_0 _25516_ (.A1(net2686),
    .A2(\inst$top.soc.cpu.gprf.mem[6][2] ),
    .B1(net2618),
    .Y(_06228_));
 sky130_fd_sc_hd__a22oi_1 _25518_ (.A1(net2505),
    .A2(\inst$top.soc.cpu.gprf.mem[4][2] ),
    .B1(net1944),
    .B2(\inst$top.soc.cpu.gprf.mem[5][2] ),
    .Y(_06230_));
 sky130_fd_sc_hd__o21ai_0 _25519_ (.A1(_06227_),
    .A2(_06228_),
    .B1(_06230_),
    .Y(_06231_));
 sky130_fd_sc_hd__nand2_1 _25520_ (.A(_06231_),
    .B(net1942),
    .Y(_06232_));
 sky130_fd_sc_hd__nor2_1 _25521_ (.A(\inst$top.soc.cpu.gprf.mem[3][2] ),
    .B(net2463),
    .Y(_06233_));
 sky130_fd_sc_hd__o21ai_0 _25524_ (.A1(net2686),
    .A2(\inst$top.soc.cpu.gprf.mem[2][2] ),
    .B1(net2618),
    .Y(_06236_));
 sky130_fd_sc_hd__a22oi_1 _25525_ (.A1(net2505),
    .A2(\inst$top.soc.cpu.gprf.mem[0][2] ),
    .B1(net1944),
    .B2(\inst$top.soc.cpu.gprf.mem[1][2] ),
    .Y(_06237_));
 sky130_fd_sc_hd__o21ai_0 _25526_ (.A1(_06233_),
    .A2(_06236_),
    .B1(_06237_),
    .Y(_06238_));
 sky130_fd_sc_hd__a21oi_1 _25527_ (.A1(_06238_),
    .A2(net2496),
    .B1(net2591),
    .Y(_06239_));
 sky130_fd_sc_hd__nor2_1 _25528_ (.A(\inst$top.soc.cpu.gprf.mem[19][2] ),
    .B(net2461),
    .Y(_06240_));
 sky130_fd_sc_hd__o21ai_0 _25529_ (.A1(net2652),
    .A2(\inst$top.soc.cpu.gprf.mem[18][2] ),
    .B1(net2616),
    .Y(_06241_));
 sky130_fd_sc_hd__a22oi_1 _25530_ (.A1(net2506),
    .A2(\inst$top.soc.cpu.gprf.mem[16][2] ),
    .B1(net1945),
    .B2(\inst$top.soc.cpu.gprf.mem[17][2] ),
    .Y(_06242_));
 sky130_fd_sc_hd__o21ai_0 _25531_ (.A1(_06240_),
    .A2(_06241_),
    .B1(_06242_),
    .Y(_06243_));
 sky130_fd_sc_hd__nor2_1 _25532_ (.A(\inst$top.soc.cpu.gprf.mem[23][2] ),
    .B(net2461),
    .Y(_06244_));
 sky130_fd_sc_hd__o21ai_0 _25533_ (.A1(net2652),
    .A2(\inst$top.soc.cpu.gprf.mem[22][2] ),
    .B1(net2616),
    .Y(_06245_));
 sky130_fd_sc_hd__a22oi_1 _25534_ (.A1(net2506),
    .A2(\inst$top.soc.cpu.gprf.mem[20][2] ),
    .B1(net1945),
    .B2(\inst$top.soc.cpu.gprf.mem[21][2] ),
    .Y(_06246_));
 sky130_fd_sc_hd__o21ai_0 _25535_ (.A1(_06244_),
    .A2(_06245_),
    .B1(_06246_),
    .Y(_06247_));
 sky130_fd_sc_hd__nor2_1 _25536_ (.A(net2652),
    .B(\inst$top.soc.cpu.gprf.mem[26][2] ),
    .Y(_06248_));
 sky130_fd_sc_hd__nor2_1 _25537_ (.A(_20261_),
    .B(_06248_),
    .Y(_06249_));
 sky130_fd_sc_hd__o21ai_0 _25538_ (.A1(net2461),
    .A2(\inst$top.soc.cpu.gprf.mem[27][2] ),
    .B1(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__a221oi_1 _25539_ (.A1(net2505),
    .A2(\inst$top.soc.cpu.gprf.mem[24][2] ),
    .B1(net1944),
    .B2(\inst$top.soc.cpu.gprf.mem[25][2] ),
    .C1(net2607),
    .Y(_06251_));
 sky130_fd_sc_hd__nor2_1 _25540_ (.A(\inst$top.soc.cpu.gprf.mem[31][2] ),
    .B(net2461),
    .Y(_06252_));
 sky130_fd_sc_hd__o21ai_0 _25541_ (.A1(net2652),
    .A2(\inst$top.soc.cpu.gprf.mem[30][2] ),
    .B1(net2616),
    .Y(_06253_));
 sky130_fd_sc_hd__nand2_1 _25542_ (.A(net2505),
    .B(\inst$top.soc.cpu.gprf.mem[28][2] ),
    .Y(_06254_));
 sky130_fd_sc_hd__nand2_1 _25543_ (.A(net1944),
    .B(\inst$top.soc.cpu.gprf.mem[29][2] ),
    .Y(_06255_));
 sky130_fd_sc_hd__o211ai_1 _25544_ (.A1(_06252_),
    .A2(_06253_),
    .B1(_06254_),
    .C1(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__o21ai_0 _25545_ (.A1(net2452),
    .A2(_06256_),
    .B1(net2597),
    .Y(_06257_));
 sky130_fd_sc_hd__a21oi_1 _25546_ (.A1(_06250_),
    .A2(_06251_),
    .B1(_06257_),
    .Y(_06258_));
 sky130_fd_sc_hd__a221oi_1 _25547_ (.A1(net2496),
    .A2(_06243_),
    .B1(net1943),
    .B2(_06247_),
    .C1(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__a32oi_1 _25548_ (.A1(_06225_),
    .A2(_06232_),
    .A3(_06239_),
    .B1(_06259_),
    .B2(net2591),
    .Y(_00022_));
 sky130_fd_sc_hd__nor2_1 _25549_ (.A(\inst$top.soc.cpu.gprf.mem[31][3] ),
    .B(net2483),
    .Y(_06260_));
 sky130_fd_sc_hd__o21ai_0 _25550_ (.A1(net2675),
    .A2(\inst$top.soc.cpu.gprf.mem[30][3] ),
    .B1(net2637),
    .Y(_06261_));
 sky130_fd_sc_hd__a221oi_1 _25552_ (.A1(net2527),
    .A2(\inst$top.soc.cpu.gprf.mem[28][3] ),
    .B1(net1967),
    .B2(\inst$top.soc.cpu.gprf.mem[29][3] ),
    .C1(net2457),
    .Y(_06263_));
 sky130_fd_sc_hd__o21ai_0 _25553_ (.A1(_06260_),
    .A2(_06261_),
    .B1(_06263_),
    .Y(_06264_));
 sky130_fd_sc_hd__nor2_1 _25554_ (.A(\inst$top.soc.cpu.gprf.mem[27][3] ),
    .B(net2483),
    .Y(_06265_));
 sky130_fd_sc_hd__o21ai_0 _25555_ (.A1(net2675),
    .A2(\inst$top.soc.cpu.gprf.mem[26][3] ),
    .B1(net2637),
    .Y(_06266_));
 sky130_fd_sc_hd__a221oi_1 _25556_ (.A1(net2527),
    .A2(\inst$top.soc.cpu.gprf.mem[24][3] ),
    .B1(net1967),
    .B2(\inst$top.soc.cpu.gprf.mem[25][3] ),
    .C1(net2612),
    .Y(_06267_));
 sky130_fd_sc_hd__o21ai_0 _25557_ (.A1(_06265_),
    .A2(_06266_),
    .B1(_06267_),
    .Y(_06268_));
 sky130_fd_sc_hd__nand3_1 _25558_ (.A(_06264_),
    .B(_06268_),
    .C(net2603),
    .Y(_06269_));
 sky130_fd_sc_hd__nor2_1 _25559_ (.A(\inst$top.soc.cpu.gprf.mem[23][3] ),
    .B(net2482),
    .Y(_06270_));
 sky130_fd_sc_hd__o21ai_0 _25560_ (.A1(net2676),
    .A2(\inst$top.soc.cpu.gprf.mem[22][3] ),
    .B1(net2635),
    .Y(_06271_));
 sky130_fd_sc_hd__a22oi_1 _25561_ (.A1(net2528),
    .A2(\inst$top.soc.cpu.gprf.mem[20][3] ),
    .B1(net1968),
    .B2(\inst$top.soc.cpu.gprf.mem[21][3] ),
    .Y(_06272_));
 sky130_fd_sc_hd__o21ai_0 _25562_ (.A1(_06270_),
    .A2(_06271_),
    .B1(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__nand2_1 _25563_ (.A(_06273_),
    .B(net1938),
    .Y(_06274_));
 sky130_fd_sc_hd__nor2_1 _25565_ (.A(\inst$top.soc.cpu.gprf.mem[19][3] ),
    .B(net2482),
    .Y(_06276_));
 sky130_fd_sc_hd__o21ai_0 _25566_ (.A1(net2675),
    .A2(\inst$top.soc.cpu.gprf.mem[18][3] ),
    .B1(net2634),
    .Y(_06277_));
 sky130_fd_sc_hd__a22oi_1 _25567_ (.A1(net2527),
    .A2(\inst$top.soc.cpu.gprf.mem[16][3] ),
    .B1(net1967),
    .B2(\inst$top.soc.cpu.gprf.mem[17][3] ),
    .Y(_06278_));
 sky130_fd_sc_hd__o21ai_0 _25568_ (.A1(_06276_),
    .A2(_06277_),
    .B1(_06278_),
    .Y(_06279_));
 sky130_fd_sc_hd__a21oi_1 _25569_ (.A1(_06279_),
    .A2(net2500),
    .B1(net2447),
    .Y(_06280_));
 sky130_fd_sc_hd__nor2_1 _25571_ (.A(\inst$top.soc.cpu.gprf.mem[7][3] ),
    .B(net2480),
    .Y(_06282_));
 sky130_fd_sc_hd__o21ai_0 _25572_ (.A1(net2675),
    .A2(\inst$top.soc.cpu.gprf.mem[6][3] ),
    .B1(net2637),
    .Y(_06283_));
 sky130_fd_sc_hd__a22oi_1 _25573_ (.A1(net2527),
    .A2(\inst$top.soc.cpu.gprf.mem[4][3] ),
    .B1(net1967),
    .B2(\inst$top.soc.cpu.gprf.mem[5][3] ),
    .Y(_06284_));
 sky130_fd_sc_hd__o21ai_0 _25574_ (.A1(_06282_),
    .A2(_06283_),
    .B1(_06284_),
    .Y(_06285_));
 sky130_fd_sc_hd__nor2_1 _25578_ (.A(\inst$top.soc.cpu.gprf.mem[3][3] ),
    .B(net2483),
    .Y(_06289_));
 sky130_fd_sc_hd__o21ai_0 _25579_ (.A1(net2675),
    .A2(\inst$top.soc.cpu.gprf.mem[2][3] ),
    .B1(net2637),
    .Y(_06290_));
 sky130_fd_sc_hd__a22oi_1 _25580_ (.A1(net2527),
    .A2(\inst$top.soc.cpu.gprf.mem[0][3] ),
    .B1(net1967),
    .B2(\inst$top.soc.cpu.gprf.mem[1][3] ),
    .Y(_06291_));
 sky130_fd_sc_hd__o21ai_0 _25581_ (.A1(_06289_),
    .A2(_06290_),
    .B1(_06291_),
    .Y(_06292_));
 sky130_fd_sc_hd__a221oi_1 _25582_ (.A1(_06285_),
    .A2(net1938),
    .B1(net2501),
    .B2(_06292_),
    .C1(net2593),
    .Y(_06293_));
 sky130_fd_sc_hd__nor2_1 _25583_ (.A(\inst$top.soc.cpu.gprf.mem[15][3] ),
    .B(net2480),
    .Y(_06294_));
 sky130_fd_sc_hd__o21ai_0 _25584_ (.A1(net2675),
    .A2(\inst$top.soc.cpu.gprf.mem[14][3] ),
    .B1(net2634),
    .Y(_06295_));
 sky130_fd_sc_hd__a221oi_1 _25585_ (.A1(net2527),
    .A2(\inst$top.soc.cpu.gprf.mem[12][3] ),
    .B1(net1967),
    .B2(\inst$top.soc.cpu.gprf.mem[13][3] ),
    .C1(net2456),
    .Y(_06296_));
 sky130_fd_sc_hd__o21ai_0 _25586_ (.A1(_06294_),
    .A2(_06295_),
    .B1(_06296_),
    .Y(_06297_));
 sky130_fd_sc_hd__nor2_1 _25587_ (.A(\inst$top.soc.cpu.gprf.mem[11][3] ),
    .B(net2480),
    .Y(_06298_));
 sky130_fd_sc_hd__o21ai_0 _25588_ (.A1(net2675),
    .A2(\inst$top.soc.cpu.gprf.mem[10][3] ),
    .B1(net2634),
    .Y(_06299_));
 sky130_fd_sc_hd__a221oi_1 _25589_ (.A1(net2527),
    .A2(\inst$top.soc.cpu.gprf.mem[8][3] ),
    .B1(net1967),
    .B2(\inst$top.soc.cpu.gprf.mem[9][3] ),
    .C1(net2612),
    .Y(_06300_));
 sky130_fd_sc_hd__o21ai_0 _25590_ (.A1(_06298_),
    .A2(_06299_),
    .B1(_06300_),
    .Y(_06301_));
 sky130_fd_sc_hd__nand3_1 _25591_ (.A(_06297_),
    .B(_06301_),
    .C(net2603),
    .Y(_06302_));
 sky130_fd_sc_hd__a32oi_1 _25592_ (.A1(_06269_),
    .A2(_06274_),
    .A3(_06280_),
    .B1(_06293_),
    .B2(_06302_),
    .Y(_00025_));
 sky130_fd_sc_hd__nor2_1 _25594_ (.A(\inst$top.soc.cpu.gprf.mem[11][4] ),
    .B(net2467),
    .Y(_06304_));
 sky130_fd_sc_hd__o21ai_0 _25595_ (.A1(net2657),
    .A2(\inst$top.soc.cpu.gprf.mem[10][4] ),
    .B1(net2621),
    .Y(_06305_));
 sky130_fd_sc_hd__a221oi_1 _25596_ (.A1(net2510),
    .A2(\inst$top.soc.cpu.gprf.mem[8][4] ),
    .B1(net1949),
    .B2(\inst$top.soc.cpu.gprf.mem[9][4] ),
    .C1(net2610),
    .Y(_06306_));
 sky130_fd_sc_hd__o21ai_0 _25597_ (.A1(_06304_),
    .A2(_06305_),
    .B1(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__nor2_1 _25598_ (.A(\inst$top.soc.cpu.gprf.mem[15][4] ),
    .B(net2466),
    .Y(_06308_));
 sky130_fd_sc_hd__o21ai_0 _25599_ (.A1(net2657),
    .A2(\inst$top.soc.cpu.gprf.mem[14][4] ),
    .B1(net2621),
    .Y(_06309_));
 sky130_fd_sc_hd__a221oi_1 _25600_ (.A1(net2510),
    .A2(\inst$top.soc.cpu.gprf.mem[12][4] ),
    .B1(net1949),
    .B2(\inst$top.soc.cpu.gprf.mem[13][4] ),
    .C1(net2453),
    .Y(_06310_));
 sky130_fd_sc_hd__o21ai_0 _25601_ (.A1(_06308_),
    .A2(_06309_),
    .B1(_06310_),
    .Y(_06311_));
 sky130_fd_sc_hd__nand3_1 _25602_ (.A(_06307_),
    .B(_06311_),
    .C(net2600),
    .Y(_06312_));
 sky130_fd_sc_hd__nor2_1 _25603_ (.A(\inst$top.soc.cpu.gprf.mem[7][4] ),
    .B(net2466),
    .Y(_06313_));
 sky130_fd_sc_hd__o21ai_0 _25604_ (.A1(net2657),
    .A2(\inst$top.soc.cpu.gprf.mem[6][4] ),
    .B1(net2621),
    .Y(_06314_));
 sky130_fd_sc_hd__a22oi_1 _25605_ (.A1(net2510),
    .A2(\inst$top.soc.cpu.gprf.mem[4][4] ),
    .B1(net1949),
    .B2(\inst$top.soc.cpu.gprf.mem[5][4] ),
    .Y(_06315_));
 sky130_fd_sc_hd__o21ai_0 _25606_ (.A1(_06313_),
    .A2(_06314_),
    .B1(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__nand2_1 _25607_ (.A(_06316_),
    .B(net1934),
    .Y(_06317_));
 sky130_fd_sc_hd__nor2_1 _25608_ (.A(\inst$top.soc.cpu.gprf.mem[3][4] ),
    .B(net2466),
    .Y(_06318_));
 sky130_fd_sc_hd__o21ai_0 _25609_ (.A1(net2657),
    .A2(\inst$top.soc.cpu.gprf.mem[2][4] ),
    .B1(net2621),
    .Y(_06319_));
 sky130_fd_sc_hd__a22oi_1 _25611_ (.A1(net2510),
    .A2(\inst$top.soc.cpu.gprf.mem[0][4] ),
    .B1(net1949),
    .B2(\inst$top.soc.cpu.gprf.mem[1][4] ),
    .Y(_06321_));
 sky130_fd_sc_hd__o21ai_0 _25612_ (.A1(_06318_),
    .A2(_06319_),
    .B1(_06321_),
    .Y(_06322_));
 sky130_fd_sc_hd__a21oi_1 _25613_ (.A1(_06322_),
    .A2(net2499),
    .B1(net2592),
    .Y(_06323_));
 sky130_fd_sc_hd__nor2_1 _25614_ (.A(\inst$top.soc.cpu.gprf.mem[23][4] ),
    .B(net2466),
    .Y(_06324_));
 sky130_fd_sc_hd__o21ai_0 _25617_ (.A1(net2657),
    .A2(\inst$top.soc.cpu.gprf.mem[22][4] ),
    .B1(net2621),
    .Y(_06327_));
 sky130_fd_sc_hd__a22oi_1 _25618_ (.A1(net2510),
    .A2(\inst$top.soc.cpu.gprf.mem[20][4] ),
    .B1(net1949),
    .B2(\inst$top.soc.cpu.gprf.mem[21][4] ),
    .Y(_06328_));
 sky130_fd_sc_hd__o21ai_0 _25619_ (.A1(_06324_),
    .A2(_06327_),
    .B1(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__nor2_1 _25620_ (.A(\inst$top.soc.cpu.gprf.mem[19][4] ),
    .B(net2466),
    .Y(_06330_));
 sky130_fd_sc_hd__o21ai_0 _25623_ (.A1(net2657),
    .A2(\inst$top.soc.cpu.gprf.mem[18][4] ),
    .B1(net2623),
    .Y(_06333_));
 sky130_fd_sc_hd__a22oi_1 _25624_ (.A1(net2510),
    .A2(\inst$top.soc.cpu.gprf.mem[16][4] ),
    .B1(net1949),
    .B2(\inst$top.soc.cpu.gprf.mem[17][4] ),
    .Y(_06334_));
 sky130_fd_sc_hd__o21ai_0 _25625_ (.A1(_06330_),
    .A2(_06333_),
    .B1(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__a221oi_1 _25626_ (.A1(_06329_),
    .A2(net1934),
    .B1(net2499),
    .B2(_06335_),
    .C1(net2446),
    .Y(_06336_));
 sky130_fd_sc_hd__nor2_1 _25627_ (.A(\inst$top.soc.cpu.gprf.mem[31][4] ),
    .B(net2466),
    .Y(_06337_));
 sky130_fd_sc_hd__o21ai_0 _25628_ (.A1(net2657),
    .A2(\inst$top.soc.cpu.gprf.mem[30][4] ),
    .B1(net2621),
    .Y(_06338_));
 sky130_fd_sc_hd__a221oi_1 _25629_ (.A1(net2510),
    .A2(\inst$top.soc.cpu.gprf.mem[28][4] ),
    .B1(net1949),
    .B2(\inst$top.soc.cpu.gprf.mem[29][4] ),
    .C1(net2451),
    .Y(_06339_));
 sky130_fd_sc_hd__o21ai_0 _25630_ (.A1(_06337_),
    .A2(_06338_),
    .B1(_06339_),
    .Y(_06340_));
 sky130_fd_sc_hd__nor2_1 _25632_ (.A(\inst$top.soc.cpu.gprf.mem[27][4] ),
    .B(net2466),
    .Y(_06342_));
 sky130_fd_sc_hd__o21ai_0 _25633_ (.A1(net2653),
    .A2(\inst$top.soc.cpu.gprf.mem[26][4] ),
    .B1(net2621),
    .Y(_06343_));
 sky130_fd_sc_hd__a221oi_1 _25634_ (.A1(net2510),
    .A2(\inst$top.soc.cpu.gprf.mem[24][4] ),
    .B1(net1949),
    .B2(\inst$top.soc.cpu.gprf.mem[25][4] ),
    .C1(net2607),
    .Y(_06344_));
 sky130_fd_sc_hd__o21ai_0 _25635_ (.A1(_06342_),
    .A2(_06343_),
    .B1(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand3_1 _25636_ (.A(_06340_),
    .B(_06345_),
    .C(net2600),
    .Y(_06346_));
 sky130_fd_sc_hd__a32oi_1 _25637_ (.A1(_06312_),
    .A2(_06317_),
    .A3(_06323_),
    .B1(_06336_),
    .B2(_06346_),
    .Y(_00026_));
 sky130_fd_sc_hd__nor2_1 _25638_ (.A(\inst$top.soc.cpu.gprf.mem[11][5] ),
    .B(net2479),
    .Y(_06347_));
 sky130_fd_sc_hd__o21ai_0 _25639_ (.A1(net2668),
    .A2(\inst$top.soc.cpu.gprf.mem[10][5] ),
    .B1(net2633),
    .Y(_06348_));
 sky130_fd_sc_hd__a221oi_1 _25640_ (.A1(net2520),
    .A2(\inst$top.soc.cpu.gprf.mem[8][5] ),
    .B1(net1960),
    .B2(\inst$top.soc.cpu.gprf.mem[9][5] ),
    .C1(net2611),
    .Y(_06349_));
 sky130_fd_sc_hd__o21ai_0 _25641_ (.A1(_06347_),
    .A2(_06348_),
    .B1(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__nor2_1 _25642_ (.A(\inst$top.soc.cpu.gprf.mem[15][5] ),
    .B(net2470),
    .Y(_06351_));
 sky130_fd_sc_hd__o21ai_0 _25643_ (.A1(net2666),
    .A2(\inst$top.soc.cpu.gprf.mem[14][5] ),
    .B1(net2633),
    .Y(_06352_));
 sky130_fd_sc_hd__a221oi_1 _25644_ (.A1(net2518),
    .A2(\inst$top.soc.cpu.gprf.mem[12][5] ),
    .B1(net1958),
    .B2(\inst$top.soc.cpu.gprf.mem[13][5] ),
    .C1(net2454),
    .Y(_06353_));
 sky130_fd_sc_hd__o21ai_0 _25645_ (.A1(_06351_),
    .A2(_06352_),
    .B1(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__nand3_1 _25646_ (.A(_06350_),
    .B(_06354_),
    .C(net2601),
    .Y(_06355_));
 sky130_fd_sc_hd__nor2_1 _25647_ (.A(\inst$top.soc.cpu.gprf.mem[7][5] ),
    .B(net2479),
    .Y(_06356_));
 sky130_fd_sc_hd__o21ai_0 _25648_ (.A1(net2666),
    .A2(\inst$top.soc.cpu.gprf.mem[6][5] ),
    .B1(net2633),
    .Y(_06357_));
 sky130_fd_sc_hd__a22oi_1 _25649_ (.A1(net2518),
    .A2(\inst$top.soc.cpu.gprf.mem[4][5] ),
    .B1(net1958),
    .B2(\inst$top.soc.cpu.gprf.mem[5][5] ),
    .Y(_06358_));
 sky130_fd_sc_hd__o21ai_0 _25650_ (.A1(_06356_),
    .A2(_06357_),
    .B1(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__nand2_1 _25651_ (.A(_06359_),
    .B(net1937),
    .Y(_06360_));
 sky130_fd_sc_hd__nor2_1 _25652_ (.A(\inst$top.soc.cpu.gprf.mem[3][5] ),
    .B(net2470),
    .Y(_06361_));
 sky130_fd_sc_hd__o21ai_0 _25653_ (.A1(net2666),
    .A2(\inst$top.soc.cpu.gprf.mem[2][5] ),
    .B1(net2633),
    .Y(_06362_));
 sky130_fd_sc_hd__a22oi_1 _25654_ (.A1(net2518),
    .A2(\inst$top.soc.cpu.gprf.mem[0][5] ),
    .B1(net1958),
    .B2(\inst$top.soc.cpu.gprf.mem[1][5] ),
    .Y(_06363_));
 sky130_fd_sc_hd__o21ai_0 _25655_ (.A1(_06361_),
    .A2(_06362_),
    .B1(_06363_),
    .Y(_06364_));
 sky130_fd_sc_hd__a21oi_1 _25656_ (.A1(_06364_),
    .A2(net2500),
    .B1(net2594),
    .Y(_06365_));
 sky130_fd_sc_hd__nor2_1 _25657_ (.A(\inst$top.soc.cpu.gprf.mem[23][5] ),
    .B(net2481),
    .Y(_06366_));
 sky130_fd_sc_hd__o21ai_0 _25658_ (.A1(net2669),
    .A2(\inst$top.soc.cpu.gprf.mem[22][5] ),
    .B1(net2635),
    .Y(_06367_));
 sky130_fd_sc_hd__a22oi_1 _25659_ (.A1(net2521),
    .A2(\inst$top.soc.cpu.gprf.mem[20][5] ),
    .B1(net1960),
    .B2(\inst$top.soc.cpu.gprf.mem[21][5] ),
    .Y(_06368_));
 sky130_fd_sc_hd__o21ai_0 _25660_ (.A1(_06366_),
    .A2(_06367_),
    .B1(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__nor2_1 _25661_ (.A(\inst$top.soc.cpu.gprf.mem[19][5] ),
    .B(net2472),
    .Y(_06370_));
 sky130_fd_sc_hd__o21ai_0 _25662_ (.A1(net2667),
    .A2(\inst$top.soc.cpu.gprf.mem[18][5] ),
    .B1(net2635),
    .Y(_06371_));
 sky130_fd_sc_hd__a22oi_1 _25663_ (.A1(net2519),
    .A2(\inst$top.soc.cpu.gprf.mem[16][5] ),
    .B1(net1959),
    .B2(\inst$top.soc.cpu.gprf.mem[17][5] ),
    .Y(_06372_));
 sky130_fd_sc_hd__o21ai_0 _25664_ (.A1(_06370_),
    .A2(_06371_),
    .B1(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__a221oi_1 _25665_ (.A1(_06369_),
    .A2(net1937),
    .B1(net2500),
    .B2(_06373_),
    .C1(net2447),
    .Y(_06374_));
 sky130_fd_sc_hd__nor2_1 _25666_ (.A(\inst$top.soc.cpu.gprf.mem[31][5] ),
    .B(net2479),
    .Y(_06375_));
 sky130_fd_sc_hd__o21ai_0 _25667_ (.A1(net2668),
    .A2(\inst$top.soc.cpu.gprf.mem[30][5] ),
    .B1(net2633),
    .Y(_06376_));
 sky130_fd_sc_hd__a221oi_1 _25668_ (.A1(net2520),
    .A2(\inst$top.soc.cpu.gprf.mem[28][5] ),
    .B1(net1960),
    .B2(\inst$top.soc.cpu.gprf.mem[29][5] ),
    .C1(net2456),
    .Y(_06377_));
 sky130_fd_sc_hd__o21ai_0 _25669_ (.A1(_06375_),
    .A2(_06376_),
    .B1(_06377_),
    .Y(_06378_));
 sky130_fd_sc_hd__nor2_1 _25670_ (.A(\inst$top.soc.cpu.gprf.mem[27][5] ),
    .B(net2479),
    .Y(_06379_));
 sky130_fd_sc_hd__o21ai_0 _25671_ (.A1(net2668),
    .A2(\inst$top.soc.cpu.gprf.mem[26][5] ),
    .B1(net2633),
    .Y(_06380_));
 sky130_fd_sc_hd__a221oi_1 _25672_ (.A1(net2520),
    .A2(\inst$top.soc.cpu.gprf.mem[24][5] ),
    .B1(net1960),
    .B2(\inst$top.soc.cpu.gprf.mem[25][5] ),
    .C1(net2611),
    .Y(_06381_));
 sky130_fd_sc_hd__o21ai_0 _25673_ (.A1(_06379_),
    .A2(_06380_),
    .B1(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__nand3_1 _25674_ (.A(_06378_),
    .B(_06382_),
    .C(net2601),
    .Y(_06383_));
 sky130_fd_sc_hd__a32oi_1 _25675_ (.A1(_06355_),
    .A2(_06360_),
    .A3(_06365_),
    .B1(_06374_),
    .B2(_06383_),
    .Y(_00027_));
 sky130_fd_sc_hd__nor2_1 _25676_ (.A(\inst$top.soc.cpu.gprf.mem[15][6] ),
    .B(net2472),
    .Y(_06384_));
 sky130_fd_sc_hd__o21ai_0 _25677_ (.A1(net2666),
    .A2(\inst$top.soc.cpu.gprf.mem[14][6] ),
    .B1(net2626),
    .Y(_06385_));
 sky130_fd_sc_hd__a221oi_1 _25678_ (.A1(net2518),
    .A2(\inst$top.soc.cpu.gprf.mem[12][6] ),
    .B1(net1958),
    .B2(\inst$top.soc.cpu.gprf.mem[13][6] ),
    .C1(net2454),
    .Y(_06386_));
 sky130_fd_sc_hd__o21ai_0 _25679_ (.A1(_06384_),
    .A2(_06385_),
    .B1(_06386_),
    .Y(_06387_));
 sky130_fd_sc_hd__nor2_1 _25680_ (.A(\inst$top.soc.cpu.gprf.mem[11][6] ),
    .B(net2470),
    .Y(_06388_));
 sky130_fd_sc_hd__o21ai_0 _25681_ (.A1(net2666),
    .A2(\inst$top.soc.cpu.gprf.mem[10][6] ),
    .B1(net2624),
    .Y(_06389_));
 sky130_fd_sc_hd__a221oi_1 _25683_ (.A1(net2518),
    .A2(\inst$top.soc.cpu.gprf.mem[8][6] ),
    .B1(net1958),
    .B2(\inst$top.soc.cpu.gprf.mem[9][6] ),
    .C1(net2610),
    .Y(_06391_));
 sky130_fd_sc_hd__o21ai_0 _25684_ (.A1(_06388_),
    .A2(_06389_),
    .B1(_06391_),
    .Y(_06392_));
 sky130_fd_sc_hd__nand3_1 _25685_ (.A(_06387_),
    .B(_06392_),
    .C(net2598),
    .Y(_06393_));
 sky130_fd_sc_hd__nor2_1 _25686_ (.A(\inst$top.soc.cpu.gprf.mem[7][6] ),
    .B(net2470),
    .Y(_06394_));
 sky130_fd_sc_hd__o21ai_0 _25687_ (.A1(net2666),
    .A2(\inst$top.soc.cpu.gprf.mem[6][6] ),
    .B1(net2624),
    .Y(_06395_));
 sky130_fd_sc_hd__a22oi_1 _25688_ (.A1(net2518),
    .A2(\inst$top.soc.cpu.gprf.mem[4][6] ),
    .B1(net1958),
    .B2(\inst$top.soc.cpu.gprf.mem[5][6] ),
    .Y(_06396_));
 sky130_fd_sc_hd__o21ai_0 _25689_ (.A1(_06394_),
    .A2(_06395_),
    .B1(_06396_),
    .Y(_06397_));
 sky130_fd_sc_hd__nand2_1 _25690_ (.A(_06397_),
    .B(net1935),
    .Y(_06398_));
 sky130_fd_sc_hd__nor2_1 _25691_ (.A(\inst$top.soc.cpu.gprf.mem[3][6] ),
    .B(net2470),
    .Y(_06399_));
 sky130_fd_sc_hd__o21ai_0 _25692_ (.A1(net2659),
    .A2(\inst$top.soc.cpu.gprf.mem[2][6] ),
    .B1(net2624),
    .Y(_06400_));
 sky130_fd_sc_hd__a22oi_1 _25694_ (.A1(net2518),
    .A2(\inst$top.soc.cpu.gprf.mem[0][6] ),
    .B1(net1958),
    .B2(\inst$top.soc.cpu.gprf.mem[1][6] ),
    .Y(_06402_));
 sky130_fd_sc_hd__o21ai_0 _25695_ (.A1(_06399_),
    .A2(_06400_),
    .B1(_06402_),
    .Y(_06403_));
 sky130_fd_sc_hd__a21oi_1 _25696_ (.A1(_06403_),
    .A2(net2497),
    .B1(net2594),
    .Y(_06404_));
 sky130_fd_sc_hd__nor2_1 _25697_ (.A(\inst$top.soc.cpu.gprf.mem[23][6] ),
    .B(net2472),
    .Y(_06405_));
 sky130_fd_sc_hd__o21ai_0 _25698_ (.A1(net2666),
    .A2(\inst$top.soc.cpu.gprf.mem[22][6] ),
    .B1(net2626),
    .Y(_06406_));
 sky130_fd_sc_hd__a22oi_1 _25701_ (.A1(net2518),
    .A2(\inst$top.soc.cpu.gprf.mem[20][6] ),
    .B1(net1958),
    .B2(\inst$top.soc.cpu.gprf.mem[21][6] ),
    .Y(_06409_));
 sky130_fd_sc_hd__o21ai_0 _25702_ (.A1(_06405_),
    .A2(_06406_),
    .B1(_06409_),
    .Y(_06410_));
 sky130_fd_sc_hd__nor2_1 _25703_ (.A(\inst$top.soc.cpu.gprf.mem[19][6] ),
    .B(net2472),
    .Y(_06411_));
 sky130_fd_sc_hd__o21ai_0 _25704_ (.A1(net2666),
    .A2(\inst$top.soc.cpu.gprf.mem[18][6] ),
    .B1(net2626),
    .Y(_06412_));
 sky130_fd_sc_hd__a22oi_1 _25707_ (.A1(net2519),
    .A2(\inst$top.soc.cpu.gprf.mem[16][6] ),
    .B1(net1959),
    .B2(\inst$top.soc.cpu.gprf.mem[17][6] ),
    .Y(_06415_));
 sky130_fd_sc_hd__o21ai_0 _25708_ (.A1(_06411_),
    .A2(_06412_),
    .B1(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__a221oi_1 _25709_ (.A1(_06410_),
    .A2(net1935),
    .B1(net2497),
    .B2(_06416_),
    .C1(net2449),
    .Y(_06417_));
 sky130_fd_sc_hd__nor2_1 _25710_ (.A(\inst$top.soc.cpu.gprf.mem[31][6] ),
    .B(net2470),
    .Y(_06418_));
 sky130_fd_sc_hd__o21ai_0 _25711_ (.A1(net2666),
    .A2(\inst$top.soc.cpu.gprf.mem[30][6] ),
    .B1(net2624),
    .Y(_06419_));
 sky130_fd_sc_hd__a221oi_1 _25712_ (.A1(net2518),
    .A2(\inst$top.soc.cpu.gprf.mem[28][6] ),
    .B1(net1958),
    .B2(\inst$top.soc.cpu.gprf.mem[29][6] ),
    .C1(net2454),
    .Y(_06420_));
 sky130_fd_sc_hd__o21ai_0 _25713_ (.A1(_06418_),
    .A2(_06419_),
    .B1(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__nor2_1 _25714_ (.A(\inst$top.soc.cpu.gprf.mem[27][6] ),
    .B(net2472),
    .Y(_06422_));
 sky130_fd_sc_hd__o21ai_0 _25715_ (.A1(net2666),
    .A2(\inst$top.soc.cpu.gprf.mem[26][6] ),
    .B1(net2626),
    .Y(_06423_));
 sky130_fd_sc_hd__a221oi_1 _25716_ (.A1(net2518),
    .A2(\inst$top.soc.cpu.gprf.mem[24][6] ),
    .B1(net1958),
    .B2(\inst$top.soc.cpu.gprf.mem[25][6] ),
    .C1(net2610),
    .Y(_06424_));
 sky130_fd_sc_hd__o21ai_0 _25717_ (.A1(_06422_),
    .A2(_06423_),
    .B1(_06424_),
    .Y(_06425_));
 sky130_fd_sc_hd__nand3_1 _25718_ (.A(_06421_),
    .B(_06425_),
    .C(net2598),
    .Y(_06426_));
 sky130_fd_sc_hd__a32oi_1 _25719_ (.A1(_06393_),
    .A2(_06398_),
    .A3(_06404_),
    .B1(_06417_),
    .B2(_06426_),
    .Y(_00028_));
 sky130_fd_sc_hd__nor2_1 _25720_ (.A(\inst$top.soc.cpu.gprf.mem[15][7] ),
    .B(net2486),
    .Y(_06427_));
 sky130_fd_sc_hd__o21ai_0 _25721_ (.A1(net2677),
    .A2(\inst$top.soc.cpu.gprf.mem[14][7] ),
    .B1(net2638),
    .Y(_06428_));
 sky130_fd_sc_hd__a221oi_1 _25722_ (.A1(net2529),
    .A2(\inst$top.soc.cpu.gprf.mem[12][7] ),
    .B1(net1969),
    .B2(\inst$top.soc.cpu.gprf.mem[13][7] ),
    .C1(net2457),
    .Y(_06429_));
 sky130_fd_sc_hd__o21ai_0 _25723_ (.A1(_06427_),
    .A2(_06428_),
    .B1(_06429_),
    .Y(_06430_));
 sky130_fd_sc_hd__nor2_1 _25724_ (.A(\inst$top.soc.cpu.gprf.mem[11][7] ),
    .B(net2483),
    .Y(_06431_));
 sky130_fd_sc_hd__o21ai_0 _25725_ (.A1(net2677),
    .A2(\inst$top.soc.cpu.gprf.mem[10][7] ),
    .B1(net2637),
    .Y(_06432_));
 sky130_fd_sc_hd__a221oi_1 _25727_ (.A1(net2529),
    .A2(\inst$top.soc.cpu.gprf.mem[8][7] ),
    .B1(net1969),
    .B2(\inst$top.soc.cpu.gprf.mem[9][7] ),
    .C1(net2611),
    .Y(_06434_));
 sky130_fd_sc_hd__o21ai_0 _25728_ (.A1(_06431_),
    .A2(_06432_),
    .B1(_06434_),
    .Y(_06435_));
 sky130_fd_sc_hd__nand3_1 _25729_ (.A(_06430_),
    .B(_06435_),
    .C(net2603),
    .Y(_06436_));
 sky130_fd_sc_hd__nor2_1 _25730_ (.A(\inst$top.soc.cpu.gprf.mem[3][7] ),
    .B(net2483),
    .Y(_06437_));
 sky130_fd_sc_hd__o21ai_0 _25731_ (.A1(net2677),
    .A2(\inst$top.soc.cpu.gprf.mem[2][7] ),
    .B1(net2637),
    .Y(_06438_));
 sky130_fd_sc_hd__a22oi_1 _25732_ (.A1(net2529),
    .A2(\inst$top.soc.cpu.gprf.mem[0][7] ),
    .B1(net1969),
    .B2(\inst$top.soc.cpu.gprf.mem[1][7] ),
    .Y(_06439_));
 sky130_fd_sc_hd__o21ai_0 _25733_ (.A1(_06437_),
    .A2(_06438_),
    .B1(_06439_),
    .Y(_06440_));
 sky130_fd_sc_hd__nand2_1 _25734_ (.A(_06440_),
    .B(net2501),
    .Y(_06441_));
 sky130_fd_sc_hd__nor2_1 _25735_ (.A(\inst$top.soc.cpu.gprf.mem[7][7] ),
    .B(net2483),
    .Y(_06442_));
 sky130_fd_sc_hd__o21ai_0 _25736_ (.A1(net2677),
    .A2(\inst$top.soc.cpu.gprf.mem[6][7] ),
    .B1(net2637),
    .Y(_06443_));
 sky130_fd_sc_hd__a22oi_1 _25737_ (.A1(net2529),
    .A2(\inst$top.soc.cpu.gprf.mem[4][7] ),
    .B1(net1969),
    .B2(\inst$top.soc.cpu.gprf.mem[5][7] ),
    .Y(_06444_));
 sky130_fd_sc_hd__o21ai_0 _25738_ (.A1(_06442_),
    .A2(_06443_),
    .B1(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__a21oi_1 _25739_ (.A1(_06445_),
    .A2(net1938),
    .B1(net2593),
    .Y(_06446_));
 sky130_fd_sc_hd__nor2_1 _25740_ (.A(\inst$top.soc.cpu.gprf.mem[19][7] ),
    .B(net2483),
    .Y(_06447_));
 sky130_fd_sc_hd__o21ai_0 _25741_ (.A1(net2677),
    .A2(\inst$top.soc.cpu.gprf.mem[18][7] ),
    .B1(net2638),
    .Y(_06448_));
 sky130_fd_sc_hd__a22oi_1 _25742_ (.A1(net2530),
    .A2(\inst$top.soc.cpu.gprf.mem[16][7] ),
    .B1(net1969),
    .B2(\inst$top.soc.cpu.gprf.mem[17][7] ),
    .Y(_06449_));
 sky130_fd_sc_hd__o21ai_0 _25743_ (.A1(_06447_),
    .A2(_06448_),
    .B1(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__nor2_1 _25746_ (.A(\inst$top.soc.cpu.gprf.mem[23][7] ),
    .B(net2483),
    .Y(_06453_));
 sky130_fd_sc_hd__o21ai_0 _25747_ (.A1(net2678),
    .A2(\inst$top.soc.cpu.gprf.mem[22][7] ),
    .B1(net2638),
    .Y(_06454_));
 sky130_fd_sc_hd__a22oi_1 _25748_ (.A1(net2530),
    .A2(\inst$top.soc.cpu.gprf.mem[20][7] ),
    .B1(net1970),
    .B2(\inst$top.soc.cpu.gprf.mem[21][7] ),
    .Y(_06455_));
 sky130_fd_sc_hd__o21ai_0 _25749_ (.A1(_06453_),
    .A2(_06454_),
    .B1(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__a221oi_1 _25750_ (.A1(_06450_),
    .A2(net2501),
    .B1(net1938),
    .B2(_06456_),
    .C1(net2448),
    .Y(_06457_));
 sky130_fd_sc_hd__nor2_1 _25751_ (.A(\inst$top.soc.cpu.gprf.mem[31][7] ),
    .B(net2483),
    .Y(_06458_));
 sky130_fd_sc_hd__o21ai_0 _25752_ (.A1(net2677),
    .A2(\inst$top.soc.cpu.gprf.mem[30][7] ),
    .B1(net2637),
    .Y(_06459_));
 sky130_fd_sc_hd__a221oi_1 _25753_ (.A1(net2529),
    .A2(\inst$top.soc.cpu.gprf.mem[28][7] ),
    .B1(net1969),
    .B2(\inst$top.soc.cpu.gprf.mem[29][7] ),
    .C1(net2457),
    .Y(_06460_));
 sky130_fd_sc_hd__o21ai_0 _25754_ (.A1(_06458_),
    .A2(_06459_),
    .B1(_06460_),
    .Y(_06461_));
 sky130_fd_sc_hd__nor2_1 _25755_ (.A(\inst$top.soc.cpu.gprf.mem[27][7] ),
    .B(net2486),
    .Y(_06462_));
 sky130_fd_sc_hd__o21ai_0 _25756_ (.A1(net2677),
    .A2(\inst$top.soc.cpu.gprf.mem[26][7] ),
    .B1(net2638),
    .Y(_06463_));
 sky130_fd_sc_hd__a221oi_1 _25757_ (.A1(net2529),
    .A2(\inst$top.soc.cpu.gprf.mem[24][7] ),
    .B1(net1969),
    .B2(\inst$top.soc.cpu.gprf.mem[25][7] ),
    .C1(net2612),
    .Y(_06464_));
 sky130_fd_sc_hd__o21ai_0 _25758_ (.A1(_06462_),
    .A2(_06463_),
    .B1(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__nand3_1 _25759_ (.A(_06461_),
    .B(_06465_),
    .C(net2603),
    .Y(_06466_));
 sky130_fd_sc_hd__a32oi_1 _25760_ (.A1(_06436_),
    .A2(_06441_),
    .A3(_06446_),
    .B1(_06457_),
    .B2(_06466_),
    .Y(_00029_));
 sky130_fd_sc_hd__nor2_1 _25761_ (.A(\inst$top.soc.cpu.gprf.mem[11][8] ),
    .B(net2467),
    .Y(_06467_));
 sky130_fd_sc_hd__o21ai_0 _25762_ (.A1(net2657),
    .A2(\inst$top.soc.cpu.gprf.mem[10][8] ),
    .B1(net2621),
    .Y(_06468_));
 sky130_fd_sc_hd__a221oi_1 _25763_ (.A1(net2512),
    .A2(\inst$top.soc.cpu.gprf.mem[8][8] ),
    .B1(net1951),
    .B2(\inst$top.soc.cpu.gprf.mem[9][8] ),
    .C1(net2610),
    .Y(_06469_));
 sky130_fd_sc_hd__o21ai_0 _25764_ (.A1(_06467_),
    .A2(_06468_),
    .B1(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__nor2_1 _25765_ (.A(\inst$top.soc.cpu.gprf.mem[15][8] ),
    .B(net2466),
    .Y(_06471_));
 sky130_fd_sc_hd__o21ai_0 _25768_ (.A1(net2657),
    .A2(\inst$top.soc.cpu.gprf.mem[14][8] ),
    .B1(net2623),
    .Y(_06474_));
 sky130_fd_sc_hd__a221oi_1 _25769_ (.A1(net2511),
    .A2(\inst$top.soc.cpu.gprf.mem[12][8] ),
    .B1(net1950),
    .B2(\inst$top.soc.cpu.gprf.mem[13][8] ),
    .C1(net2453),
    .Y(_06475_));
 sky130_fd_sc_hd__o21ai_0 _25770_ (.A1(_06471_),
    .A2(_06474_),
    .B1(_06475_),
    .Y(_06476_));
 sky130_fd_sc_hd__nand3_1 _25771_ (.A(_06470_),
    .B(_06476_),
    .C(net2598),
    .Y(_06477_));
 sky130_fd_sc_hd__nor2_1 _25772_ (.A(\inst$top.soc.cpu.gprf.mem[7][8] ),
    .B(net2468),
    .Y(_06478_));
 sky130_fd_sc_hd__o21ai_0 _25773_ (.A1(net2658),
    .A2(\inst$top.soc.cpu.gprf.mem[6][8] ),
    .B1(net2622),
    .Y(_06479_));
 sky130_fd_sc_hd__a22oi_1 _25774_ (.A1(net2511),
    .A2(\inst$top.soc.cpu.gprf.mem[4][8] ),
    .B1(net1950),
    .B2(\inst$top.soc.cpu.gprf.mem[5][8] ),
    .Y(_06480_));
 sky130_fd_sc_hd__o21ai_0 _25775_ (.A1(_06478_),
    .A2(_06479_),
    .B1(_06480_),
    .Y(_06481_));
 sky130_fd_sc_hd__nand2_1 _25776_ (.A(_06481_),
    .B(net1934),
    .Y(_06482_));
 sky130_fd_sc_hd__nor2_1 _25777_ (.A(\inst$top.soc.cpu.gprf.mem[3][8] ),
    .B(net2469),
    .Y(_06483_));
 sky130_fd_sc_hd__o21ai_0 _25778_ (.A1(net2658),
    .A2(\inst$top.soc.cpu.gprf.mem[2][8] ),
    .B1(net2622),
    .Y(_06484_));
 sky130_fd_sc_hd__a22oi_1 _25779_ (.A1(net2513),
    .A2(\inst$top.soc.cpu.gprf.mem[0][8] ),
    .B1(net1952),
    .B2(\inst$top.soc.cpu.gprf.mem[1][8] ),
    .Y(_06485_));
 sky130_fd_sc_hd__o21ai_0 _25780_ (.A1(_06483_),
    .A2(_06484_),
    .B1(_06485_),
    .Y(_06486_));
 sky130_fd_sc_hd__a21oi_1 _25782_ (.A1(_06486_),
    .A2(net2499),
    .B1(net2596),
    .Y(_06488_));
 sky130_fd_sc_hd__nor2_1 _25783_ (.A(\inst$top.soc.cpu.gprf.mem[19][8] ),
    .B(net2469),
    .Y(_06489_));
 sky130_fd_sc_hd__o21ai_0 _25784_ (.A1(net2660),
    .A2(\inst$top.soc.cpu.gprf.mem[18][8] ),
    .B1(net2625),
    .Y(_06490_));
 sky130_fd_sc_hd__a22oi_1 _25785_ (.A1(net2513),
    .A2(\inst$top.soc.cpu.gprf.mem[16][8] ),
    .B1(net1952),
    .B2(\inst$top.soc.cpu.gprf.mem[17][8] ),
    .Y(_06491_));
 sky130_fd_sc_hd__o21ai_0 _25786_ (.A1(_06489_),
    .A2(_06490_),
    .B1(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__nor2_1 _25787_ (.A(\inst$top.soc.cpu.gprf.mem[23][8] ),
    .B(net2469),
    .Y(_06493_));
 sky130_fd_sc_hd__o21ai_0 _25788_ (.A1(net2660),
    .A2(\inst$top.soc.cpu.gprf.mem[22][8] ),
    .B1(net2625),
    .Y(_06494_));
 sky130_fd_sc_hd__a22oi_1 _25789_ (.A1(net2513),
    .A2(\inst$top.soc.cpu.gprf.mem[20][8] ),
    .B1(net1952),
    .B2(\inst$top.soc.cpu.gprf.mem[21][8] ),
    .Y(_06495_));
 sky130_fd_sc_hd__o21ai_0 _25790_ (.A1(_06493_),
    .A2(_06494_),
    .B1(_06495_),
    .Y(_06496_));
 sky130_fd_sc_hd__a221oi_1 _25791_ (.A1(_06492_),
    .A2(net2497),
    .B1(net1935),
    .B2(_06496_),
    .C1(net2446),
    .Y(_06497_));
 sky130_fd_sc_hd__nor2_1 _25792_ (.A(\inst$top.soc.cpu.gprf.mem[31][8] ),
    .B(net2468),
    .Y(_06498_));
 sky130_fd_sc_hd__o21ai_0 _25793_ (.A1(net2658),
    .A2(\inst$top.soc.cpu.gprf.mem[30][8] ),
    .B1(net2622),
    .Y(_06499_));
 sky130_fd_sc_hd__a221oi_1 _25794_ (.A1(net2511),
    .A2(\inst$top.soc.cpu.gprf.mem[28][8] ),
    .B1(net1950),
    .B2(\inst$top.soc.cpu.gprf.mem[29][8] ),
    .C1(net2453),
    .Y(_06500_));
 sky130_fd_sc_hd__o21ai_0 _25795_ (.A1(_06498_),
    .A2(_06499_),
    .B1(_06500_),
    .Y(_06501_));
 sky130_fd_sc_hd__nor2_1 _25796_ (.A(\inst$top.soc.cpu.gprf.mem[27][8] ),
    .B(net2469),
    .Y(_06502_));
 sky130_fd_sc_hd__o21ai_0 _25797_ (.A1(net2658),
    .A2(\inst$top.soc.cpu.gprf.mem[26][8] ),
    .B1(net2622),
    .Y(_06503_));
 sky130_fd_sc_hd__a221oi_1 _25798_ (.A1(net2513),
    .A2(\inst$top.soc.cpu.gprf.mem[24][8] ),
    .B1(net1952),
    .B2(\inst$top.soc.cpu.gprf.mem[25][8] ),
    .C1(net2610),
    .Y(_06504_));
 sky130_fd_sc_hd__o21ai_0 _25799_ (.A1(_06502_),
    .A2(_06503_),
    .B1(_06504_),
    .Y(_06505_));
 sky130_fd_sc_hd__nand3_1 _25800_ (.A(_06501_),
    .B(_06505_),
    .C(net2598),
    .Y(_06506_));
 sky130_fd_sc_hd__a32oi_1 _25801_ (.A1(_06477_),
    .A2(_06482_),
    .A3(_06488_),
    .B1(_06497_),
    .B2(_06506_),
    .Y(_00030_));
 sky130_fd_sc_hd__nor2_1 _25802_ (.A(\inst$top.soc.cpu.gprf.mem[31][9] ),
    .B(net2472),
    .Y(_06507_));
 sky130_fd_sc_hd__o21ai_0 _25803_ (.A1(net2667),
    .A2(\inst$top.soc.cpu.gprf.mem[30][9] ),
    .B1(net2626),
    .Y(_06508_));
 sky130_fd_sc_hd__a221oi_1 _25805_ (.A1(net2519),
    .A2(\inst$top.soc.cpu.gprf.mem[28][9] ),
    .B1(net1959),
    .B2(\inst$top.soc.cpu.gprf.mem[29][9] ),
    .C1(net2454),
    .Y(_06510_));
 sky130_fd_sc_hd__o21ai_0 _25806_ (.A1(_06507_),
    .A2(_06508_),
    .B1(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__nor2_1 _25807_ (.A(\inst$top.soc.cpu.gprf.mem[27][9] ),
    .B(net2471),
    .Y(_06512_));
 sky130_fd_sc_hd__o21ai_0 _25808_ (.A1(net2667),
    .A2(\inst$top.soc.cpu.gprf.mem[26][9] ),
    .B1(net2635),
    .Y(_06513_));
 sky130_fd_sc_hd__a221oi_1 _25810_ (.A1(net2521),
    .A2(\inst$top.soc.cpu.gprf.mem[24][9] ),
    .B1(net1961),
    .B2(\inst$top.soc.cpu.gprf.mem[25][9] ),
    .C1(net2610),
    .Y(_06515_));
 sky130_fd_sc_hd__o21ai_0 _25811_ (.A1(_06512_),
    .A2(_06513_),
    .B1(_06515_),
    .Y(_06516_));
 sky130_fd_sc_hd__nand3_1 _25812_ (.A(_06511_),
    .B(_06516_),
    .C(net2601),
    .Y(_06517_));
 sky130_fd_sc_hd__nor2_1 _25813_ (.A(\inst$top.soc.cpu.gprf.mem[19][9] ),
    .B(net2477),
    .Y(_06518_));
 sky130_fd_sc_hd__o21ai_0 _25814_ (.A1(net2667),
    .A2(\inst$top.soc.cpu.gprf.mem[18][9] ),
    .B1(net2631),
    .Y(_06519_));
 sky130_fd_sc_hd__a22oi_1 _25816_ (.A1(net2523),
    .A2(\inst$top.soc.cpu.gprf.mem[16][9] ),
    .B1(net1963),
    .B2(\inst$top.soc.cpu.gprf.mem[17][9] ),
    .Y(_06521_));
 sky130_fd_sc_hd__o21ai_0 _25817_ (.A1(_06518_),
    .A2(_06519_),
    .B1(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__a21oi_1 _25819_ (.A1(_06522_),
    .A2(net2497),
    .B1(net2446),
    .Y(_06524_));
 sky130_fd_sc_hd__nor2_1 _25821_ (.A(\inst$top.soc.cpu.gprf.mem[23][9] ),
    .B(net2481),
    .Y(_06526_));
 sky130_fd_sc_hd__o21ai_0 _25824_ (.A1(net2669),
    .A2(\inst$top.soc.cpu.gprf.mem[22][9] ),
    .B1(net2635),
    .Y(_06529_));
 sky130_fd_sc_hd__a22oi_1 _25827_ (.A1(net2521),
    .A2(\inst$top.soc.cpu.gprf.mem[20][9] ),
    .B1(net1961),
    .B2(\inst$top.soc.cpu.gprf.mem[21][9] ),
    .Y(_06532_));
 sky130_fd_sc_hd__o21ai_0 _25828_ (.A1(_06526_),
    .A2(_06529_),
    .B1(_06532_),
    .Y(_06533_));
 sky130_fd_sc_hd__nand2_1 _25829_ (.A(_06533_),
    .B(net1937),
    .Y(_06534_));
 sky130_fd_sc_hd__nor2_1 _25830_ (.A(\inst$top.soc.cpu.gprf.mem[3][9] ),
    .B(net2472),
    .Y(_06535_));
 sky130_fd_sc_hd__o21ai_0 _25831_ (.A1(net2667),
    .A2(\inst$top.soc.cpu.gprf.mem[2][9] ),
    .B1(net2626),
    .Y(_06536_));
 sky130_fd_sc_hd__a22oi_1 _25832_ (.A1(net2519),
    .A2(\inst$top.soc.cpu.gprf.mem[0][9] ),
    .B1(net1959),
    .B2(\inst$top.soc.cpu.gprf.mem[1][9] ),
    .Y(_06537_));
 sky130_fd_sc_hd__o21ai_0 _25833_ (.A1(_06535_),
    .A2(_06536_),
    .B1(_06537_),
    .Y(_06538_));
 sky130_fd_sc_hd__nor2_1 _25834_ (.A(\inst$top.soc.cpu.gprf.mem[7][9] ),
    .B(net2472),
    .Y(_06539_));
 sky130_fd_sc_hd__o21ai_0 _25835_ (.A1(net2667),
    .A2(\inst$top.soc.cpu.gprf.mem[6][9] ),
    .B1(net2626),
    .Y(_06540_));
 sky130_fd_sc_hd__a22oi_1 _25836_ (.A1(net2519),
    .A2(\inst$top.soc.cpu.gprf.mem[4][9] ),
    .B1(net1959),
    .B2(\inst$top.soc.cpu.gprf.mem[5][9] ),
    .Y(_06541_));
 sky130_fd_sc_hd__o21ai_0 _25837_ (.A1(_06539_),
    .A2(_06540_),
    .B1(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__a221oi_1 _25838_ (.A1(_06538_),
    .A2(net2497),
    .B1(net1935),
    .B2(_06542_),
    .C1(net2594),
    .Y(_06543_));
 sky130_fd_sc_hd__nor2_1 _25839_ (.A(\inst$top.soc.cpu.gprf.mem[15][9] ),
    .B(net2481),
    .Y(_06544_));
 sky130_fd_sc_hd__o21ai_0 _25840_ (.A1(net2669),
    .A2(\inst$top.soc.cpu.gprf.mem[14][9] ),
    .B1(net2635),
    .Y(_06545_));
 sky130_fd_sc_hd__a221oi_1 _25841_ (.A1(net2521),
    .A2(\inst$top.soc.cpu.gprf.mem[12][9] ),
    .B1(net1961),
    .B2(\inst$top.soc.cpu.gprf.mem[13][9] ),
    .C1(net2456),
    .Y(_06546_));
 sky130_fd_sc_hd__o21ai_0 _25842_ (.A1(_06544_),
    .A2(_06545_),
    .B1(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__nor2_1 _25843_ (.A(\inst$top.soc.cpu.gprf.mem[11][9] ),
    .B(net2481),
    .Y(_06548_));
 sky130_fd_sc_hd__o21ai_0 _25844_ (.A1(net2669),
    .A2(\inst$top.soc.cpu.gprf.mem[10][9] ),
    .B1(net2635),
    .Y(_06549_));
 sky130_fd_sc_hd__a221oi_1 _25845_ (.A1(net2521),
    .A2(\inst$top.soc.cpu.gprf.mem[8][9] ),
    .B1(net1961),
    .B2(\inst$top.soc.cpu.gprf.mem[9][9] ),
    .C1(net2611),
    .Y(_06550_));
 sky130_fd_sc_hd__o21ai_0 _25846_ (.A1(_06548_),
    .A2(_06549_),
    .B1(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__nand3_1 _25847_ (.A(_06547_),
    .B(_06551_),
    .C(net2601),
    .Y(_06552_));
 sky130_fd_sc_hd__a32oi_1 _25848_ (.A1(_06517_),
    .A2(_06524_),
    .A3(_06534_),
    .B1(_06543_),
    .B2(_06552_),
    .Y(_00031_));
 sky130_fd_sc_hd__nor2_1 _25849_ (.A(\inst$top.soc.cpu.gprf.mem[11][10] ),
    .B(net2477),
    .Y(_06553_));
 sky130_fd_sc_hd__o21ai_0 _25850_ (.A1(net2671),
    .A2(\inst$top.soc.cpu.gprf.mem[10][10] ),
    .B1(net2631),
    .Y(_06554_));
 sky130_fd_sc_hd__a221oi_1 _25851_ (.A1(net2523),
    .A2(\inst$top.soc.cpu.gprf.mem[8][10] ),
    .B1(net1963),
    .B2(\inst$top.soc.cpu.gprf.mem[9][10] ),
    .C1(net2609),
    .Y(_06555_));
 sky130_fd_sc_hd__o21ai_0 _25852_ (.A1(_06553_),
    .A2(_06554_),
    .B1(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__nor2_1 _25854_ (.A(\inst$top.soc.cpu.gprf.mem[15][10] ),
    .B(net2477),
    .Y(_06558_));
 sky130_fd_sc_hd__o21ai_0 _25855_ (.A1(net2671),
    .A2(\inst$top.soc.cpu.gprf.mem[14][10] ),
    .B1(net2631),
    .Y(_06559_));
 sky130_fd_sc_hd__a221oi_1 _25856_ (.A1(net2523),
    .A2(\inst$top.soc.cpu.gprf.mem[12][10] ),
    .B1(net1963),
    .B2(\inst$top.soc.cpu.gprf.mem[13][10] ),
    .C1(net2454),
    .Y(_06560_));
 sky130_fd_sc_hd__o21ai_0 _25857_ (.A1(_06558_),
    .A2(_06559_),
    .B1(_06560_),
    .Y(_06561_));
 sky130_fd_sc_hd__nand3_1 _25859_ (.A(_06556_),
    .B(_06561_),
    .C(net2602),
    .Y(_06563_));
 sky130_fd_sc_hd__nor2_1 _25860_ (.A(\inst$top.soc.cpu.gprf.mem[7][10] ),
    .B(net2477),
    .Y(_06564_));
 sky130_fd_sc_hd__o21ai_0 _25861_ (.A1(net2662),
    .A2(\inst$top.soc.cpu.gprf.mem[6][10] ),
    .B1(net2631),
    .Y(_06565_));
 sky130_fd_sc_hd__a22oi_1 _25862_ (.A1(net2523),
    .A2(\inst$top.soc.cpu.gprf.mem[4][10] ),
    .B1(net1963),
    .B2(\inst$top.soc.cpu.gprf.mem[5][10] ),
    .Y(_06566_));
 sky130_fd_sc_hd__o21ai_0 _25863_ (.A1(_06564_),
    .A2(_06565_),
    .B1(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__nand2_1 _25864_ (.A(_06567_),
    .B(net1935),
    .Y(_06568_));
 sky130_fd_sc_hd__nor2_1 _25865_ (.A(\inst$top.soc.cpu.gprf.mem[3][10] ),
    .B(net2477),
    .Y(_06569_));
 sky130_fd_sc_hd__o21ai_0 _25866_ (.A1(net2671),
    .A2(\inst$top.soc.cpu.gprf.mem[2][10] ),
    .B1(net2631),
    .Y(_06570_));
 sky130_fd_sc_hd__a22oi_1 _25867_ (.A1(net2523),
    .A2(\inst$top.soc.cpu.gprf.mem[0][10] ),
    .B1(net1963),
    .B2(\inst$top.soc.cpu.gprf.mem[1][10] ),
    .Y(_06571_));
 sky130_fd_sc_hd__o21ai_0 _25868_ (.A1(_06569_),
    .A2(_06570_),
    .B1(_06571_),
    .Y(_06572_));
 sky130_fd_sc_hd__a21oi_1 _25869_ (.A1(_06572_),
    .A2(net2497),
    .B1(net2594),
    .Y(_06573_));
 sky130_fd_sc_hd__nor2_1 _25870_ (.A(\inst$top.soc.cpu.gprf.mem[19][10] ),
    .B(net2477),
    .Y(_06574_));
 sky130_fd_sc_hd__o21ai_0 _25871_ (.A1(net2662),
    .A2(\inst$top.soc.cpu.gprf.mem[18][10] ),
    .B1(net2631),
    .Y(_06575_));
 sky130_fd_sc_hd__a22oi_1 _25872_ (.A1(net2515),
    .A2(\inst$top.soc.cpu.gprf.mem[16][10] ),
    .B1(net1954),
    .B2(\inst$top.soc.cpu.gprf.mem[17][10] ),
    .Y(_06576_));
 sky130_fd_sc_hd__o21ai_0 _25873_ (.A1(_06574_),
    .A2(_06575_),
    .B1(_06576_),
    .Y(_06577_));
 sky130_fd_sc_hd__nor2_1 _25874_ (.A(\inst$top.soc.cpu.gprf.mem[23][10] ),
    .B(net2477),
    .Y(_06578_));
 sky130_fd_sc_hd__o21ai_0 _25875_ (.A1(net2662),
    .A2(\inst$top.soc.cpu.gprf.mem[22][10] ),
    .B1(net2631),
    .Y(_06579_));
 sky130_fd_sc_hd__a22oi_1 _25876_ (.A1(net2515),
    .A2(\inst$top.soc.cpu.gprf.mem[20][10] ),
    .B1(net1954),
    .B2(\inst$top.soc.cpu.gprf.mem[21][10] ),
    .Y(_06580_));
 sky130_fd_sc_hd__o21ai_0 _25877_ (.A1(_06578_),
    .A2(_06579_),
    .B1(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__a221oi_1 _25878_ (.A1(_06577_),
    .A2(net2498),
    .B1(net1936),
    .B2(_06581_),
    .C1(net2446),
    .Y(_06582_));
 sky130_fd_sc_hd__nor2_1 _25879_ (.A(\inst$top.soc.cpu.gprf.mem[31][10] ),
    .B(net2477),
    .Y(_06583_));
 sky130_fd_sc_hd__o21ai_0 _25882_ (.A1(net2662),
    .A2(\inst$top.soc.cpu.gprf.mem[30][10] ),
    .B1(net2631),
    .Y(_06586_));
 sky130_fd_sc_hd__a221oi_1 _25884_ (.A1(net2515),
    .A2(\inst$top.soc.cpu.gprf.mem[28][10] ),
    .B1(net1963),
    .B2(\inst$top.soc.cpu.gprf.mem[29][10] ),
    .C1(net2454),
    .Y(_06588_));
 sky130_fd_sc_hd__o21ai_0 _25885_ (.A1(_06583_),
    .A2(_06586_),
    .B1(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__nor2_1 _25886_ (.A(\inst$top.soc.cpu.gprf.mem[27][10] ),
    .B(net2477),
    .Y(_06590_));
 sky130_fd_sc_hd__o21ai_0 _25887_ (.A1(net2671),
    .A2(\inst$top.soc.cpu.gprf.mem[26][10] ),
    .B1(net2631),
    .Y(_06591_));
 sky130_fd_sc_hd__a221oi_1 _25889_ (.A1(net2523),
    .A2(\inst$top.soc.cpu.gprf.mem[24][10] ),
    .B1(net1963),
    .B2(\inst$top.soc.cpu.gprf.mem[25][10] ),
    .C1(net2609),
    .Y(_06593_));
 sky130_fd_sc_hd__o21ai_0 _25890_ (.A1(_06590_),
    .A2(_06591_),
    .B1(_06593_),
    .Y(_06594_));
 sky130_fd_sc_hd__nand3_1 _25892_ (.A(_06589_),
    .B(_06594_),
    .C(net2599),
    .Y(_06596_));
 sky130_fd_sc_hd__a32oi_1 _25893_ (.A1(_06563_),
    .A2(_06568_),
    .A3(_06573_),
    .B1(_06582_),
    .B2(_06596_),
    .Y(_00001_));
 sky130_fd_sc_hd__nor2_1 _25894_ (.A(\inst$top.soc.cpu.gprf.mem[15][11] ),
    .B(net2474),
    .Y(_06597_));
 sky130_fd_sc_hd__o21ai_0 _25895_ (.A1(net2661),
    .A2(\inst$top.soc.cpu.gprf.mem[14][11] ),
    .B1(net2628),
    .Y(_06598_));
 sky130_fd_sc_hd__a221oi_1 _25896_ (.A1(net2514),
    .A2(\inst$top.soc.cpu.gprf.mem[12][11] ),
    .B1(net1953),
    .B2(\inst$top.soc.cpu.gprf.mem[13][11] ),
    .C1(net2455),
    .Y(_06599_));
 sky130_fd_sc_hd__o21ai_0 _25897_ (.A1(_06597_),
    .A2(_06598_),
    .B1(_06599_),
    .Y(_06600_));
 sky130_fd_sc_hd__nor2_1 _25898_ (.A(\inst$top.soc.cpu.gprf.mem[11][11] ),
    .B(net2474),
    .Y(_06601_));
 sky130_fd_sc_hd__o21ai_0 _25899_ (.A1(net2661),
    .A2(\inst$top.soc.cpu.gprf.mem[10][11] ),
    .B1(net2628),
    .Y(_06602_));
 sky130_fd_sc_hd__a221oi_1 _25900_ (.A1(net2515),
    .A2(\inst$top.soc.cpu.gprf.mem[8][11] ),
    .B1(net1954),
    .B2(\inst$top.soc.cpu.gprf.mem[9][11] ),
    .C1(net2609),
    .Y(_06603_));
 sky130_fd_sc_hd__o21ai_0 _25901_ (.A1(_06601_),
    .A2(_06602_),
    .B1(_06603_),
    .Y(_06604_));
 sky130_fd_sc_hd__nand3_1 _25902_ (.A(_06600_),
    .B(_06604_),
    .C(net2598),
    .Y(_06605_));
 sky130_fd_sc_hd__nor2_1 _25903_ (.A(\inst$top.soc.cpu.gprf.mem[7][11] ),
    .B(net2474),
    .Y(_06606_));
 sky130_fd_sc_hd__o21ai_0 _25906_ (.A1(net2664),
    .A2(\inst$top.soc.cpu.gprf.mem[6][11] ),
    .B1(net2632),
    .Y(_06609_));
 sky130_fd_sc_hd__a22oi_1 _25908_ (.A1(net2514),
    .A2(\inst$top.soc.cpu.gprf.mem[4][11] ),
    .B1(net1956),
    .B2(\inst$top.soc.cpu.gprf.mem[5][11] ),
    .Y(_06611_));
 sky130_fd_sc_hd__o21ai_0 _25909_ (.A1(_06606_),
    .A2(_06609_),
    .B1(_06611_),
    .Y(_06612_));
 sky130_fd_sc_hd__nand2_1 _25910_ (.A(_06612_),
    .B(net1934),
    .Y(_06613_));
 sky130_fd_sc_hd__nor2_1 _25911_ (.A(\inst$top.soc.cpu.gprf.mem[3][11] ),
    .B(net2474),
    .Y(_06614_));
 sky130_fd_sc_hd__o21ai_0 _25912_ (.A1(net2661),
    .A2(\inst$top.soc.cpu.gprf.mem[2][11] ),
    .B1(net2628),
    .Y(_06615_));
 sky130_fd_sc_hd__a22oi_1 _25913_ (.A1(net2514),
    .A2(\inst$top.soc.cpu.gprf.mem[0][11] ),
    .B1(net1956),
    .B2(\inst$top.soc.cpu.gprf.mem[1][11] ),
    .Y(_06616_));
 sky130_fd_sc_hd__o21ai_0 _25914_ (.A1(_06614_),
    .A2(_06615_),
    .B1(_06616_),
    .Y(_06617_));
 sky130_fd_sc_hd__a21oi_1 _25915_ (.A1(_06617_),
    .A2(net2499),
    .B1(net2596),
    .Y(_06618_));
 sky130_fd_sc_hd__nor2_1 _25916_ (.A(\inst$top.soc.cpu.gprf.mem[23][11] ),
    .B(net2474),
    .Y(_06619_));
 sky130_fd_sc_hd__o21ai_0 _25917_ (.A1(net2664),
    .A2(\inst$top.soc.cpu.gprf.mem[22][11] ),
    .B1(net2628),
    .Y(_06620_));
 sky130_fd_sc_hd__a22oi_1 _25918_ (.A1(net2514),
    .A2(\inst$top.soc.cpu.gprf.mem[20][11] ),
    .B1(net1956),
    .B2(\inst$top.soc.cpu.gprf.mem[21][11] ),
    .Y(_06621_));
 sky130_fd_sc_hd__o21ai_0 _25919_ (.A1(_06619_),
    .A2(_06620_),
    .B1(_06621_),
    .Y(_06622_));
 sky130_fd_sc_hd__nor2_1 _25920_ (.A(\inst$top.soc.cpu.gprf.mem[19][11] ),
    .B(net2474),
    .Y(_06623_));
 sky130_fd_sc_hd__o21ai_0 _25921_ (.A1(net2664),
    .A2(\inst$top.soc.cpu.gprf.mem[18][11] ),
    .B1(net2628),
    .Y(_06624_));
 sky130_fd_sc_hd__a22oi_1 _25922_ (.A1(net2517),
    .A2(\inst$top.soc.cpu.gprf.mem[16][11] ),
    .B1(net1954),
    .B2(\inst$top.soc.cpu.gprf.mem[17][11] ),
    .Y(_06625_));
 sky130_fd_sc_hd__o21ai_0 _25923_ (.A1(_06623_),
    .A2(_06624_),
    .B1(_06625_),
    .Y(_06626_));
 sky130_fd_sc_hd__a221oi_1 _25924_ (.A1(_06622_),
    .A2(net1936),
    .B1(net2499),
    .B2(_06626_),
    .C1(net2446),
    .Y(_06627_));
 sky130_fd_sc_hd__nor2_1 _25925_ (.A(\inst$top.soc.cpu.gprf.mem[31][11] ),
    .B(net2474),
    .Y(_06628_));
 sky130_fd_sc_hd__o21ai_0 _25926_ (.A1(net2662),
    .A2(\inst$top.soc.cpu.gprf.mem[30][11] ),
    .B1(net2628),
    .Y(_06629_));
 sky130_fd_sc_hd__a221oi_1 _25927_ (.A1(net2515),
    .A2(\inst$top.soc.cpu.gprf.mem[28][11] ),
    .B1(net1954),
    .B2(\inst$top.soc.cpu.gprf.mem[29][11] ),
    .C1(net2453),
    .Y(_06630_));
 sky130_fd_sc_hd__o21ai_0 _25928_ (.A1(_06628_),
    .A2(_06629_),
    .B1(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__nor2_1 _25929_ (.A(\inst$top.soc.cpu.gprf.mem[27][11] ),
    .B(net2474),
    .Y(_06632_));
 sky130_fd_sc_hd__o21ai_0 _25930_ (.A1(net2661),
    .A2(\inst$top.soc.cpu.gprf.mem[26][11] ),
    .B1(net2627),
    .Y(_06633_));
 sky130_fd_sc_hd__a221oi_1 _25931_ (.A1(net2514),
    .A2(\inst$top.soc.cpu.gprf.mem[24][11] ),
    .B1(net1953),
    .B2(\inst$top.soc.cpu.gprf.mem[25][11] ),
    .C1(net2609),
    .Y(_06634_));
 sky130_fd_sc_hd__o21ai_0 _25932_ (.A1(_06632_),
    .A2(_06633_),
    .B1(_06634_),
    .Y(_06635_));
 sky130_fd_sc_hd__nand3_1 _25933_ (.A(_06631_),
    .B(_06635_),
    .C(net2599),
    .Y(_06636_));
 sky130_fd_sc_hd__a32oi_1 _25934_ (.A1(_06605_),
    .A2(_06613_),
    .A3(_06618_),
    .B1(_06627_),
    .B2(_06636_),
    .Y(_00002_));
 sky130_fd_sc_hd__nor2_1 _25935_ (.A(\inst$top.soc.cpu.gprf.mem[11][12] ),
    .B(net2492),
    .Y(_06637_));
 sky130_fd_sc_hd__o21ai_0 _25938_ (.A1(net2683),
    .A2(\inst$top.soc.cpu.gprf.mem[10][12] ),
    .B1(net2649),
    .Y(_06640_));
 sky130_fd_sc_hd__a221oi_1 _25940_ (.A1(net2533),
    .A2(\inst$top.soc.cpu.gprf.mem[8][12] ),
    .B1(net1973),
    .B2(\inst$top.soc.cpu.gprf.mem[9][12] ),
    .C1(net2613),
    .Y(_06642_));
 sky130_fd_sc_hd__o21ai_0 _25941_ (.A1(_06637_),
    .A2(_06640_),
    .B1(_06642_),
    .Y(_06643_));
 sky130_fd_sc_hd__nor2_1 _25942_ (.A(\inst$top.soc.cpu.gprf.mem[15][12] ),
    .B(net2493),
    .Y(_06644_));
 sky130_fd_sc_hd__o21ai_0 _25943_ (.A1(net2683),
    .A2(\inst$top.soc.cpu.gprf.mem[14][12] ),
    .B1(net2649),
    .Y(_06645_));
 sky130_fd_sc_hd__a221oi_1 _25945_ (.A1(net2533),
    .A2(\inst$top.soc.cpu.gprf.mem[12][12] ),
    .B1(net1973),
    .B2(\inst$top.soc.cpu.gprf.mem[13][12] ),
    .C1(net2458),
    .Y(_06647_));
 sky130_fd_sc_hd__o21ai_0 _25946_ (.A1(_06644_),
    .A2(_06645_),
    .B1(_06647_),
    .Y(_06648_));
 sky130_fd_sc_hd__nand3_1 _25947_ (.A(_06643_),
    .B(_06648_),
    .C(net2604),
    .Y(_06649_));
 sky130_fd_sc_hd__nor2_1 _25948_ (.A(\inst$top.soc.cpu.gprf.mem[7][12] ),
    .B(net2492),
    .Y(_06650_));
 sky130_fd_sc_hd__o21ai_0 _25949_ (.A1(net2681),
    .A2(\inst$top.soc.cpu.gprf.mem[6][12] ),
    .B1(net2648),
    .Y(_06651_));
 sky130_fd_sc_hd__a22oi_1 _25950_ (.A1(net2532),
    .A2(\inst$top.soc.cpu.gprf.mem[4][12] ),
    .B1(net1972),
    .B2(\inst$top.soc.cpu.gprf.mem[5][12] ),
    .Y(_06652_));
 sky130_fd_sc_hd__o21ai_0 _25951_ (.A1(_06650_),
    .A2(_06651_),
    .B1(_06652_),
    .Y(_06653_));
 sky130_fd_sc_hd__nand2_1 _25953_ (.A(_06653_),
    .B(net1939),
    .Y(_06655_));
 sky130_fd_sc_hd__nor2_1 _25954_ (.A(\inst$top.soc.cpu.gprf.mem[3][12] ),
    .B(net2492),
    .Y(_06656_));
 sky130_fd_sc_hd__o21ai_0 _25955_ (.A1(net2683),
    .A2(\inst$top.soc.cpu.gprf.mem[2][12] ),
    .B1(net2648),
    .Y(_06657_));
 sky130_fd_sc_hd__a22oi_1 _25956_ (.A1(net2532),
    .A2(\inst$top.soc.cpu.gprf.mem[0][12] ),
    .B1(net1972),
    .B2(\inst$top.soc.cpu.gprf.mem[1][12] ),
    .Y(_06658_));
 sky130_fd_sc_hd__o21ai_0 _25957_ (.A1(_06656_),
    .A2(_06657_),
    .B1(_06658_),
    .Y(_06659_));
 sky130_fd_sc_hd__a21oi_1 _25959_ (.A1(_06659_),
    .A2(net2502),
    .B1(net2594),
    .Y(_06661_));
 sky130_fd_sc_hd__nor2_1 _25960_ (.A(\inst$top.soc.cpu.gprf.mem[19][12] ),
    .B(net2492),
    .Y(_06662_));
 sky130_fd_sc_hd__o21ai_0 _25961_ (.A1(net2683),
    .A2(\inst$top.soc.cpu.gprf.mem[18][12] ),
    .B1(net2648),
    .Y(_06663_));
 sky130_fd_sc_hd__a22oi_1 _25962_ (.A1(net2533),
    .A2(\inst$top.soc.cpu.gprf.mem[16][12] ),
    .B1(net1973),
    .B2(\inst$top.soc.cpu.gprf.mem[17][12] ),
    .Y(_06664_));
 sky130_fd_sc_hd__o21ai_0 _25963_ (.A1(_06662_),
    .A2(_06663_),
    .B1(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__nor2_1 _25964_ (.A(\inst$top.soc.cpu.gprf.mem[23][12] ),
    .B(net2493),
    .Y(_06666_));
 sky130_fd_sc_hd__o21ai_0 _25965_ (.A1(net2683),
    .A2(\inst$top.soc.cpu.gprf.mem[22][12] ),
    .B1(net2648),
    .Y(_06667_));
 sky130_fd_sc_hd__a22oi_1 _25966_ (.A1(net2533),
    .A2(\inst$top.soc.cpu.gprf.mem[20][12] ),
    .B1(net1973),
    .B2(\inst$top.soc.cpu.gprf.mem[21][12] ),
    .Y(_06668_));
 sky130_fd_sc_hd__o21ai_0 _25967_ (.A1(_06666_),
    .A2(_06667_),
    .B1(_06668_),
    .Y(_06669_));
 sky130_fd_sc_hd__a221oi_1 _25968_ (.A1(_06665_),
    .A2(net2502),
    .B1(net1939),
    .B2(_06669_),
    .C1(net2447),
    .Y(_06670_));
 sky130_fd_sc_hd__nor2_1 _25970_ (.A(\inst$top.soc.cpu.gprf.mem[31][12] ),
    .B(net2492),
    .Y(_06672_));
 sky130_fd_sc_hd__o21ai_0 _25971_ (.A1(net2683),
    .A2(\inst$top.soc.cpu.gprf.mem[30][12] ),
    .B1(net2648),
    .Y(_06673_));
 sky130_fd_sc_hd__a221oi_1 _25974_ (.A1(net2533),
    .A2(\inst$top.soc.cpu.gprf.mem[28][12] ),
    .B1(net1973),
    .B2(\inst$top.soc.cpu.gprf.mem[29][12] ),
    .C1(net2458),
    .Y(_06676_));
 sky130_fd_sc_hd__o21ai_0 _25975_ (.A1(_06672_),
    .A2(_06673_),
    .B1(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__nor2_1 _25976_ (.A(\inst$top.soc.cpu.gprf.mem[27][12] ),
    .B(net2492),
    .Y(_06678_));
 sky130_fd_sc_hd__o21ai_0 _25979_ (.A1(net2681),
    .A2(\inst$top.soc.cpu.gprf.mem[26][12] ),
    .B1(net2648),
    .Y(_06681_));
 sky130_fd_sc_hd__a221oi_1 _25982_ (.A1(net2532),
    .A2(\inst$top.soc.cpu.gprf.mem[24][12] ),
    .B1(net1972),
    .B2(\inst$top.soc.cpu.gprf.mem[25][12] ),
    .C1(net2614),
    .Y(_06684_));
 sky130_fd_sc_hd__o21ai_0 _25983_ (.A1(_06678_),
    .A2(_06681_),
    .B1(_06684_),
    .Y(_06685_));
 sky130_fd_sc_hd__nand3_1 _25984_ (.A(_06677_),
    .B(_06685_),
    .C(net2604),
    .Y(_06686_));
 sky130_fd_sc_hd__a32oi_1 _25985_ (.A1(_06649_),
    .A2(_06655_),
    .A3(_06661_),
    .B1(_06670_),
    .B2(_06686_),
    .Y(_00003_));
 sky130_fd_sc_hd__nor2_1 _25986_ (.A(\inst$top.soc.cpu.gprf.mem[15][13] ),
    .B(net2466),
    .Y(_06687_));
 sky130_fd_sc_hd__o21ai_0 _25987_ (.A1(net2659),
    .A2(\inst$top.soc.cpu.gprf.mem[14][13] ),
    .B1(net2623),
    .Y(_06688_));
 sky130_fd_sc_hd__a221oi_1 _25988_ (.A1(net2512),
    .A2(\inst$top.soc.cpu.gprf.mem[12][13] ),
    .B1(net1951),
    .B2(\inst$top.soc.cpu.gprf.mem[13][13] ),
    .C1(net2453),
    .Y(_06689_));
 sky130_fd_sc_hd__o21ai_0 _25989_ (.A1(_06687_),
    .A2(_06688_),
    .B1(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__nor2_1 _25990_ (.A(\inst$top.soc.cpu.gprf.mem[11][13] ),
    .B(net2467),
    .Y(_06691_));
 sky130_fd_sc_hd__o21ai_0 _25991_ (.A1(net2659),
    .A2(\inst$top.soc.cpu.gprf.mem[10][13] ),
    .B1(net2624),
    .Y(_06692_));
 sky130_fd_sc_hd__a221oi_1 _25992_ (.A1(net2512),
    .A2(\inst$top.soc.cpu.gprf.mem[8][13] ),
    .B1(net1951),
    .B2(\inst$top.soc.cpu.gprf.mem[9][13] ),
    .C1(net2610),
    .Y(_06693_));
 sky130_fd_sc_hd__o21ai_0 _25993_ (.A1(_06691_),
    .A2(_06692_),
    .B1(_06693_),
    .Y(_06694_));
 sky130_fd_sc_hd__nand3_1 _25994_ (.A(_06690_),
    .B(_06694_),
    .C(net2598),
    .Y(_06695_));
 sky130_fd_sc_hd__nor2_1 _25996_ (.A(\inst$top.soc.cpu.gprf.mem[7][13] ),
    .B(net2470),
    .Y(_06697_));
 sky130_fd_sc_hd__o21ai_0 _25997_ (.A1(net2659),
    .A2(\inst$top.soc.cpu.gprf.mem[6][13] ),
    .B1(net2624),
    .Y(_06698_));
 sky130_fd_sc_hd__a22oi_1 _25999_ (.A1(net2512),
    .A2(\inst$top.soc.cpu.gprf.mem[4][13] ),
    .B1(net1951),
    .B2(\inst$top.soc.cpu.gprf.mem[5][13] ),
    .Y(_06700_));
 sky130_fd_sc_hd__o21ai_0 _26000_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__nand2_1 _26001_ (.A(_06701_),
    .B(net1935),
    .Y(_06702_));
 sky130_fd_sc_hd__nor2_1 _26002_ (.A(\inst$top.soc.cpu.gprf.mem[3][13] ),
    .B(net2470),
    .Y(_06703_));
 sky130_fd_sc_hd__o21ai_0 _26005_ (.A1(net2659),
    .A2(\inst$top.soc.cpu.gprf.mem[2][13] ),
    .B1(net2624),
    .Y(_06706_));
 sky130_fd_sc_hd__a22oi_1 _26006_ (.A1(net2512),
    .A2(\inst$top.soc.cpu.gprf.mem[0][13] ),
    .B1(net1951),
    .B2(\inst$top.soc.cpu.gprf.mem[1][13] ),
    .Y(_06707_));
 sky130_fd_sc_hd__o21ai_0 _26007_ (.A1(_06703_),
    .A2(_06706_),
    .B1(_06707_),
    .Y(_06708_));
 sky130_fd_sc_hd__a21oi_1 _26008_ (.A1(_06708_),
    .A2(net2497),
    .B1(net2592),
    .Y(_06709_));
 sky130_fd_sc_hd__nor2_1 _26010_ (.A(\inst$top.soc.cpu.gprf.mem[23][13] ),
    .B(net2467),
    .Y(_06711_));
 sky130_fd_sc_hd__o21ai_0 _26011_ (.A1(net2659),
    .A2(\inst$top.soc.cpu.gprf.mem[22][13] ),
    .B1(net2624),
    .Y(_06712_));
 sky130_fd_sc_hd__a22oi_1 _26012_ (.A1(net2512),
    .A2(\inst$top.soc.cpu.gprf.mem[20][13] ),
    .B1(net1951),
    .B2(\inst$top.soc.cpu.gprf.mem[21][13] ),
    .Y(_06713_));
 sky130_fd_sc_hd__o21ai_0 _26013_ (.A1(_06711_),
    .A2(_06712_),
    .B1(_06713_),
    .Y(_06714_));
 sky130_fd_sc_hd__nor2_1 _26015_ (.A(\inst$top.soc.cpu.gprf.mem[19][13] ),
    .B(net2467),
    .Y(_06716_));
 sky130_fd_sc_hd__o21ai_0 _26016_ (.A1(net2659),
    .A2(\inst$top.soc.cpu.gprf.mem[18][13] ),
    .B1(net2621),
    .Y(_06717_));
 sky130_fd_sc_hd__a22oi_1 _26017_ (.A1(net2512),
    .A2(\inst$top.soc.cpu.gprf.mem[16][13] ),
    .B1(net1951),
    .B2(\inst$top.soc.cpu.gprf.mem[17][13] ),
    .Y(_06718_));
 sky130_fd_sc_hd__o21ai_0 _26018_ (.A1(_06716_),
    .A2(_06717_),
    .B1(_06718_),
    .Y(_06719_));
 sky130_fd_sc_hd__a221oi_1 _26019_ (.A1(_06714_),
    .A2(net1935),
    .B1(net2497),
    .B2(_06719_),
    .C1(net2446),
    .Y(_06720_));
 sky130_fd_sc_hd__nor2_1 _26020_ (.A(\inst$top.soc.cpu.gprf.mem[31][13] ),
    .B(net2470),
    .Y(_06721_));
 sky130_fd_sc_hd__o21ai_0 _26021_ (.A1(net2659),
    .A2(\inst$top.soc.cpu.gprf.mem[30][13] ),
    .B1(net2624),
    .Y(_06722_));
 sky130_fd_sc_hd__a221oi_1 _26022_ (.A1(net2512),
    .A2(\inst$top.soc.cpu.gprf.mem[28][13] ),
    .B1(net1951),
    .B2(\inst$top.soc.cpu.gprf.mem[29][13] ),
    .C1(net2453),
    .Y(_06723_));
 sky130_fd_sc_hd__o21ai_0 _26023_ (.A1(_06721_),
    .A2(_06722_),
    .B1(_06723_),
    .Y(_06724_));
 sky130_fd_sc_hd__nor2_1 _26024_ (.A(\inst$top.soc.cpu.gprf.mem[27][13] ),
    .B(net2470),
    .Y(_06725_));
 sky130_fd_sc_hd__o21ai_0 _26025_ (.A1(net2659),
    .A2(\inst$top.soc.cpu.gprf.mem[26][13] ),
    .B1(net2624),
    .Y(_06726_));
 sky130_fd_sc_hd__a221oi_1 _26026_ (.A1(net2512),
    .A2(\inst$top.soc.cpu.gprf.mem[24][13] ),
    .B1(net1951),
    .B2(\inst$top.soc.cpu.gprf.mem[25][13] ),
    .C1(net2610),
    .Y(_06727_));
 sky130_fd_sc_hd__o21ai_0 _26027_ (.A1(_06725_),
    .A2(_06726_),
    .B1(_06727_),
    .Y(_06728_));
 sky130_fd_sc_hd__nand3_1 _26028_ (.A(_06724_),
    .B(_06728_),
    .C(net2598),
    .Y(_06729_));
 sky130_fd_sc_hd__a32oi_1 _26029_ (.A1(_06695_),
    .A2(_06702_),
    .A3(_06709_),
    .B1(_06720_),
    .B2(_06729_),
    .Y(_00004_));
 sky130_fd_sc_hd__nor2_1 _26031_ (.A(\inst$top.soc.cpu.gprf.mem[11][14] ),
    .B(net2485),
    .Y(_06731_));
 sky130_fd_sc_hd__o21ai_0 _26032_ (.A1(net2678),
    .A2(\inst$top.soc.cpu.gprf.mem[10][14] ),
    .B1(net2640),
    .Y(_06732_));
 sky130_fd_sc_hd__a221oi_1 _26033_ (.A1(net2530),
    .A2(\inst$top.soc.cpu.gprf.mem[8][14] ),
    .B1(net1970),
    .B2(\inst$top.soc.cpu.gprf.mem[9][14] ),
    .C1(net2612),
    .Y(_06733_));
 sky130_fd_sc_hd__o21ai_0 _26034_ (.A1(_06731_),
    .A2(_06732_),
    .B1(_06733_),
    .Y(_06734_));
 sky130_fd_sc_hd__nor2_1 _26035_ (.A(\inst$top.soc.cpu.gprf.mem[15][14] ),
    .B(net2486),
    .Y(_06735_));
 sky130_fd_sc_hd__o21ai_0 _26036_ (.A1(net2678),
    .A2(\inst$top.soc.cpu.gprf.mem[14][14] ),
    .B1(net2638),
    .Y(_06736_));
 sky130_fd_sc_hd__a221oi_1 _26037_ (.A1(net2529),
    .A2(\inst$top.soc.cpu.gprf.mem[12][14] ),
    .B1(net1970),
    .B2(\inst$top.soc.cpu.gprf.mem[13][14] ),
    .C1(net2457),
    .Y(_06737_));
 sky130_fd_sc_hd__o21ai_0 _26038_ (.A1(_06735_),
    .A2(_06736_),
    .B1(_06737_),
    .Y(_06738_));
 sky130_fd_sc_hd__nand3_1 _26039_ (.A(_06734_),
    .B(_06738_),
    .C(net2603),
    .Y(_06739_));
 sky130_fd_sc_hd__nor2_1 _26040_ (.A(\inst$top.soc.cpu.gprf.mem[7][14] ),
    .B(net2483),
    .Y(_06740_));
 sky130_fd_sc_hd__o21ai_0 _26041_ (.A1(net2677),
    .A2(\inst$top.soc.cpu.gprf.mem[6][14] ),
    .B1(net2637),
    .Y(_06741_));
 sky130_fd_sc_hd__a22oi_1 _26042_ (.A1(net2529),
    .A2(\inst$top.soc.cpu.gprf.mem[4][14] ),
    .B1(net1969),
    .B2(\inst$top.soc.cpu.gprf.mem[5][14] ),
    .Y(_06742_));
 sky130_fd_sc_hd__o21ai_0 _26043_ (.A1(_06740_),
    .A2(_06741_),
    .B1(_06742_),
    .Y(_06743_));
 sky130_fd_sc_hd__nand2_1 _26044_ (.A(_06743_),
    .B(net1938),
    .Y(_06744_));
 sky130_fd_sc_hd__nor2_1 _26046_ (.A(\inst$top.soc.cpu.gprf.mem[3][14] ),
    .B(net2484),
    .Y(_06746_));
 sky130_fd_sc_hd__o21ai_0 _26047_ (.A1(net2679),
    .A2(\inst$top.soc.cpu.gprf.mem[2][14] ),
    .B1(net2639),
    .Y(_06747_));
 sky130_fd_sc_hd__a22oi_1 _26048_ (.A1(net2527),
    .A2(\inst$top.soc.cpu.gprf.mem[0][14] ),
    .B1(net1967),
    .B2(\inst$top.soc.cpu.gprf.mem[1][14] ),
    .Y(_06748_));
 sky130_fd_sc_hd__o21ai_0 _26049_ (.A1(_06746_),
    .A2(_06747_),
    .B1(_06748_),
    .Y(_06749_));
 sky130_fd_sc_hd__a21oi_1 _26050_ (.A1(_06749_),
    .A2(net2501),
    .B1(net2593),
    .Y(_06750_));
 sky130_fd_sc_hd__nor2_1 _26051_ (.A(\inst$top.soc.cpu.gprf.mem[23][14] ),
    .B(net2486),
    .Y(_06751_));
 sky130_fd_sc_hd__o21ai_0 _26054_ (.A1(net2678),
    .A2(\inst$top.soc.cpu.gprf.mem[22][14] ),
    .B1(net2638),
    .Y(_06754_));
 sky130_fd_sc_hd__a22oi_1 _26055_ (.A1(net2529),
    .A2(\inst$top.soc.cpu.gprf.mem[20][14] ),
    .B1(net1969),
    .B2(\inst$top.soc.cpu.gprf.mem[21][14] ),
    .Y(_06755_));
 sky130_fd_sc_hd__o21ai_0 _26056_ (.A1(_06751_),
    .A2(_06754_),
    .B1(_06755_),
    .Y(_06756_));
 sky130_fd_sc_hd__nor2_1 _26057_ (.A(\inst$top.soc.cpu.gprf.mem[19][14] ),
    .B(net2485),
    .Y(_06757_));
 sky130_fd_sc_hd__o21ai_0 _26060_ (.A1(net2679),
    .A2(\inst$top.soc.cpu.gprf.mem[18][14] ),
    .B1(net2640),
    .Y(_06760_));
 sky130_fd_sc_hd__a22oi_1 _26061_ (.A1(net2530),
    .A2(\inst$top.soc.cpu.gprf.mem[16][14] ),
    .B1(net1970),
    .B2(\inst$top.soc.cpu.gprf.mem[17][14] ),
    .Y(_06761_));
 sky130_fd_sc_hd__o21ai_0 _26062_ (.A1(_06757_),
    .A2(_06760_),
    .B1(_06761_),
    .Y(_06762_));
 sky130_fd_sc_hd__a221oi_1 _26064_ (.A1(_06756_),
    .A2(net1938),
    .B1(net2501),
    .B2(_06762_),
    .C1(net2448),
    .Y(_06764_));
 sky130_fd_sc_hd__nor2_1 _26065_ (.A(\inst$top.soc.cpu.gprf.mem[31][14] ),
    .B(net2484),
    .Y(_06765_));
 sky130_fd_sc_hd__o21ai_0 _26066_ (.A1(net2677),
    .A2(\inst$top.soc.cpu.gprf.mem[30][14] ),
    .B1(net2638),
    .Y(_06766_));
 sky130_fd_sc_hd__a221oi_1 _26067_ (.A1(net2529),
    .A2(\inst$top.soc.cpu.gprf.mem[28][14] ),
    .B1(net1969),
    .B2(\inst$top.soc.cpu.gprf.mem[29][14] ),
    .C1(net2457),
    .Y(_06767_));
 sky130_fd_sc_hd__o21ai_0 _26068_ (.A1(_06765_),
    .A2(_06766_),
    .B1(_06767_),
    .Y(_06768_));
 sky130_fd_sc_hd__nor2_1 _26070_ (.A(\inst$top.soc.cpu.gprf.mem[27][14] ),
    .B(net2484),
    .Y(_06770_));
 sky130_fd_sc_hd__o21ai_0 _26071_ (.A1(net2676),
    .A2(\inst$top.soc.cpu.gprf.mem[26][14] ),
    .B1(net2639),
    .Y(_06771_));
 sky130_fd_sc_hd__a221oi_1 _26072_ (.A1(net2528),
    .A2(\inst$top.soc.cpu.gprf.mem[24][14] ),
    .B1(net1968),
    .B2(\inst$top.soc.cpu.gprf.mem[25][14] ),
    .C1(net2612),
    .Y(_06772_));
 sky130_fd_sc_hd__o21ai_0 _26073_ (.A1(_06770_),
    .A2(_06771_),
    .B1(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__nand3_1 _26074_ (.A(_06768_),
    .B(_06773_),
    .C(net2604),
    .Y(_06774_));
 sky130_fd_sc_hd__a32oi_1 _26075_ (.A1(_06739_),
    .A2(_06744_),
    .A3(_06750_),
    .B1(_06764_),
    .B2(_06774_),
    .Y(_00005_));
 sky130_fd_sc_hd__nor2_1 _26076_ (.A(\inst$top.soc.cpu.gprf.mem[31][15] ),
    .B(net2485),
    .Y(_06775_));
 sky130_fd_sc_hd__o21ai_0 _26077_ (.A1(net2678),
    .A2(\inst$top.soc.cpu.gprf.mem[30][15] ),
    .B1(net2640),
    .Y(_06776_));
 sky130_fd_sc_hd__a221oi_1 _26078_ (.A1(net2530),
    .A2(\inst$top.soc.cpu.gprf.mem[28][15] ),
    .B1(net1970),
    .B2(\inst$top.soc.cpu.gprf.mem[29][15] ),
    .C1(net2457),
    .Y(_06777_));
 sky130_fd_sc_hd__o21ai_0 _26079_ (.A1(_06775_),
    .A2(_06776_),
    .B1(_06777_),
    .Y(_06778_));
 sky130_fd_sc_hd__nor2_1 _26080_ (.A(\inst$top.soc.cpu.gprf.mem[27][15] ),
    .B(net2484),
    .Y(_06779_));
 sky130_fd_sc_hd__o21ai_0 _26081_ (.A1(net2678),
    .A2(\inst$top.soc.cpu.gprf.mem[26][15] ),
    .B1(net2639),
    .Y(_06780_));
 sky130_fd_sc_hd__a221oi_1 _26082_ (.A1(net2530),
    .A2(\inst$top.soc.cpu.gprf.mem[24][15] ),
    .B1(net1970),
    .B2(\inst$top.soc.cpu.gprf.mem[25][15] ),
    .C1(net2612),
    .Y(_06781_));
 sky130_fd_sc_hd__o21ai_0 _26083_ (.A1(_06779_),
    .A2(_06780_),
    .B1(_06781_),
    .Y(_06782_));
 sky130_fd_sc_hd__nand3_1 _26084_ (.A(_06778_),
    .B(_06782_),
    .C(net2603),
    .Y(_06783_));
 sky130_fd_sc_hd__nor2_1 _26085_ (.A(\inst$top.soc.cpu.gprf.mem[19][15] ),
    .B(net2484),
    .Y(_06784_));
 sky130_fd_sc_hd__o21ai_0 _26086_ (.A1(net2678),
    .A2(\inst$top.soc.cpu.gprf.mem[18][15] ),
    .B1(net2639),
    .Y(_06785_));
 sky130_fd_sc_hd__a22oi_1 _26087_ (.A1(net2530),
    .A2(\inst$top.soc.cpu.gprf.mem[16][15] ),
    .B1(net1970),
    .B2(\inst$top.soc.cpu.gprf.mem[17][15] ),
    .Y(_06786_));
 sky130_fd_sc_hd__o21ai_0 _26088_ (.A1(_06784_),
    .A2(_06785_),
    .B1(_06786_),
    .Y(_06787_));
 sky130_fd_sc_hd__nand2_1 _26089_ (.A(_06787_),
    .B(net2501),
    .Y(_06788_));
 sky130_fd_sc_hd__nor2_1 _26090_ (.A(\inst$top.soc.cpu.gprf.mem[23][15] ),
    .B(net2485),
    .Y(_06789_));
 sky130_fd_sc_hd__o21ai_0 _26091_ (.A1(net2679),
    .A2(\inst$top.soc.cpu.gprf.mem[22][15] ),
    .B1(net2640),
    .Y(_06790_));
 sky130_fd_sc_hd__a22oi_1 _26093_ (.A1(net2536),
    .A2(\inst$top.soc.cpu.gprf.mem[20][15] ),
    .B1(net1970),
    .B2(\inst$top.soc.cpu.gprf.mem[21][15] ),
    .Y(_06792_));
 sky130_fd_sc_hd__o21ai_0 _26094_ (.A1(_06789_),
    .A2(_06790_),
    .B1(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__a21oi_1 _26095_ (.A1(_06793_),
    .A2(net1938),
    .B1(net2447),
    .Y(_06794_));
 sky130_fd_sc_hd__nor2_1 _26096_ (.A(\inst$top.soc.cpu.gprf.mem[3][15] ),
    .B(net2484),
    .Y(_06795_));
 sky130_fd_sc_hd__o21ai_0 _26097_ (.A1(net2679),
    .A2(\inst$top.soc.cpu.gprf.mem[2][15] ),
    .B1(net2639),
    .Y(_06796_));
 sky130_fd_sc_hd__a22oi_1 _26098_ (.A1(net2528),
    .A2(\inst$top.soc.cpu.gprf.mem[0][15] ),
    .B1(net1968),
    .B2(\inst$top.soc.cpu.gprf.mem[1][15] ),
    .Y(_06797_));
 sky130_fd_sc_hd__o21ai_0 _26099_ (.A1(_06795_),
    .A2(_06796_),
    .B1(_06797_),
    .Y(_06798_));
 sky130_fd_sc_hd__nor2_1 _26100_ (.A(\inst$top.soc.cpu.gprf.mem[7][15] ),
    .B(net2484),
    .Y(_06799_));
 sky130_fd_sc_hd__o21ai_0 _26101_ (.A1(net2679),
    .A2(\inst$top.soc.cpu.gprf.mem[6][15] ),
    .B1(net2639),
    .Y(_06800_));
 sky130_fd_sc_hd__a22oi_1 _26102_ (.A1(net2528),
    .A2(\inst$top.soc.cpu.gprf.mem[4][15] ),
    .B1(net1968),
    .B2(\inst$top.soc.cpu.gprf.mem[5][15] ),
    .Y(_06801_));
 sky130_fd_sc_hd__o21ai_0 _26103_ (.A1(_06799_),
    .A2(_06800_),
    .B1(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__a221oi_1 _26104_ (.A1(_06798_),
    .A2(net2501),
    .B1(net1938),
    .B2(_06802_),
    .C1(net2593),
    .Y(_06803_));
 sky130_fd_sc_hd__nor2_1 _26105_ (.A(\inst$top.soc.cpu.gprf.mem[15][15] ),
    .B(net2484),
    .Y(_06804_));
 sky130_fd_sc_hd__o21ai_0 _26106_ (.A1(net2678),
    .A2(\inst$top.soc.cpu.gprf.mem[14][15] ),
    .B1(net2639),
    .Y(_06805_));
 sky130_fd_sc_hd__a221oi_1 _26107_ (.A1(net2530),
    .A2(\inst$top.soc.cpu.gprf.mem[12][15] ),
    .B1(net1970),
    .B2(\inst$top.soc.cpu.gprf.mem[13][15] ),
    .C1(net2457),
    .Y(_06806_));
 sky130_fd_sc_hd__o21ai_0 _26108_ (.A1(_06804_),
    .A2(_06805_),
    .B1(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__nor2_1 _26109_ (.A(\inst$top.soc.cpu.gprf.mem[11][15] ),
    .B(net2485),
    .Y(_06808_));
 sky130_fd_sc_hd__o21ai_0 _26110_ (.A1(net2678),
    .A2(\inst$top.soc.cpu.gprf.mem[10][15] ),
    .B1(net2640),
    .Y(_06809_));
 sky130_fd_sc_hd__a221oi_1 _26111_ (.A1(net2530),
    .A2(\inst$top.soc.cpu.gprf.mem[8][15] ),
    .B1(net1976),
    .B2(\inst$top.soc.cpu.gprf.mem[9][15] ),
    .C1(net2612),
    .Y(_06810_));
 sky130_fd_sc_hd__o21ai_0 _26112_ (.A1(_06808_),
    .A2(_06809_),
    .B1(_06810_),
    .Y(_06811_));
 sky130_fd_sc_hd__nand3_1 _26113_ (.A(_06807_),
    .B(_06811_),
    .C(net2603),
    .Y(_06812_));
 sky130_fd_sc_hd__a32oi_1 _26114_ (.A1(_06783_),
    .A2(_06788_),
    .A3(_06794_),
    .B1(_06803_),
    .B2(_06812_),
    .Y(_00006_));
 sky130_fd_sc_hd__nor2_1 _26115_ (.A(\inst$top.soc.cpu.gprf.mem[11][16] ),
    .B(net2489),
    .Y(_06813_));
 sky130_fd_sc_hd__o21ai_0 _26116_ (.A1(net2681),
    .A2(\inst$top.soc.cpu.gprf.mem[10][16] ),
    .B1(net2644),
    .Y(_06814_));
 sky130_fd_sc_hd__a221oi_1 _26117_ (.A1(net2532),
    .A2(\inst$top.soc.cpu.gprf.mem[8][16] ),
    .B1(net1972),
    .B2(\inst$top.soc.cpu.gprf.mem[9][16] ),
    .C1(net2613),
    .Y(_06815_));
 sky130_fd_sc_hd__o21ai_0 _26118_ (.A1(_06813_),
    .A2(_06814_),
    .B1(_06815_),
    .Y(_06816_));
 sky130_fd_sc_hd__nor2_1 _26119_ (.A(\inst$top.soc.cpu.gprf.mem[15][16] ),
    .B(net2488),
    .Y(_06817_));
 sky130_fd_sc_hd__o21ai_0 _26120_ (.A1(net2673),
    .A2(\inst$top.soc.cpu.gprf.mem[14][16] ),
    .B1(net2643),
    .Y(_06818_));
 sky130_fd_sc_hd__a221oi_1 _26122_ (.A1(net2525),
    .A2(\inst$top.soc.cpu.gprf.mem[12][16] ),
    .B1(net1972),
    .B2(\inst$top.soc.cpu.gprf.mem[13][16] ),
    .C1(net2459),
    .Y(_06820_));
 sky130_fd_sc_hd__o21ai_0 _26123_ (.A1(_06817_),
    .A2(_06818_),
    .B1(_06820_),
    .Y(_06821_));
 sky130_fd_sc_hd__nand3_1 _26124_ (.A(_06816_),
    .B(_06821_),
    .C(net2601),
    .Y(_06822_));
 sky130_fd_sc_hd__nor2_1 _26125_ (.A(\inst$top.soc.cpu.gprf.mem[7][16] ),
    .B(net2489),
    .Y(_06823_));
 sky130_fd_sc_hd__o21ai_0 _26126_ (.A1(net2681),
    .A2(\inst$top.soc.cpu.gprf.mem[6][16] ),
    .B1(net2644),
    .Y(_06824_));
 sky130_fd_sc_hd__a22oi_1 _26127_ (.A1(net2532),
    .A2(\inst$top.soc.cpu.gprf.mem[4][16] ),
    .B1(net1972),
    .B2(\inst$top.soc.cpu.gprf.mem[5][16] ),
    .Y(_06825_));
 sky130_fd_sc_hd__o21ai_0 _26128_ (.A1(_06823_),
    .A2(_06824_),
    .B1(_06825_),
    .Y(_06826_));
 sky130_fd_sc_hd__nand2_1 _26129_ (.A(_06826_),
    .B(net1940),
    .Y(_06827_));
 sky130_fd_sc_hd__nor2_1 _26130_ (.A(\inst$top.soc.cpu.gprf.mem[3][16] ),
    .B(net2489),
    .Y(_06828_));
 sky130_fd_sc_hd__o21ai_0 _26131_ (.A1(net2673),
    .A2(\inst$top.soc.cpu.gprf.mem[2][16] ),
    .B1(net2644),
    .Y(_06829_));
 sky130_fd_sc_hd__a22oi_1 _26132_ (.A1(net2525),
    .A2(\inst$top.soc.cpu.gprf.mem[0][16] ),
    .B1(net1965),
    .B2(\inst$top.soc.cpu.gprf.mem[1][16] ),
    .Y(_06830_));
 sky130_fd_sc_hd__o21ai_0 _26133_ (.A1(_06828_),
    .A2(_06829_),
    .B1(_06830_),
    .Y(_06831_));
 sky130_fd_sc_hd__a21oi_1 _26134_ (.A1(_06831_),
    .A2(net2503),
    .B1(net2594),
    .Y(_06832_));
 sky130_fd_sc_hd__nor2_1 _26135_ (.A(\inst$top.soc.cpu.gprf.mem[19][16] ),
    .B(net2489),
    .Y(_06833_));
 sky130_fd_sc_hd__o21ai_0 _26136_ (.A1(net2673),
    .A2(\inst$top.soc.cpu.gprf.mem[18][16] ),
    .B1(net2644),
    .Y(_06834_));
 sky130_fd_sc_hd__a22oi_1 _26139_ (.A1(net2525),
    .A2(\inst$top.soc.cpu.gprf.mem[16][16] ),
    .B1(net1965),
    .B2(\inst$top.soc.cpu.gprf.mem[17][16] ),
    .Y(_06837_));
 sky130_fd_sc_hd__o21ai_0 _26140_ (.A1(_06833_),
    .A2(_06834_),
    .B1(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__nor2_1 _26141_ (.A(\inst$top.soc.cpu.gprf.mem[23][16] ),
    .B(net2488),
    .Y(_06839_));
 sky130_fd_sc_hd__o21ai_0 _26142_ (.A1(net2673),
    .A2(\inst$top.soc.cpu.gprf.mem[22][16] ),
    .B1(net2643),
    .Y(_06840_));
 sky130_fd_sc_hd__a22oi_1 _26145_ (.A1(net2525),
    .A2(\inst$top.soc.cpu.gprf.mem[20][16] ),
    .B1(net1965),
    .B2(\inst$top.soc.cpu.gprf.mem[21][16] ),
    .Y(_06843_));
 sky130_fd_sc_hd__o21ai_0 _26146_ (.A1(_06839_),
    .A2(_06840_),
    .B1(_06843_),
    .Y(_06844_));
 sky130_fd_sc_hd__a221oi_1 _26147_ (.A1(_06838_),
    .A2(net2500),
    .B1(net1940),
    .B2(_06844_),
    .C1(net2447),
    .Y(_06845_));
 sky130_fd_sc_hd__nor2_1 _26148_ (.A(\inst$top.soc.cpu.gprf.mem[31][16] ),
    .B(net2488),
    .Y(_06846_));
 sky130_fd_sc_hd__o21ai_0 _26149_ (.A1(net2673),
    .A2(\inst$top.soc.cpu.gprf.mem[30][16] ),
    .B1(net2643),
    .Y(_06847_));
 sky130_fd_sc_hd__a221oi_1 _26150_ (.A1(net2525),
    .A2(\inst$top.soc.cpu.gprf.mem[28][16] ),
    .B1(net1965),
    .B2(\inst$top.soc.cpu.gprf.mem[29][16] ),
    .C1(net2459),
    .Y(_06848_));
 sky130_fd_sc_hd__o21ai_0 _26151_ (.A1(_06846_),
    .A2(_06847_),
    .B1(_06848_),
    .Y(_06849_));
 sky130_fd_sc_hd__nor2_1 _26152_ (.A(\inst$top.soc.cpu.gprf.mem[27][16] ),
    .B(net2488),
    .Y(_06850_));
 sky130_fd_sc_hd__o21ai_0 _26153_ (.A1(net2673),
    .A2(\inst$top.soc.cpu.gprf.mem[26][16] ),
    .B1(net2643),
    .Y(_06851_));
 sky130_fd_sc_hd__a221oi_1 _26154_ (.A1(net2525),
    .A2(\inst$top.soc.cpu.gprf.mem[24][16] ),
    .B1(net1965),
    .B2(\inst$top.soc.cpu.gprf.mem[25][16] ),
    .C1(net2613),
    .Y(_06852_));
 sky130_fd_sc_hd__o21ai_0 _26155_ (.A1(_06850_),
    .A2(_06851_),
    .B1(_06852_),
    .Y(_06853_));
 sky130_fd_sc_hd__nand3_1 _26156_ (.A(_06849_),
    .B(_06853_),
    .C(net2602),
    .Y(_06854_));
 sky130_fd_sc_hd__a32oi_1 _26157_ (.A1(_06822_),
    .A2(_06827_),
    .A3(_06832_),
    .B1(_06845_),
    .B2(_06854_),
    .Y(_00007_));
 sky130_fd_sc_hd__nor2_1 _26158_ (.A(\inst$top.soc.cpu.gprf.mem[31][17] ),
    .B(net2493),
    .Y(_06855_));
 sky130_fd_sc_hd__o21ai_0 _26159_ (.A1(net2683),
    .A2(\inst$top.soc.cpu.gprf.mem[30][17] ),
    .B1(net2649),
    .Y(_06856_));
 sky130_fd_sc_hd__a221oi_1 _26160_ (.A1(net2533),
    .A2(\inst$top.soc.cpu.gprf.mem[28][17] ),
    .B1(net1973),
    .B2(\inst$top.soc.cpu.gprf.mem[29][17] ),
    .C1(net2457),
    .Y(_06857_));
 sky130_fd_sc_hd__o21ai_0 _26161_ (.A1(_06855_),
    .A2(_06856_),
    .B1(_06857_),
    .Y(_06858_));
 sky130_fd_sc_hd__nor2_1 _26162_ (.A(\inst$top.soc.cpu.gprf.mem[27][17] ),
    .B(net2490),
    .Y(_06859_));
 sky130_fd_sc_hd__o21ai_0 _26163_ (.A1(net2682),
    .A2(\inst$top.soc.cpu.gprf.mem[26][17] ),
    .B1(net2646),
    .Y(_06860_));
 sky130_fd_sc_hd__a221oi_1 _26165_ (.A1(net2534),
    .A2(\inst$top.soc.cpu.gprf.mem[24][17] ),
    .B1(net1974),
    .B2(\inst$top.soc.cpu.gprf.mem[25][17] ),
    .C1(net2613),
    .Y(_06862_));
 sky130_fd_sc_hd__o21ai_0 _26166_ (.A1(_06859_),
    .A2(_06860_),
    .B1(_06862_),
    .Y(_06863_));
 sky130_fd_sc_hd__nand3_1 _26167_ (.A(_06858_),
    .B(_06863_),
    .C(net2604),
    .Y(_06864_));
 sky130_fd_sc_hd__nor2_1 _26168_ (.A(\inst$top.soc.cpu.gprf.mem[19][17] ),
    .B(net2490),
    .Y(_06865_));
 sky130_fd_sc_hd__o21ai_0 _26169_ (.A1(net2682),
    .A2(\inst$top.soc.cpu.gprf.mem[18][17] ),
    .B1(net2646),
    .Y(_06866_));
 sky130_fd_sc_hd__a22oi_1 _26170_ (.A1(net2534),
    .A2(\inst$top.soc.cpu.gprf.mem[16][17] ),
    .B1(net1974),
    .B2(\inst$top.soc.cpu.gprf.mem[17][17] ),
    .Y(_06867_));
 sky130_fd_sc_hd__o21ai_0 _26171_ (.A1(_06865_),
    .A2(_06866_),
    .B1(_06867_),
    .Y(_06868_));
 sky130_fd_sc_hd__a21oi_1 _26172_ (.A1(_06868_),
    .A2(net2502),
    .B1(net2447),
    .Y(_06869_));
 sky130_fd_sc_hd__nor2_1 _26173_ (.A(\inst$top.soc.cpu.gprf.mem[23][17] ),
    .B(net2493),
    .Y(_06870_));
 sky130_fd_sc_hd__o21ai_0 _26174_ (.A1(net2683),
    .A2(\inst$top.soc.cpu.gprf.mem[22][17] ),
    .B1(net2648),
    .Y(_06871_));
 sky130_fd_sc_hd__a22oi_1 _26175_ (.A1(net2533),
    .A2(\inst$top.soc.cpu.gprf.mem[20][17] ),
    .B1(net1973),
    .B2(\inst$top.soc.cpu.gprf.mem[21][17] ),
    .Y(_06872_));
 sky130_fd_sc_hd__o21ai_0 _26176_ (.A1(_06870_),
    .A2(_06871_),
    .B1(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__nand2_1 _26177_ (.A(_06873_),
    .B(net1939),
    .Y(_06874_));
 sky130_fd_sc_hd__nor2_1 _26178_ (.A(\inst$top.soc.cpu.gprf.mem[3][17] ),
    .B(net2490),
    .Y(_06875_));
 sky130_fd_sc_hd__o21ai_0 _26179_ (.A1(net2682),
    .A2(\inst$top.soc.cpu.gprf.mem[2][17] ),
    .B1(net2646),
    .Y(_06876_));
 sky130_fd_sc_hd__a22oi_1 _26180_ (.A1(net2531),
    .A2(\inst$top.soc.cpu.gprf.mem[0][17] ),
    .B1(net1971),
    .B2(\inst$top.soc.cpu.gprf.mem[1][17] ),
    .Y(_06877_));
 sky130_fd_sc_hd__o21ai_0 _26181_ (.A1(_06875_),
    .A2(_06876_),
    .B1(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__nor2_1 _26182_ (.A(\inst$top.soc.cpu.gprf.mem[7][17] ),
    .B(net2490),
    .Y(_06879_));
 sky130_fd_sc_hd__o21ai_0 _26183_ (.A1(net2682),
    .A2(\inst$top.soc.cpu.gprf.mem[6][17] ),
    .B1(net2646),
    .Y(_06880_));
 sky130_fd_sc_hd__a22oi_1 _26184_ (.A1(net2532),
    .A2(\inst$top.soc.cpu.gprf.mem[4][17] ),
    .B1(net1971),
    .B2(\inst$top.soc.cpu.gprf.mem[5][17] ),
    .Y(_06881_));
 sky130_fd_sc_hd__o21ai_0 _26185_ (.A1(_06879_),
    .A2(_06880_),
    .B1(_06881_),
    .Y(_06882_));
 sky130_fd_sc_hd__a221oi_1 _26186_ (.A1(_06878_),
    .A2(net2501),
    .B1(net1939),
    .B2(_06882_),
    .C1(net2593),
    .Y(_06883_));
 sky130_fd_sc_hd__nor2_1 _26187_ (.A(\inst$top.soc.cpu.gprf.mem[15][17] ),
    .B(net2491),
    .Y(_06884_));
 sky130_fd_sc_hd__o21ai_0 _26188_ (.A1(net2682),
    .A2(\inst$top.soc.cpu.gprf.mem[14][17] ),
    .B1(net2646),
    .Y(_06885_));
 sky130_fd_sc_hd__a221oi_1 _26189_ (.A1(net2534),
    .A2(\inst$top.soc.cpu.gprf.mem[12][17] ),
    .B1(net1974),
    .B2(\inst$top.soc.cpu.gprf.mem[13][17] ),
    .C1(net2458),
    .Y(_06886_));
 sky130_fd_sc_hd__o21ai_0 _26190_ (.A1(_06884_),
    .A2(_06885_),
    .B1(_06886_),
    .Y(_06887_));
 sky130_fd_sc_hd__nor2_1 _26191_ (.A(\inst$top.soc.cpu.gprf.mem[11][17] ),
    .B(net2491),
    .Y(_06888_));
 sky130_fd_sc_hd__o21ai_0 _26192_ (.A1(net2682),
    .A2(\inst$top.soc.cpu.gprf.mem[10][17] ),
    .B1(net2647),
    .Y(_06889_));
 sky130_fd_sc_hd__a221oi_1 _26193_ (.A1(net2534),
    .A2(\inst$top.soc.cpu.gprf.mem[8][17] ),
    .B1(net1974),
    .B2(\inst$top.soc.cpu.gprf.mem[9][17] ),
    .C1(net2614),
    .Y(_06890_));
 sky130_fd_sc_hd__o21ai_0 _26194_ (.A1(_06888_),
    .A2(_06889_),
    .B1(_06890_),
    .Y(_06891_));
 sky130_fd_sc_hd__nand3_1 _26195_ (.A(_06887_),
    .B(_06891_),
    .C(net2604),
    .Y(_06892_));
 sky130_fd_sc_hd__a32oi_1 _26196_ (.A1(_06864_),
    .A2(_06869_),
    .A3(_06874_),
    .B1(_06883_),
    .B2(_06892_),
    .Y(_00008_));
 sky130_fd_sc_hd__nor2_1 _26197_ (.A(\inst$top.soc.cpu.gprf.mem[11][18] ),
    .B(net2473),
    .Y(_06893_));
 sky130_fd_sc_hd__o21ai_0 _26198_ (.A1(net2661),
    .A2(\inst$top.soc.cpu.gprf.mem[10][18] ),
    .B1(net2627),
    .Y(_06894_));
 sky130_fd_sc_hd__a221oi_1 _26199_ (.A1(net2514),
    .A2(\inst$top.soc.cpu.gprf.mem[8][18] ),
    .B1(net1953),
    .B2(\inst$top.soc.cpu.gprf.mem[9][18] ),
    .C1(net2608),
    .Y(_06895_));
 sky130_fd_sc_hd__o21ai_0 _26200_ (.A1(_06893_),
    .A2(_06894_),
    .B1(_06895_),
    .Y(_06896_));
 sky130_fd_sc_hd__nor2_1 _26201_ (.A(\inst$top.soc.cpu.gprf.mem[15][18] ),
    .B(net2464),
    .Y(_06897_));
 sky130_fd_sc_hd__o21ai_0 _26204_ (.A1(net2656),
    .A2(\inst$top.soc.cpu.gprf.mem[14][18] ),
    .B1(net2619),
    .Y(_06900_));
 sky130_fd_sc_hd__a221oi_1 _26205_ (.A1(net2509),
    .A2(\inst$top.soc.cpu.gprf.mem[12][18] ),
    .B1(net1948),
    .B2(\inst$top.soc.cpu.gprf.mem[13][18] ),
    .C1(net2451),
    .Y(_06901_));
 sky130_fd_sc_hd__o21ai_0 _26206_ (.A1(_06897_),
    .A2(_06900_),
    .B1(_06901_),
    .Y(_06902_));
 sky130_fd_sc_hd__nand3_1 _26207_ (.A(_06896_),
    .B(_06902_),
    .C(net2600),
    .Y(_06903_));
 sky130_fd_sc_hd__nor2_1 _26208_ (.A(\inst$top.soc.cpu.gprf.mem[7][18] ),
    .B(net2468),
    .Y(_06904_));
 sky130_fd_sc_hd__o21ai_0 _26209_ (.A1(net2654),
    .A2(\inst$top.soc.cpu.gprf.mem[6][18] ),
    .B1(net2622),
    .Y(_06905_));
 sky130_fd_sc_hd__a22oi_1 _26210_ (.A1(net2511),
    .A2(\inst$top.soc.cpu.gprf.mem[4][18] ),
    .B1(net1950),
    .B2(\inst$top.soc.cpu.gprf.mem[5][18] ),
    .Y(_06906_));
 sky130_fd_sc_hd__o21ai_0 _26211_ (.A1(_06904_),
    .A2(_06905_),
    .B1(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__nand2_1 _26212_ (.A(_06907_),
    .B(net1934),
    .Y(_06908_));
 sky130_fd_sc_hd__nor2_1 _26213_ (.A(\inst$top.soc.cpu.gprf.mem[3][18] ),
    .B(net2464),
    .Y(_06909_));
 sky130_fd_sc_hd__o21ai_0 _26214_ (.A1(net2654),
    .A2(\inst$top.soc.cpu.gprf.mem[2][18] ),
    .B1(net2618),
    .Y(_06910_));
 sky130_fd_sc_hd__a22oi_1 _26216_ (.A1(net2507),
    .A2(\inst$top.soc.cpu.gprf.mem[0][18] ),
    .B1(net1946),
    .B2(\inst$top.soc.cpu.gprf.mem[1][18] ),
    .Y(_06912_));
 sky130_fd_sc_hd__o21ai_0 _26217_ (.A1(_06909_),
    .A2(_06910_),
    .B1(_06912_),
    .Y(_06913_));
 sky130_fd_sc_hd__a21oi_1 _26218_ (.A1(_06913_),
    .A2(net2504),
    .B1(net2592),
    .Y(_06914_));
 sky130_fd_sc_hd__nor2_1 _26219_ (.A(\inst$top.soc.cpu.gprf.mem[19][18] ),
    .B(net2464),
    .Y(_06915_));
 sky130_fd_sc_hd__o21ai_0 _26220_ (.A1(net2656),
    .A2(\inst$top.soc.cpu.gprf.mem[18][18] ),
    .B1(net2619),
    .Y(_06916_));
 sky130_fd_sc_hd__a22oi_1 _26221_ (.A1(net2509),
    .A2(\inst$top.soc.cpu.gprf.mem[16][18] ),
    .B1(net1948),
    .B2(\inst$top.soc.cpu.gprf.mem[17][18] ),
    .Y(_06917_));
 sky130_fd_sc_hd__o21ai_0 _26222_ (.A1(_06915_),
    .A2(_06916_),
    .B1(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__nor2_1 _26223_ (.A(\inst$top.soc.cpu.gprf.mem[23][18] ),
    .B(net2464),
    .Y(_06919_));
 sky130_fd_sc_hd__o21ai_0 _26224_ (.A1(net2654),
    .A2(\inst$top.soc.cpu.gprf.mem[22][18] ),
    .B1(net2618),
    .Y(_06920_));
 sky130_fd_sc_hd__a22oi_1 _26225_ (.A1(net2507),
    .A2(\inst$top.soc.cpu.gprf.mem[20][18] ),
    .B1(net1946),
    .B2(\inst$top.soc.cpu.gprf.mem[21][18] ),
    .Y(_06921_));
 sky130_fd_sc_hd__o21ai_0 _26226_ (.A1(_06919_),
    .A2(_06920_),
    .B1(_06921_),
    .Y(_06922_));
 sky130_fd_sc_hd__a221oi_1 _26227_ (.A1(net2507),
    .A2(\inst$top.soc.cpu.gprf.mem[28][18] ),
    .B1(net1946),
    .B2(\inst$top.soc.cpu.gprf.mem[29][18] ),
    .C1(net2451),
    .Y(_06923_));
 sky130_fd_sc_hd__nor2_1 _26228_ (.A(net2654),
    .B(\inst$top.soc.cpu.gprf.mem[30][18] ),
    .Y(_06924_));
 sky130_fd_sc_hd__nor2_1 _26229_ (.A(_20261_),
    .B(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__o21ai_0 _26230_ (.A1(net2462),
    .A2(\inst$top.soc.cpu.gprf.mem[31][18] ),
    .B1(_06925_),
    .Y(_06926_));
 sky130_fd_sc_hd__nor2_1 _26231_ (.A(\inst$top.soc.cpu.gprf.mem[27][18] ),
    .B(net2462),
    .Y(_06927_));
 sky130_fd_sc_hd__o21ai_0 _26232_ (.A1(net2653),
    .A2(\inst$top.soc.cpu.gprf.mem[26][18] ),
    .B1(net2617),
    .Y(_06928_));
 sky130_fd_sc_hd__nor2_1 _26233_ (.A(_06927_),
    .B(_06928_),
    .Y(_06929_));
 sky130_fd_sc_hd__inv_1 _26234_ (.A(\inst$top.soc.cpu.gprf.mem[24][18] ),
    .Y(_06930_));
 sky130_fd_sc_hd__o21ai_0 _26235_ (.A1(_06930_),
    .A2(_20236_),
    .B1(net2451),
    .Y(_06931_));
 sky130_fd_sc_hd__a211oi_1 _26236_ (.A1(\inst$top.soc.cpu.gprf.mem[25][18] ),
    .A2(net1946),
    .B1(_06929_),
    .C1(_06931_),
    .Y(_06932_));
 sky130_fd_sc_hd__a211oi_1 _26237_ (.A1(_06923_),
    .A2(_06926_),
    .B1(_06038_),
    .C1(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__a221oi_1 _26238_ (.A1(net2496),
    .A2(_06918_),
    .B1(net1943),
    .B2(_06922_),
    .C1(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__a32oi_1 _26239_ (.A1(_06903_),
    .A2(_06908_),
    .A3(_06914_),
    .B1(_06934_),
    .B2(net2592),
    .Y(_00009_));
 sky130_fd_sc_hd__nor2_1 _26240_ (.A(\inst$top.soc.cpu.gprf.mem[15][19] ),
    .B(net2491),
    .Y(_06935_));
 sky130_fd_sc_hd__o21ai_0 _26241_ (.A1(net2682),
    .A2(\inst$top.soc.cpu.gprf.mem[14][19] ),
    .B1(net2647),
    .Y(_06936_));
 sky130_fd_sc_hd__a221oi_1 _26243_ (.A1(net2534),
    .A2(\inst$top.soc.cpu.gprf.mem[12][19] ),
    .B1(net1974),
    .B2(\inst$top.soc.cpu.gprf.mem[13][19] ),
    .C1(net2457),
    .Y(_06938_));
 sky130_fd_sc_hd__o21ai_0 _26244_ (.A1(_06935_),
    .A2(_06936_),
    .B1(_06938_),
    .Y(_06939_));
 sky130_fd_sc_hd__nor2_1 _26245_ (.A(\inst$top.soc.cpu.gprf.mem[11][19] ),
    .B(net2490),
    .Y(_06940_));
 sky130_fd_sc_hd__o21ai_0 _26246_ (.A1(net2684),
    .A2(\inst$top.soc.cpu.gprf.mem[10][19] ),
    .B1(net2647),
    .Y(_06941_));
 sky130_fd_sc_hd__a221oi_1 _26247_ (.A1(net2534),
    .A2(\inst$top.soc.cpu.gprf.mem[8][19] ),
    .B1(net1974),
    .B2(\inst$top.soc.cpu.gprf.mem[9][19] ),
    .C1(net2613),
    .Y(_06942_));
 sky130_fd_sc_hd__o21ai_0 _26248_ (.A1(_06940_),
    .A2(_06941_),
    .B1(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__nand3_1 _26249_ (.A(_06939_),
    .B(_06943_),
    .C(net2604),
    .Y(_06944_));
 sky130_fd_sc_hd__nor2_1 _26250_ (.A(\inst$top.soc.cpu.gprf.mem[7][19] ),
    .B(net2490),
    .Y(_06945_));
 sky130_fd_sc_hd__o21ai_0 _26251_ (.A1(net2682),
    .A2(\inst$top.soc.cpu.gprf.mem[6][19] ),
    .B1(net2646),
    .Y(_06946_));
 sky130_fd_sc_hd__a22oi_1 _26252_ (.A1(net2531),
    .A2(\inst$top.soc.cpu.gprf.mem[4][19] ),
    .B1(net1971),
    .B2(\inst$top.soc.cpu.gprf.mem[5][19] ),
    .Y(_06947_));
 sky130_fd_sc_hd__o21ai_0 _26253_ (.A1(_06945_),
    .A2(_06946_),
    .B1(_06947_),
    .Y(_06948_));
 sky130_fd_sc_hd__nand2_1 _26254_ (.A(_06948_),
    .B(net1939),
    .Y(_06949_));
 sky130_fd_sc_hd__nor2_1 _26255_ (.A(\inst$top.soc.cpu.gprf.mem[3][19] ),
    .B(net2490),
    .Y(_06950_));
 sky130_fd_sc_hd__o21ai_0 _26256_ (.A1(net2680),
    .A2(\inst$top.soc.cpu.gprf.mem[2][19] ),
    .B1(net2646),
    .Y(_06951_));
 sky130_fd_sc_hd__a22oi_1 _26257_ (.A1(net2531),
    .A2(\inst$top.soc.cpu.gprf.mem[0][19] ),
    .B1(net1971),
    .B2(\inst$top.soc.cpu.gprf.mem[1][19] ),
    .Y(_06952_));
 sky130_fd_sc_hd__o21ai_0 _26258_ (.A1(_06950_),
    .A2(_06951_),
    .B1(_06952_),
    .Y(_06953_));
 sky130_fd_sc_hd__a21oi_1 _26259_ (.A1(_06953_),
    .A2(net2502),
    .B1(net2593),
    .Y(_06954_));
 sky130_fd_sc_hd__nor2_1 _26260_ (.A(\inst$top.soc.cpu.gprf.mem[23][19] ),
    .B(net2491),
    .Y(_06955_));
 sky130_fd_sc_hd__o21ai_0 _26261_ (.A1(net2684),
    .A2(\inst$top.soc.cpu.gprf.mem[22][19] ),
    .B1(net2647),
    .Y(_06956_));
 sky130_fd_sc_hd__a22oi_1 _26262_ (.A1(net2534),
    .A2(\inst$top.soc.cpu.gprf.mem[20][19] ),
    .B1(net1974),
    .B2(\inst$top.soc.cpu.gprf.mem[21][19] ),
    .Y(_06957_));
 sky130_fd_sc_hd__o21ai_0 _26263_ (.A1(_06955_),
    .A2(_06956_),
    .B1(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__nor2_1 _26264_ (.A(\inst$top.soc.cpu.gprf.mem[19][19] ),
    .B(net2491),
    .Y(_06959_));
 sky130_fd_sc_hd__o21ai_0 _26265_ (.A1(net2684),
    .A2(\inst$top.soc.cpu.gprf.mem[18][19] ),
    .B1(net2647),
    .Y(_06960_));
 sky130_fd_sc_hd__a22oi_1 _26266_ (.A1(net2534),
    .A2(\inst$top.soc.cpu.gprf.mem[16][19] ),
    .B1(net1974),
    .B2(\inst$top.soc.cpu.gprf.mem[17][19] ),
    .Y(_06961_));
 sky130_fd_sc_hd__o21ai_0 _26267_ (.A1(_06959_),
    .A2(_06960_),
    .B1(_06961_),
    .Y(_06962_));
 sky130_fd_sc_hd__a221oi_1 _26268_ (.A1(_06958_),
    .A2(net1939),
    .B1(net2502),
    .B2(_06962_),
    .C1(net2448),
    .Y(_06963_));
 sky130_fd_sc_hd__nor2_1 _26269_ (.A(\inst$top.soc.cpu.gprf.mem[31][19] ),
    .B(net2490),
    .Y(_06964_));
 sky130_fd_sc_hd__o21ai_0 _26270_ (.A1(net2682),
    .A2(\inst$top.soc.cpu.gprf.mem[30][19] ),
    .B1(net2646),
    .Y(_06965_));
 sky130_fd_sc_hd__a221oi_1 _26271_ (.A1(net2534),
    .A2(\inst$top.soc.cpu.gprf.mem[28][19] ),
    .B1(net1974),
    .B2(\inst$top.soc.cpu.gprf.mem[29][19] ),
    .C1(net2458),
    .Y(_06966_));
 sky130_fd_sc_hd__o21ai_0 _26272_ (.A1(_06964_),
    .A2(_06965_),
    .B1(_06966_),
    .Y(_06967_));
 sky130_fd_sc_hd__nor2_1 _26273_ (.A(\inst$top.soc.cpu.gprf.mem[27][19] ),
    .B(net2491),
    .Y(_06968_));
 sky130_fd_sc_hd__o21ai_0 _26274_ (.A1(net2682),
    .A2(\inst$top.soc.cpu.gprf.mem[26][19] ),
    .B1(net2647),
    .Y(_06969_));
 sky130_fd_sc_hd__a221oi_1 _26275_ (.A1(net2534),
    .A2(\inst$top.soc.cpu.gprf.mem[24][19] ),
    .B1(net1974),
    .B2(\inst$top.soc.cpu.gprf.mem[25][19] ),
    .C1(net2613),
    .Y(_06970_));
 sky130_fd_sc_hd__o21ai_0 _26276_ (.A1(_06968_),
    .A2(_06969_),
    .B1(_06970_),
    .Y(_06971_));
 sky130_fd_sc_hd__nand3_1 _26277_ (.A(_06967_),
    .B(_06971_),
    .C(net2604),
    .Y(_06972_));
 sky130_fd_sc_hd__a32oi_1 _26278_ (.A1(_06944_),
    .A2(_06949_),
    .A3(_06954_),
    .B1(_06963_),
    .B2(_06972_),
    .Y(_00010_));
 sky130_fd_sc_hd__nor2_1 _26279_ (.A(\inst$top.soc.cpu.gprf.mem[11][20] ),
    .B(net2475),
    .Y(_06973_));
 sky130_fd_sc_hd__o21ai_0 _26280_ (.A1(net2663),
    .A2(\inst$top.soc.cpu.gprf.mem[10][20] ),
    .B1(net2629),
    .Y(_06974_));
 sky130_fd_sc_hd__a221oi_1 _26281_ (.A1(net2522),
    .A2(\inst$top.soc.cpu.gprf.mem[8][20] ),
    .B1(net1962),
    .B2(\inst$top.soc.cpu.gprf.mem[9][20] ),
    .C1(net2609),
    .Y(_06975_));
 sky130_fd_sc_hd__o21ai_0 _26282_ (.A1(_06973_),
    .A2(_06974_),
    .B1(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__nor2_1 _26284_ (.A(\inst$top.soc.cpu.gprf.mem[15][20] ),
    .B(net2476),
    .Y(_06978_));
 sky130_fd_sc_hd__o21ai_0 _26285_ (.A1(net2670),
    .A2(\inst$top.soc.cpu.gprf.mem[14][20] ),
    .B1(net2630),
    .Y(_06979_));
 sky130_fd_sc_hd__a221oi_1 _26286_ (.A1(net2522),
    .A2(\inst$top.soc.cpu.gprf.mem[12][20] ),
    .B1(net1962),
    .B2(\inst$top.soc.cpu.gprf.mem[13][20] ),
    .C1(net2455),
    .Y(_06980_));
 sky130_fd_sc_hd__o21ai_0 _26287_ (.A1(_06978_),
    .A2(_06979_),
    .B1(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__nand3_1 _26289_ (.A(_06976_),
    .B(_06981_),
    .C(net2599),
    .Y(_06983_));
 sky130_fd_sc_hd__nor2_1 _26290_ (.A(\inst$top.soc.cpu.gprf.mem[7][20] ),
    .B(net2476),
    .Y(_06984_));
 sky130_fd_sc_hd__o21ai_0 _26291_ (.A1(net2670),
    .A2(\inst$top.soc.cpu.gprf.mem[6][20] ),
    .B1(net2630),
    .Y(_06985_));
 sky130_fd_sc_hd__a22oi_1 _26292_ (.A1(net2523),
    .A2(\inst$top.soc.cpu.gprf.mem[4][20] ),
    .B1(net1962),
    .B2(\inst$top.soc.cpu.gprf.mem[5][20] ),
    .Y(_06986_));
 sky130_fd_sc_hd__o21ai_0 _26293_ (.A1(_06984_),
    .A2(_06985_),
    .B1(_06986_),
    .Y(_06987_));
 sky130_fd_sc_hd__nand2_1 _26294_ (.A(_06987_),
    .B(net1936),
    .Y(_06988_));
 sky130_fd_sc_hd__nor2_1 _26295_ (.A(\inst$top.soc.cpu.gprf.mem[3][20] ),
    .B(net2475),
    .Y(_06989_));
 sky130_fd_sc_hd__o21ai_0 _26296_ (.A1(net2670),
    .A2(\inst$top.soc.cpu.gprf.mem[2][20] ),
    .B1(net2630),
    .Y(_06990_));
 sky130_fd_sc_hd__a22oi_1 _26297_ (.A1(net2522),
    .A2(\inst$top.soc.cpu.gprf.mem[0][20] ),
    .B1(net1962),
    .B2(\inst$top.soc.cpu.gprf.mem[1][20] ),
    .Y(_06991_));
 sky130_fd_sc_hd__o21ai_0 _26298_ (.A1(_06989_),
    .A2(_06990_),
    .B1(_06991_),
    .Y(_06992_));
 sky130_fd_sc_hd__a21oi_1 _26299_ (.A1(_06992_),
    .A2(net2498),
    .B1(net2594),
    .Y(_06993_));
 sky130_fd_sc_hd__nor2_1 _26300_ (.A(\inst$top.soc.cpu.gprf.mem[19][20] ),
    .B(net2475),
    .Y(_06994_));
 sky130_fd_sc_hd__o21ai_0 _26301_ (.A1(net2663),
    .A2(\inst$top.soc.cpu.gprf.mem[18][20] ),
    .B1(net2629),
    .Y(_06995_));
 sky130_fd_sc_hd__a22oi_1 _26302_ (.A1(net2522),
    .A2(\inst$top.soc.cpu.gprf.mem[16][20] ),
    .B1(net1962),
    .B2(\inst$top.soc.cpu.gprf.mem[17][20] ),
    .Y(_06996_));
 sky130_fd_sc_hd__o21ai_0 _26303_ (.A1(_06994_),
    .A2(_06995_),
    .B1(_06996_),
    .Y(_06997_));
 sky130_fd_sc_hd__nor2_1 _26304_ (.A(\inst$top.soc.cpu.gprf.mem[23][20] ),
    .B(net2476),
    .Y(_06998_));
 sky130_fd_sc_hd__o21ai_0 _26305_ (.A1(net2670),
    .A2(\inst$top.soc.cpu.gprf.mem[22][20] ),
    .B1(net2630),
    .Y(_06999_));
 sky130_fd_sc_hd__a22oi_1 _26306_ (.A1(net2522),
    .A2(\inst$top.soc.cpu.gprf.mem[20][20] ),
    .B1(net1962),
    .B2(\inst$top.soc.cpu.gprf.mem[21][20] ),
    .Y(_07000_));
 sky130_fd_sc_hd__o21ai_0 _26307_ (.A1(_06998_),
    .A2(_06999_),
    .B1(_07000_),
    .Y(_07001_));
 sky130_fd_sc_hd__a221oi_1 _26308_ (.A1(_06997_),
    .A2(net2498),
    .B1(net1936),
    .B2(_07001_),
    .C1(net2449),
    .Y(_07002_));
 sky130_fd_sc_hd__nor2_1 _26309_ (.A(\inst$top.soc.cpu.gprf.mem[31][20] ),
    .B(net2475),
    .Y(_07003_));
 sky130_fd_sc_hd__o21ai_0 _26310_ (.A1(net2670),
    .A2(\inst$top.soc.cpu.gprf.mem[30][20] ),
    .B1(net2630),
    .Y(_07004_));
 sky130_fd_sc_hd__a221oi_1 _26311_ (.A1(net2522),
    .A2(\inst$top.soc.cpu.gprf.mem[28][20] ),
    .B1(net1962),
    .B2(\inst$top.soc.cpu.gprf.mem[29][20] ),
    .C1(net2455),
    .Y(_07005_));
 sky130_fd_sc_hd__o21ai_0 _26312_ (.A1(_07003_),
    .A2(_07004_),
    .B1(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__nor2_1 _26313_ (.A(\inst$top.soc.cpu.gprf.mem[27][20] ),
    .B(net2476),
    .Y(_07007_));
 sky130_fd_sc_hd__o21ai_0 _26314_ (.A1(net2670),
    .A2(\inst$top.soc.cpu.gprf.mem[26][20] ),
    .B1(net2630),
    .Y(_07008_));
 sky130_fd_sc_hd__a221oi_1 _26315_ (.A1(net2523),
    .A2(\inst$top.soc.cpu.gprf.mem[24][20] ),
    .B1(net1963),
    .B2(\inst$top.soc.cpu.gprf.mem[25][20] ),
    .C1(net2609),
    .Y(_07009_));
 sky130_fd_sc_hd__o21ai_0 _26316_ (.A1(_07007_),
    .A2(_07008_),
    .B1(_07009_),
    .Y(_07010_));
 sky130_fd_sc_hd__nand3_1 _26317_ (.A(_07006_),
    .B(_07010_),
    .C(net2598),
    .Y(_07011_));
 sky130_fd_sc_hd__a32oi_1 _26318_ (.A1(_06983_),
    .A2(_06988_),
    .A3(_06993_),
    .B1(_07002_),
    .B2(_07011_),
    .Y(_00012_));
 sky130_fd_sc_hd__nor2_1 _26319_ (.A(\inst$top.soc.cpu.gprf.mem[15][21] ),
    .B(net2490),
    .Y(_07012_));
 sky130_fd_sc_hd__o21ai_0 _26320_ (.A1(net2680),
    .A2(\inst$top.soc.cpu.gprf.mem[14][21] ),
    .B1(net2646),
    .Y(_07013_));
 sky130_fd_sc_hd__a221oi_1 _26321_ (.A1(net2531),
    .A2(\inst$top.soc.cpu.gprf.mem[12][21] ),
    .B1(net1971),
    .B2(\inst$top.soc.cpu.gprf.mem[13][21] ),
    .C1(net2457),
    .Y(_07014_));
 sky130_fd_sc_hd__o21ai_0 _26322_ (.A1(_07012_),
    .A2(_07013_),
    .B1(_07014_),
    .Y(_07015_));
 sky130_fd_sc_hd__nor2_1 _26323_ (.A(\inst$top.soc.cpu.gprf.mem[11][21] ),
    .B(net2489),
    .Y(_07016_));
 sky130_fd_sc_hd__o21ai_0 _26324_ (.A1(net2680),
    .A2(\inst$top.soc.cpu.gprf.mem[10][21] ),
    .B1(net2645),
    .Y(_07017_));
 sky130_fd_sc_hd__a221oi_1 _26325_ (.A1(net2531),
    .A2(\inst$top.soc.cpu.gprf.mem[8][21] ),
    .B1(net1971),
    .B2(\inst$top.soc.cpu.gprf.mem[9][21] ),
    .C1(net2613),
    .Y(_07018_));
 sky130_fd_sc_hd__o21ai_0 _26326_ (.A1(_07016_),
    .A2(_07017_),
    .B1(_07018_),
    .Y(_07019_));
 sky130_fd_sc_hd__nand3_1 _26327_ (.A(_07015_),
    .B(_07019_),
    .C(net2604),
    .Y(_07020_));
 sky130_fd_sc_hd__nor2_1 _26328_ (.A(\inst$top.soc.cpu.gprf.mem[7][21] ),
    .B(net2487),
    .Y(_07021_));
 sky130_fd_sc_hd__o21ai_0 _26329_ (.A1(net2680),
    .A2(\inst$top.soc.cpu.gprf.mem[6][21] ),
    .B1(net2642),
    .Y(_07022_));
 sky130_fd_sc_hd__a22oi_1 _26330_ (.A1(net2531),
    .A2(\inst$top.soc.cpu.gprf.mem[4][21] ),
    .B1(net1971),
    .B2(\inst$top.soc.cpu.gprf.mem[5][21] ),
    .Y(_07023_));
 sky130_fd_sc_hd__o21ai_0 _26331_ (.A1(_07021_),
    .A2(_07022_),
    .B1(_07023_),
    .Y(_07024_));
 sky130_fd_sc_hd__nand2_1 _26332_ (.A(_07024_),
    .B(net1940),
    .Y(_07025_));
 sky130_fd_sc_hd__nor2_1 _26333_ (.A(\inst$top.soc.cpu.gprf.mem[3][21] ),
    .B(net2489),
    .Y(_07026_));
 sky130_fd_sc_hd__o21ai_0 _26334_ (.A1(net2680),
    .A2(\inst$top.soc.cpu.gprf.mem[2][21] ),
    .B1(net2642),
    .Y(_07027_));
 sky130_fd_sc_hd__a22oi_1 _26335_ (.A1(net2531),
    .A2(\inst$top.soc.cpu.gprf.mem[0][21] ),
    .B1(net1971),
    .B2(\inst$top.soc.cpu.gprf.mem[1][21] ),
    .Y(_07028_));
 sky130_fd_sc_hd__o21ai_0 _26336_ (.A1(_07026_),
    .A2(_07027_),
    .B1(_07028_),
    .Y(_07029_));
 sky130_fd_sc_hd__a21oi_1 _26337_ (.A1(_07029_),
    .A2(net2503),
    .B1(net2593),
    .Y(_07030_));
 sky130_fd_sc_hd__nor2_1 _26338_ (.A(\inst$top.soc.cpu.gprf.mem[23][21] ),
    .B(net2489),
    .Y(_07031_));
 sky130_fd_sc_hd__o21ai_0 _26339_ (.A1(net2681),
    .A2(\inst$top.soc.cpu.gprf.mem[22][21] ),
    .B1(net2644),
    .Y(_07032_));
 sky130_fd_sc_hd__a22oi_1 _26340_ (.A1(net2531),
    .A2(\inst$top.soc.cpu.gprf.mem[20][21] ),
    .B1(net1971),
    .B2(\inst$top.soc.cpu.gprf.mem[21][21] ),
    .Y(_07033_));
 sky130_fd_sc_hd__o21ai_0 _26341_ (.A1(_07031_),
    .A2(_07032_),
    .B1(_07033_),
    .Y(_07034_));
 sky130_fd_sc_hd__nor2_1 _26342_ (.A(\inst$top.soc.cpu.gprf.mem[19][21] ),
    .B(net2489),
    .Y(_07035_));
 sky130_fd_sc_hd__o21ai_0 _26343_ (.A1(net2672),
    .A2(\inst$top.soc.cpu.gprf.mem[18][21] ),
    .B1(net2642),
    .Y(_07036_));
 sky130_fd_sc_hd__a22oi_1 _26344_ (.A1(net2524),
    .A2(\inst$top.soc.cpu.gprf.mem[16][21] ),
    .B1(net1964),
    .B2(\inst$top.soc.cpu.gprf.mem[17][21] ),
    .Y(_07037_));
 sky130_fd_sc_hd__o21ai_0 _26345_ (.A1(_07035_),
    .A2(_07036_),
    .B1(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__a221oi_1 _26346_ (.A1(_07034_),
    .A2(net1940),
    .B1(net2503),
    .B2(_07038_),
    .C1(net2447),
    .Y(_07039_));
 sky130_fd_sc_hd__nor2_1 _26347_ (.A(\inst$top.soc.cpu.gprf.mem[31][21] ),
    .B(net2487),
    .Y(_07040_));
 sky130_fd_sc_hd__o21ai_0 _26350_ (.A1(net2680),
    .A2(\inst$top.soc.cpu.gprf.mem[30][21] ),
    .B1(net2645),
    .Y(_07043_));
 sky130_fd_sc_hd__a221oi_1 _26352_ (.A1(net2531),
    .A2(\inst$top.soc.cpu.gprf.mem[28][21] ),
    .B1(net1972),
    .B2(\inst$top.soc.cpu.gprf.mem[29][21] ),
    .C1(net2458),
    .Y(_07045_));
 sky130_fd_sc_hd__o21ai_0 _26353_ (.A1(_07040_),
    .A2(_07043_),
    .B1(_07045_),
    .Y(_07046_));
 sky130_fd_sc_hd__nor2_1 _26354_ (.A(\inst$top.soc.cpu.gprf.mem[27][21] ),
    .B(net2490),
    .Y(_07047_));
 sky130_fd_sc_hd__o21ai_0 _26355_ (.A1(net2680),
    .A2(\inst$top.soc.cpu.gprf.mem[26][21] ),
    .B1(net2646),
    .Y(_07048_));
 sky130_fd_sc_hd__a221oi_1 _26357_ (.A1(net2531),
    .A2(\inst$top.soc.cpu.gprf.mem[24][21] ),
    .B1(net1971),
    .B2(\inst$top.soc.cpu.gprf.mem[25][21] ),
    .C1(net2614),
    .Y(_07050_));
 sky130_fd_sc_hd__o21ai_0 _26358_ (.A1(_07047_),
    .A2(_07048_),
    .B1(_07050_),
    .Y(_07051_));
 sky130_fd_sc_hd__nand3_1 _26360_ (.A(_07046_),
    .B(_07051_),
    .C(net2605),
    .Y(_07053_));
 sky130_fd_sc_hd__a32oi_1 _26361_ (.A1(_07020_),
    .A2(_07025_),
    .A3(_07030_),
    .B1(_07039_),
    .B2(_07053_),
    .Y(_00013_));
 sky130_fd_sc_hd__nor2_1 _26362_ (.A(\inst$top.soc.cpu.gprf.mem[11][22] ),
    .B(net2464),
    .Y(_07054_));
 sky130_fd_sc_hd__o21ai_0 _26365_ (.A1(net2656),
    .A2(\inst$top.soc.cpu.gprf.mem[10][22] ),
    .B1(net2619),
    .Y(_07057_));
 sky130_fd_sc_hd__a221oi_1 _26367_ (.A1(net2509),
    .A2(\inst$top.soc.cpu.gprf.mem[8][22] ),
    .B1(net1948),
    .B2(\inst$top.soc.cpu.gprf.mem[9][22] ),
    .C1(net2607),
    .Y(_07059_));
 sky130_fd_sc_hd__o21ai_0 _26368_ (.A1(_07054_),
    .A2(_07057_),
    .B1(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__nor2_1 _26369_ (.A(\inst$top.soc.cpu.gprf.mem[15][22] ),
    .B(net2464),
    .Y(_07061_));
 sky130_fd_sc_hd__o21ai_0 _26370_ (.A1(net2656),
    .A2(\inst$top.soc.cpu.gprf.mem[14][22] ),
    .B1(net2619),
    .Y(_07062_));
 sky130_fd_sc_hd__a221oi_1 _26371_ (.A1(net2509),
    .A2(\inst$top.soc.cpu.gprf.mem[12][22] ),
    .B1(net1948),
    .B2(\inst$top.soc.cpu.gprf.mem[13][22] ),
    .C1(net2451),
    .Y(_07063_));
 sky130_fd_sc_hd__o21ai_0 _26372_ (.A1(_07061_),
    .A2(_07062_),
    .B1(_07063_),
    .Y(_07064_));
 sky130_fd_sc_hd__nand3_1 _26373_ (.A(_07060_),
    .B(_07064_),
    .C(net2600),
    .Y(_07065_));
 sky130_fd_sc_hd__nor2_1 _26374_ (.A(\inst$top.soc.cpu.gprf.mem[7][22] ),
    .B(net2473),
    .Y(_07066_));
 sky130_fd_sc_hd__o21ai_0 _26375_ (.A1(net2656),
    .A2(\inst$top.soc.cpu.gprf.mem[6][22] ),
    .B1(net2628),
    .Y(_07067_));
 sky130_fd_sc_hd__a22oi_1 _26376_ (.A1(net2509),
    .A2(\inst$top.soc.cpu.gprf.mem[4][22] ),
    .B1(net1953),
    .B2(\inst$top.soc.cpu.gprf.mem[5][22] ),
    .Y(_07068_));
 sky130_fd_sc_hd__o21ai_0 _26377_ (.A1(_07066_),
    .A2(_07067_),
    .B1(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__nand2_1 _26378_ (.A(_07069_),
    .B(net1936),
    .Y(_07070_));
 sky130_fd_sc_hd__nor2_1 _26379_ (.A(\inst$top.soc.cpu.gprf.mem[3][22] ),
    .B(net2473),
    .Y(_07071_));
 sky130_fd_sc_hd__o21ai_0 _26380_ (.A1(net2656),
    .A2(\inst$top.soc.cpu.gprf.mem[2][22] ),
    .B1(net2627),
    .Y(_07072_));
 sky130_fd_sc_hd__a22oi_1 _26381_ (.A1(net2509),
    .A2(\inst$top.soc.cpu.gprf.mem[0][22] ),
    .B1(net1953),
    .B2(\inst$top.soc.cpu.gprf.mem[1][22] ),
    .Y(_07073_));
 sky130_fd_sc_hd__o21ai_0 _26382_ (.A1(_07071_),
    .A2(_07072_),
    .B1(_07073_),
    .Y(_07074_));
 sky130_fd_sc_hd__a21oi_1 _26383_ (.A1(_07074_),
    .A2(net2499),
    .B1(net2592),
    .Y(_07075_));
 sky130_fd_sc_hd__nor2_1 _26384_ (.A(\inst$top.soc.cpu.gprf.mem[23][22] ),
    .B(net2473),
    .Y(_07076_));
 sky130_fd_sc_hd__o21ai_0 _26385_ (.A1(net2661),
    .A2(\inst$top.soc.cpu.gprf.mem[22][22] ),
    .B1(net2627),
    .Y(_07077_));
 sky130_fd_sc_hd__a22oi_1 _26386_ (.A1(net2514),
    .A2(\inst$top.soc.cpu.gprf.mem[20][22] ),
    .B1(net1953),
    .B2(\inst$top.soc.cpu.gprf.mem[21][22] ),
    .Y(_07078_));
 sky130_fd_sc_hd__o21ai_0 _26387_ (.A1(_07076_),
    .A2(_07077_),
    .B1(_07078_),
    .Y(_07079_));
 sky130_fd_sc_hd__nor2_1 _26388_ (.A(\inst$top.soc.cpu.gprf.mem[19][22] ),
    .B(net2473),
    .Y(_07080_));
 sky130_fd_sc_hd__o21ai_0 _26389_ (.A1(net2661),
    .A2(\inst$top.soc.cpu.gprf.mem[18][22] ),
    .B1(net2627),
    .Y(_07081_));
 sky130_fd_sc_hd__a22oi_1 _26390_ (.A1(net2514),
    .A2(\inst$top.soc.cpu.gprf.mem[16][22] ),
    .B1(net1953),
    .B2(\inst$top.soc.cpu.gprf.mem[17][22] ),
    .Y(_07082_));
 sky130_fd_sc_hd__o21ai_0 _26391_ (.A1(_07080_),
    .A2(_07081_),
    .B1(_07082_),
    .Y(_07083_));
 sky130_fd_sc_hd__a221oi_1 _26392_ (.A1(_07079_),
    .A2(net1934),
    .B1(net2499),
    .B2(_07083_),
    .C1(net2446),
    .Y(_07084_));
 sky130_fd_sc_hd__nor2_1 _26393_ (.A(\inst$top.soc.cpu.gprf.mem[31][22] ),
    .B(net2473),
    .Y(_07085_));
 sky130_fd_sc_hd__o21ai_0 _26394_ (.A1(net2661),
    .A2(\inst$top.soc.cpu.gprf.mem[30][22] ),
    .B1(net2627),
    .Y(_07086_));
 sky130_fd_sc_hd__a221oi_1 _26395_ (.A1(net2514),
    .A2(\inst$top.soc.cpu.gprf.mem[28][22] ),
    .B1(net1953),
    .B2(\inst$top.soc.cpu.gprf.mem[29][22] ),
    .C1(net2452),
    .Y(_07087_));
 sky130_fd_sc_hd__o21ai_0 _26396_ (.A1(_07085_),
    .A2(_07086_),
    .B1(_07087_),
    .Y(_07088_));
 sky130_fd_sc_hd__nor2_1 _26397_ (.A(\inst$top.soc.cpu.gprf.mem[27][22] ),
    .B(net2464),
    .Y(_07089_));
 sky130_fd_sc_hd__o21ai_0 _26398_ (.A1(net2656),
    .A2(\inst$top.soc.cpu.gprf.mem[26][22] ),
    .B1(net2627),
    .Y(_07090_));
 sky130_fd_sc_hd__a221oi_1 _26399_ (.A1(net2509),
    .A2(\inst$top.soc.cpu.gprf.mem[24][22] ),
    .B1(net1953),
    .B2(\inst$top.soc.cpu.gprf.mem[25][22] ),
    .C1(net2608),
    .Y(_07091_));
 sky130_fd_sc_hd__o21ai_0 _26400_ (.A1(_07089_),
    .A2(_07090_),
    .B1(_07091_),
    .Y(_07092_));
 sky130_fd_sc_hd__nand3_1 _26401_ (.A(_07088_),
    .B(_07092_),
    .C(net2600),
    .Y(_07093_));
 sky130_fd_sc_hd__a32oi_1 _26402_ (.A1(_07065_),
    .A2(_07070_),
    .A3(_07075_),
    .B1(_07084_),
    .B2(_07093_),
    .Y(_00014_));
 sky130_fd_sc_hd__nor2_1 _26403_ (.A(\inst$top.soc.cpu.gprf.mem[31][23] ),
    .B(net2475),
    .Y(_07094_));
 sky130_fd_sc_hd__o21ai_0 _26404_ (.A1(net2663),
    .A2(\inst$top.soc.cpu.gprf.mem[30][23] ),
    .B1(net2629),
    .Y(_07095_));
 sky130_fd_sc_hd__a221oi_1 _26405_ (.A1(net2516),
    .A2(\inst$top.soc.cpu.gprf.mem[28][23] ),
    .B1(net1955),
    .B2(\inst$top.soc.cpu.gprf.mem[29][23] ),
    .C1(net2453),
    .Y(_07096_));
 sky130_fd_sc_hd__o21ai_0 _26406_ (.A1(_07094_),
    .A2(_07095_),
    .B1(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__nor2_1 _26407_ (.A(\inst$top.soc.cpu.gprf.mem[27][23] ),
    .B(net2475),
    .Y(_07098_));
 sky130_fd_sc_hd__o21ai_0 _26408_ (.A1(net2663),
    .A2(\inst$top.soc.cpu.gprf.mem[26][23] ),
    .B1(net2629),
    .Y(_07099_));
 sky130_fd_sc_hd__a221oi_1 _26409_ (.A1(net2516),
    .A2(\inst$top.soc.cpu.gprf.mem[24][23] ),
    .B1(net1955),
    .B2(\inst$top.soc.cpu.gprf.mem[25][23] ),
    .C1(net2609),
    .Y(_07100_));
 sky130_fd_sc_hd__o21ai_0 _26410_ (.A1(_07098_),
    .A2(_07099_),
    .B1(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__nand3_1 _26411_ (.A(_07097_),
    .B(_07101_),
    .C(net2599),
    .Y(_07102_));
 sky130_fd_sc_hd__nor2_1 _26412_ (.A(\inst$top.soc.cpu.gprf.mem[19][23] ),
    .B(net2478),
    .Y(_07103_));
 sky130_fd_sc_hd__o21ai_0 _26413_ (.A1(net2662),
    .A2(\inst$top.soc.cpu.gprf.mem[18][23] ),
    .B1(net2628),
    .Y(_07104_));
 sky130_fd_sc_hd__a22oi_1 _26414_ (.A1(net2516),
    .A2(\inst$top.soc.cpu.gprf.mem[16][23] ),
    .B1(net1954),
    .B2(\inst$top.soc.cpu.gprf.mem[17][23] ),
    .Y(_07105_));
 sky130_fd_sc_hd__o21ai_0 _26415_ (.A1(_07103_),
    .A2(_07104_),
    .B1(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__nand2_1 _26416_ (.A(_07106_),
    .B(net2498),
    .Y(_07107_));
 sky130_fd_sc_hd__nor2_1 _26417_ (.A(\inst$top.soc.cpu.gprf.mem[23][23] ),
    .B(net2475),
    .Y(_07108_));
 sky130_fd_sc_hd__o21ai_0 _26418_ (.A1(net2663),
    .A2(\inst$top.soc.cpu.gprf.mem[22][23] ),
    .B1(net2629),
    .Y(_07109_));
 sky130_fd_sc_hd__a22oi_1 _26419_ (.A1(net2516),
    .A2(\inst$top.soc.cpu.gprf.mem[20][23] ),
    .B1(net1955),
    .B2(\inst$top.soc.cpu.gprf.mem[21][23] ),
    .Y(_07110_));
 sky130_fd_sc_hd__o21ai_0 _26420_ (.A1(_07108_),
    .A2(_07109_),
    .B1(_07110_),
    .Y(_07111_));
 sky130_fd_sc_hd__a21oi_1 _26421_ (.A1(_07111_),
    .A2(net1936),
    .B1(net2446),
    .Y(_07112_));
 sky130_fd_sc_hd__nor2_1 _26422_ (.A(\inst$top.soc.cpu.gprf.mem[3][23] ),
    .B(net2475),
    .Y(_07113_));
 sky130_fd_sc_hd__o21ai_0 _26423_ (.A1(net2663),
    .A2(\inst$top.soc.cpu.gprf.mem[2][23] ),
    .B1(net2629),
    .Y(_07114_));
 sky130_fd_sc_hd__a22oi_1 _26424_ (.A1(net2516),
    .A2(\inst$top.soc.cpu.gprf.mem[0][23] ),
    .B1(net1955),
    .B2(\inst$top.soc.cpu.gprf.mem[1][23] ),
    .Y(_07115_));
 sky130_fd_sc_hd__o21ai_0 _26425_ (.A1(_07113_),
    .A2(_07114_),
    .B1(_07115_),
    .Y(_07116_));
 sky130_fd_sc_hd__nor2_1 _26426_ (.A(\inst$top.soc.cpu.gprf.mem[7][23] ),
    .B(net2475),
    .Y(_07117_));
 sky130_fd_sc_hd__o21ai_0 _26427_ (.A1(net2663),
    .A2(\inst$top.soc.cpu.gprf.mem[6][23] ),
    .B1(net2629),
    .Y(_07118_));
 sky130_fd_sc_hd__a22oi_1 _26428_ (.A1(net2516),
    .A2(\inst$top.soc.cpu.gprf.mem[4][23] ),
    .B1(net1955),
    .B2(\inst$top.soc.cpu.gprf.mem[5][23] ),
    .Y(_07119_));
 sky130_fd_sc_hd__o21ai_0 _26429_ (.A1(_07117_),
    .A2(_07118_),
    .B1(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__a221oi_1 _26430_ (.A1(_07116_),
    .A2(net2498),
    .B1(net1935),
    .B2(_07120_),
    .C1(net2592),
    .Y(_07121_));
 sky130_fd_sc_hd__nor2_1 _26431_ (.A(\inst$top.soc.cpu.gprf.mem[15][23] ),
    .B(net2474),
    .Y(_07122_));
 sky130_fd_sc_hd__o21ai_0 _26432_ (.A1(net2663),
    .A2(\inst$top.soc.cpu.gprf.mem[14][23] ),
    .B1(net2632),
    .Y(_07123_));
 sky130_fd_sc_hd__a221oi_1 _26433_ (.A1(net2515),
    .A2(\inst$top.soc.cpu.gprf.mem[12][23] ),
    .B1(net1955),
    .B2(\inst$top.soc.cpu.gprf.mem[13][23] ),
    .C1(net2453),
    .Y(_07124_));
 sky130_fd_sc_hd__o21ai_0 _26434_ (.A1(_07122_),
    .A2(_07123_),
    .B1(_07124_),
    .Y(_07125_));
 sky130_fd_sc_hd__nor2_1 _26435_ (.A(\inst$top.soc.cpu.gprf.mem[11][23] ),
    .B(net2475),
    .Y(_07126_));
 sky130_fd_sc_hd__o21ai_0 _26436_ (.A1(net2662),
    .A2(\inst$top.soc.cpu.gprf.mem[10][23] ),
    .B1(net2629),
    .Y(_07127_));
 sky130_fd_sc_hd__a221oi_1 _26437_ (.A1(net2515),
    .A2(\inst$top.soc.cpu.gprf.mem[8][23] ),
    .B1(net1954),
    .B2(\inst$top.soc.cpu.gprf.mem[9][23] ),
    .C1(net2609),
    .Y(_07128_));
 sky130_fd_sc_hd__o21ai_0 _26438_ (.A1(_07126_),
    .A2(_07127_),
    .B1(_07128_),
    .Y(_07129_));
 sky130_fd_sc_hd__nand3_1 _26439_ (.A(_07125_),
    .B(_07129_),
    .C(net2599),
    .Y(_07130_));
 sky130_fd_sc_hd__a32oi_1 _26440_ (.A1(_07102_),
    .A2(_07107_),
    .A3(_07112_),
    .B1(_07121_),
    .B2(_07130_),
    .Y(_00015_));
 sky130_fd_sc_hd__nor2_1 _26441_ (.A(\inst$top.soc.cpu.gprf.mem[11][24] ),
    .B(net2492),
    .Y(_07131_));
 sky130_fd_sc_hd__o21ai_0 _26442_ (.A1(net2684),
    .A2(\inst$top.soc.cpu.gprf.mem[10][24] ),
    .B1(net2649),
    .Y(_07132_));
 sky130_fd_sc_hd__a221oi_1 _26443_ (.A1(net2535),
    .A2(\inst$top.soc.cpu.gprf.mem[8][24] ),
    .B1(net1975),
    .B2(\inst$top.soc.cpu.gprf.mem[9][24] ),
    .C1(net2613),
    .Y(_07133_));
 sky130_fd_sc_hd__o21ai_0 _26444_ (.A1(_07131_),
    .A2(_07132_),
    .B1(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__nor2_1 _26445_ (.A(\inst$top.soc.cpu.gprf.mem[15][24] ),
    .B(net2493),
    .Y(_07135_));
 sky130_fd_sc_hd__o21ai_0 _26446_ (.A1(net2684),
    .A2(\inst$top.soc.cpu.gprf.mem[14][24] ),
    .B1(net2649),
    .Y(_07136_));
 sky130_fd_sc_hd__a221oi_1 _26447_ (.A1(net2533),
    .A2(\inst$top.soc.cpu.gprf.mem[12][24] ),
    .B1(net1973),
    .B2(\inst$top.soc.cpu.gprf.mem[13][24] ),
    .C1(net2458),
    .Y(_07137_));
 sky130_fd_sc_hd__o21ai_0 _26448_ (.A1(_07135_),
    .A2(_07136_),
    .B1(_07137_),
    .Y(_07138_));
 sky130_fd_sc_hd__nand3_1 _26449_ (.A(_07134_),
    .B(_07138_),
    .C(net2604),
    .Y(_07139_));
 sky130_fd_sc_hd__nor2_1 _26450_ (.A(\inst$top.soc.cpu.gprf.mem[7][24] ),
    .B(net2492),
    .Y(_07140_));
 sky130_fd_sc_hd__o21ai_0 _26451_ (.A1(net2681),
    .A2(\inst$top.soc.cpu.gprf.mem[6][24] ),
    .B1(net2643),
    .Y(_07141_));
 sky130_fd_sc_hd__a22oi_1 _26452_ (.A1(net2532),
    .A2(\inst$top.soc.cpu.gprf.mem[4][24] ),
    .B1(net1972),
    .B2(\inst$top.soc.cpu.gprf.mem[5][24] ),
    .Y(_07142_));
 sky130_fd_sc_hd__o21ai_0 _26453_ (.A1(_07140_),
    .A2(_07141_),
    .B1(_07142_),
    .Y(_07143_));
 sky130_fd_sc_hd__nand2_1 _26454_ (.A(_07143_),
    .B(net1939),
    .Y(_07144_));
 sky130_fd_sc_hd__nor2_1 _26455_ (.A(\inst$top.soc.cpu.gprf.mem[3][24] ),
    .B(net2492),
    .Y(_07145_));
 sky130_fd_sc_hd__o21ai_0 _26456_ (.A1(net2680),
    .A2(\inst$top.soc.cpu.gprf.mem[2][24] ),
    .B1(net2648),
    .Y(_07146_));
 sky130_fd_sc_hd__a22oi_1 _26457_ (.A1(net2535),
    .A2(\inst$top.soc.cpu.gprf.mem[0][24] ),
    .B1(net1975),
    .B2(\inst$top.soc.cpu.gprf.mem[1][24] ),
    .Y(_07147_));
 sky130_fd_sc_hd__o21ai_0 _26458_ (.A1(_07145_),
    .A2(_07146_),
    .B1(_07147_),
    .Y(_07148_));
 sky130_fd_sc_hd__a21oi_1 _26459_ (.A1(_07148_),
    .A2(net2502),
    .B1(net2593),
    .Y(_07149_));
 sky130_fd_sc_hd__nor2_1 _26460_ (.A(\inst$top.soc.cpu.gprf.mem[19][24] ),
    .B(net2493),
    .Y(_07150_));
 sky130_fd_sc_hd__o21ai_0 _26461_ (.A1(net2683),
    .A2(\inst$top.soc.cpu.gprf.mem[18][24] ),
    .B1(net2649),
    .Y(_07151_));
 sky130_fd_sc_hd__a22oi_1 _26462_ (.A1(net2533),
    .A2(\inst$top.soc.cpu.gprf.mem[16][24] ),
    .B1(net1973),
    .B2(\inst$top.soc.cpu.gprf.mem[17][24] ),
    .Y(_07152_));
 sky130_fd_sc_hd__o21ai_0 _26463_ (.A1(_07150_),
    .A2(_07151_),
    .B1(_07152_),
    .Y(_07153_));
 sky130_fd_sc_hd__nor2_1 _26464_ (.A(\inst$top.soc.cpu.gprf.mem[23][24] ),
    .B(net2493),
    .Y(_07154_));
 sky130_fd_sc_hd__o21ai_0 _26465_ (.A1(net2683),
    .A2(\inst$top.soc.cpu.gprf.mem[22][24] ),
    .B1(net2648),
    .Y(_07155_));
 sky130_fd_sc_hd__a22oi_1 _26466_ (.A1(net2533),
    .A2(\inst$top.soc.cpu.gprf.mem[20][24] ),
    .B1(net1973),
    .B2(\inst$top.soc.cpu.gprf.mem[21][24] ),
    .Y(_07156_));
 sky130_fd_sc_hd__o21ai_0 _26467_ (.A1(_07154_),
    .A2(_07155_),
    .B1(_07156_),
    .Y(_07157_));
 sky130_fd_sc_hd__a221oi_1 _26468_ (.A1(_07153_),
    .A2(net2501),
    .B1(net1938),
    .B2(_07157_),
    .C1(net2448),
    .Y(_07158_));
 sky130_fd_sc_hd__nor2_1 _26469_ (.A(\inst$top.soc.cpu.gprf.mem[31][24] ),
    .B(net2488),
    .Y(_07159_));
 sky130_fd_sc_hd__o21ai_0 _26470_ (.A1(net2681),
    .A2(\inst$top.soc.cpu.gprf.mem[30][24] ),
    .B1(net2644),
    .Y(_07160_));
 sky130_fd_sc_hd__a221oi_1 _26471_ (.A1(net2532),
    .A2(\inst$top.soc.cpu.gprf.mem[28][24] ),
    .B1(net1975),
    .B2(\inst$top.soc.cpu.gprf.mem[29][24] ),
    .C1(net2456),
    .Y(_07161_));
 sky130_fd_sc_hd__o21ai_0 _26472_ (.A1(_07159_),
    .A2(_07160_),
    .B1(_07161_),
    .Y(_07162_));
 sky130_fd_sc_hd__nor2_1 _26473_ (.A(\inst$top.soc.cpu.gprf.mem[27][24] ),
    .B(net2492),
    .Y(_07163_));
 sky130_fd_sc_hd__o21ai_0 _26474_ (.A1(net2680),
    .A2(\inst$top.soc.cpu.gprf.mem[26][24] ),
    .B1(net2648),
    .Y(_07164_));
 sky130_fd_sc_hd__a221oi_1 _26475_ (.A1(net2532),
    .A2(\inst$top.soc.cpu.gprf.mem[24][24] ),
    .B1(net1972),
    .B2(\inst$top.soc.cpu.gprf.mem[25][24] ),
    .C1(net2614),
    .Y(_07165_));
 sky130_fd_sc_hd__o21ai_0 _26476_ (.A1(_07163_),
    .A2(_07164_),
    .B1(_07165_),
    .Y(_07166_));
 sky130_fd_sc_hd__nand3_1 _26477_ (.A(_07162_),
    .B(_07166_),
    .C(net2605),
    .Y(_07167_));
 sky130_fd_sc_hd__a32oi_1 _26478_ (.A1(_07139_),
    .A2(_07144_),
    .A3(_07149_),
    .B1(_07158_),
    .B2(_07167_),
    .Y(_00016_));
 sky130_fd_sc_hd__nor2_1 _26479_ (.A(\inst$top.soc.cpu.gprf.mem[31][25] ),
    .B(net2471),
    .Y(_07168_));
 sky130_fd_sc_hd__o21ai_0 _26480_ (.A1(net2660),
    .A2(\inst$top.soc.cpu.gprf.mem[30][25] ),
    .B1(net2625),
    .Y(_07169_));
 sky130_fd_sc_hd__a221oi_1 _26481_ (.A1(net2513),
    .A2(\inst$top.soc.cpu.gprf.mem[28][25] ),
    .B1(net1952),
    .B2(\inst$top.soc.cpu.gprf.mem[29][25] ),
    .C1(net2453),
    .Y(_07170_));
 sky130_fd_sc_hd__o21ai_0 _26482_ (.A1(_07168_),
    .A2(_07169_),
    .B1(_07170_),
    .Y(_07171_));
 sky130_fd_sc_hd__nor2_1 _26483_ (.A(\inst$top.soc.cpu.gprf.mem[27][25] ),
    .B(net2471),
    .Y(_07172_));
 sky130_fd_sc_hd__o21ai_0 _26484_ (.A1(net2660),
    .A2(\inst$top.soc.cpu.gprf.mem[26][25] ),
    .B1(net2625),
    .Y(_07173_));
 sky130_fd_sc_hd__a221oi_1 _26485_ (.A1(net2513),
    .A2(\inst$top.soc.cpu.gprf.mem[24][25] ),
    .B1(net1952),
    .B2(\inst$top.soc.cpu.gprf.mem[25][25] ),
    .C1(net2610),
    .Y(_07174_));
 sky130_fd_sc_hd__o21ai_0 _26486_ (.A1(_07172_),
    .A2(_07173_),
    .B1(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__nand3_1 _26487_ (.A(_07171_),
    .B(_07175_),
    .C(net2598),
    .Y(_07176_));
 sky130_fd_sc_hd__nor2_1 _26488_ (.A(\inst$top.soc.cpu.gprf.mem[19][25] ),
    .B(net2471),
    .Y(_07177_));
 sky130_fd_sc_hd__o21ai_0 _26489_ (.A1(net2660),
    .A2(\inst$top.soc.cpu.gprf.mem[18][25] ),
    .B1(net2625),
    .Y(_07178_));
 sky130_fd_sc_hd__a22oi_1 _26490_ (.A1(net2519),
    .A2(\inst$top.soc.cpu.gprf.mem[16][25] ),
    .B1(net1959),
    .B2(\inst$top.soc.cpu.gprf.mem[17][25] ),
    .Y(_07179_));
 sky130_fd_sc_hd__o21ai_0 _26491_ (.A1(_07177_),
    .A2(_07178_),
    .B1(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__a21oi_1 _26492_ (.A1(_07180_),
    .A2(net2497),
    .B1(net2446),
    .Y(_07181_));
 sky130_fd_sc_hd__nor2_1 _26493_ (.A(\inst$top.soc.cpu.gprf.mem[23][25] ),
    .B(net2471),
    .Y(_07182_));
 sky130_fd_sc_hd__o21ai_0 _26494_ (.A1(net2667),
    .A2(\inst$top.soc.cpu.gprf.mem[22][25] ),
    .B1(net2625),
    .Y(_07183_));
 sky130_fd_sc_hd__a22oi_1 _26495_ (.A1(net2519),
    .A2(\inst$top.soc.cpu.gprf.mem[20][25] ),
    .B1(net1959),
    .B2(\inst$top.soc.cpu.gprf.mem[21][25] ),
    .Y(_07184_));
 sky130_fd_sc_hd__o21ai_0 _26496_ (.A1(_07182_),
    .A2(_07183_),
    .B1(_07184_),
    .Y(_07185_));
 sky130_fd_sc_hd__nand2_1 _26497_ (.A(_07185_),
    .B(net1935),
    .Y(_07186_));
 sky130_fd_sc_hd__nor2_1 _26498_ (.A(\inst$top.soc.cpu.gprf.mem[3][25] ),
    .B(net2471),
    .Y(_07187_));
 sky130_fd_sc_hd__o21ai_0 _26499_ (.A1(net2660),
    .A2(\inst$top.soc.cpu.gprf.mem[2][25] ),
    .B1(net2625),
    .Y(_07188_));
 sky130_fd_sc_hd__a22oi_1 _26500_ (.A1(net2513),
    .A2(\inst$top.soc.cpu.gprf.mem[0][25] ),
    .B1(net1952),
    .B2(\inst$top.soc.cpu.gprf.mem[1][25] ),
    .Y(_07189_));
 sky130_fd_sc_hd__o21ai_0 _26501_ (.A1(_07187_),
    .A2(_07188_),
    .B1(_07189_),
    .Y(_07190_));
 sky130_fd_sc_hd__nor2_1 _26502_ (.A(\inst$top.soc.cpu.gprf.mem[7][25] ),
    .B(net2471),
    .Y(_07191_));
 sky130_fd_sc_hd__o21ai_0 _26503_ (.A1(net2667),
    .A2(\inst$top.soc.cpu.gprf.mem[6][25] ),
    .B1(net2625),
    .Y(_07192_));
 sky130_fd_sc_hd__a22oi_1 _26504_ (.A1(net2526),
    .A2(\inst$top.soc.cpu.gprf.mem[4][25] ),
    .B1(net1959),
    .B2(\inst$top.soc.cpu.gprf.mem[5][25] ),
    .Y(_07193_));
 sky130_fd_sc_hd__o21ai_0 _26505_ (.A1(_07191_),
    .A2(_07192_),
    .B1(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__a221oi_1 _26506_ (.A1(_07190_),
    .A2(net2497),
    .B1(net1935),
    .B2(_07194_),
    .C1(net2592),
    .Y(_07195_));
 sky130_fd_sc_hd__nor2_1 _26507_ (.A(\inst$top.soc.cpu.gprf.mem[15][25] ),
    .B(net2471),
    .Y(_07196_));
 sky130_fd_sc_hd__o21ai_0 _26508_ (.A1(net2667),
    .A2(\inst$top.soc.cpu.gprf.mem[14][25] ),
    .B1(net2626),
    .Y(_07197_));
 sky130_fd_sc_hd__a221oi_1 _26509_ (.A1(net2519),
    .A2(\inst$top.soc.cpu.gprf.mem[12][25] ),
    .B1(net1966),
    .B2(\inst$top.soc.cpu.gprf.mem[13][25] ),
    .C1(net2454),
    .Y(_07198_));
 sky130_fd_sc_hd__o21ai_0 _26510_ (.A1(_07196_),
    .A2(_07197_),
    .B1(_07198_),
    .Y(_07199_));
 sky130_fd_sc_hd__nor2_1 _26511_ (.A(\inst$top.soc.cpu.gprf.mem[11][25] ),
    .B(net2471),
    .Y(_07200_));
 sky130_fd_sc_hd__o21ai_0 _26512_ (.A1(net2667),
    .A2(\inst$top.soc.cpu.gprf.mem[10][25] ),
    .B1(net2625),
    .Y(_07201_));
 sky130_fd_sc_hd__a221oi_1 _26513_ (.A1(net2519),
    .A2(\inst$top.soc.cpu.gprf.mem[8][25] ),
    .B1(net1959),
    .B2(\inst$top.soc.cpu.gprf.mem[9][25] ),
    .C1(net2610),
    .Y(_07202_));
 sky130_fd_sc_hd__o21ai_0 _26514_ (.A1(_07200_),
    .A2(_07201_),
    .B1(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__nand3_1 _26515_ (.A(_07199_),
    .B(_07203_),
    .C(net2601),
    .Y(_07204_));
 sky130_fd_sc_hd__a32oi_2 _26516_ (.A1(_07176_),
    .A2(_07181_),
    .A3(_07186_),
    .B1(_07195_),
    .B2(_07204_),
    .Y(_00017_));
 sky130_fd_sc_hd__nor2_1 _26517_ (.A(\inst$top.soc.cpu.gprf.mem[11][26] ),
    .B(net2462),
    .Y(_07205_));
 sky130_fd_sc_hd__o21ai_0 _26518_ (.A1(net2653),
    .A2(\inst$top.soc.cpu.gprf.mem[10][26] ),
    .B1(net2617),
    .Y(_07206_));
 sky130_fd_sc_hd__a221oi_1 _26519_ (.A1(net2506),
    .A2(\inst$top.soc.cpu.gprf.mem[8][26] ),
    .B1(net1945),
    .B2(\inst$top.soc.cpu.gprf.mem[9][26] ),
    .C1(net2607),
    .Y(_07207_));
 sky130_fd_sc_hd__o21ai_0 _26520_ (.A1(_07205_),
    .A2(_07206_),
    .B1(_07207_),
    .Y(_07208_));
 sky130_fd_sc_hd__nor2_1 _26521_ (.A(\inst$top.soc.cpu.gprf.mem[15][26] ),
    .B(net2466),
    .Y(_07209_));
 sky130_fd_sc_hd__o21ai_0 _26522_ (.A1(net2653),
    .A2(\inst$top.soc.cpu.gprf.mem[14][26] ),
    .B1(net2621),
    .Y(_07210_));
 sky130_fd_sc_hd__a221oi_1 _26523_ (.A1(net2510),
    .A2(\inst$top.soc.cpu.gprf.mem[12][26] ),
    .B1(net1949),
    .B2(\inst$top.soc.cpu.gprf.mem[13][26] ),
    .C1(net2451),
    .Y(_07211_));
 sky130_fd_sc_hd__o21ai_0 _26524_ (.A1(_07209_),
    .A2(_07210_),
    .B1(_07211_),
    .Y(_07212_));
 sky130_fd_sc_hd__nand3_1 _26525_ (.A(_07208_),
    .B(_07212_),
    .C(net2600),
    .Y(_07213_));
 sky130_fd_sc_hd__nor2_1 _26526_ (.A(\inst$top.soc.cpu.gprf.mem[7][26] ),
    .B(net2468),
    .Y(_07214_));
 sky130_fd_sc_hd__o21ai_0 _26527_ (.A1(net2654),
    .A2(\inst$top.soc.cpu.gprf.mem[6][26] ),
    .B1(net2622),
    .Y(_07215_));
 sky130_fd_sc_hd__a22oi_1 _26528_ (.A1(net2507),
    .A2(\inst$top.soc.cpu.gprf.mem[4][26] ),
    .B1(net1950),
    .B2(\inst$top.soc.cpu.gprf.mem[5][26] ),
    .Y(_07216_));
 sky130_fd_sc_hd__o21ai_0 _26529_ (.A1(_07214_),
    .A2(_07215_),
    .B1(_07216_),
    .Y(_07217_));
 sky130_fd_sc_hd__nand2_1 _26530_ (.A(_07217_),
    .B(net1934),
    .Y(_07218_));
 sky130_fd_sc_hd__nor2_1 _26531_ (.A(\inst$top.soc.cpu.gprf.mem[3][26] ),
    .B(net2462),
    .Y(_07219_));
 sky130_fd_sc_hd__o21ai_0 _26532_ (.A1(net2654),
    .A2(\inst$top.soc.cpu.gprf.mem[2][26] ),
    .B1(net2617),
    .Y(_07220_));
 sky130_fd_sc_hd__a22oi_1 _26533_ (.A1(net2507),
    .A2(\inst$top.soc.cpu.gprf.mem[0][26] ),
    .B1(net1946),
    .B2(\inst$top.soc.cpu.gprf.mem[1][26] ),
    .Y(_07221_));
 sky130_fd_sc_hd__o21ai_0 _26534_ (.A1(_07219_),
    .A2(_07220_),
    .B1(_07221_),
    .Y(_07222_));
 sky130_fd_sc_hd__a21oi_1 _26535_ (.A1(_07222_),
    .A2(net2496),
    .B1(net2592),
    .Y(_07223_));
 sky130_fd_sc_hd__nor2_1 _26536_ (.A(\inst$top.soc.cpu.gprf.mem[19][26] ),
    .B(net2468),
    .Y(_07224_));
 sky130_fd_sc_hd__o21ai_0 _26537_ (.A1(net2658),
    .A2(\inst$top.soc.cpu.gprf.mem[18][26] ),
    .B1(net2622),
    .Y(_07225_));
 sky130_fd_sc_hd__a22oi_1 _26538_ (.A1(net2511),
    .A2(\inst$top.soc.cpu.gprf.mem[16][26] ),
    .B1(net1950),
    .B2(\inst$top.soc.cpu.gprf.mem[17][26] ),
    .Y(_07226_));
 sky130_fd_sc_hd__o21ai_0 _26539_ (.A1(_07224_),
    .A2(_07225_),
    .B1(_07226_),
    .Y(_07227_));
 sky130_fd_sc_hd__nor2_1 _26540_ (.A(\inst$top.soc.cpu.gprf.mem[23][26] ),
    .B(net2468),
    .Y(_07228_));
 sky130_fd_sc_hd__o21ai_0 _26541_ (.A1(net2658),
    .A2(\inst$top.soc.cpu.gprf.mem[22][26] ),
    .B1(net2622),
    .Y(_07229_));
 sky130_fd_sc_hd__a22oi_1 _26542_ (.A1(net2510),
    .A2(\inst$top.soc.cpu.gprf.mem[20][26] ),
    .B1(net1949),
    .B2(\inst$top.soc.cpu.gprf.mem[21][26] ),
    .Y(_07230_));
 sky130_fd_sc_hd__o21ai_0 _26543_ (.A1(_07228_),
    .A2(_07229_),
    .B1(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__a221oi_1 _26544_ (.A1(net2511),
    .A2(\inst$top.soc.cpu.gprf.mem[28][26] ),
    .B1(net1950),
    .B2(\inst$top.soc.cpu.gprf.mem[29][26] ),
    .C1(net2451),
    .Y(_07232_));
 sky130_fd_sc_hd__nor2_1 _26545_ (.A(net2658),
    .B(\inst$top.soc.cpu.gprf.mem[30][26] ),
    .Y(_07233_));
 sky130_fd_sc_hd__nor2_1 _26546_ (.A(_20261_),
    .B(_07233_),
    .Y(_07234_));
 sky130_fd_sc_hd__o21ai_0 _26547_ (.A1(net2468),
    .A2(\inst$top.soc.cpu.gprf.mem[31][26] ),
    .B1(_07234_),
    .Y(_07235_));
 sky130_fd_sc_hd__nor2_1 _26548_ (.A(\inst$top.soc.cpu.gprf.mem[27][26] ),
    .B(net2468),
    .Y(_07236_));
 sky130_fd_sc_hd__o21ai_0 _26549_ (.A1(net2658),
    .A2(\inst$top.soc.cpu.gprf.mem[26][26] ),
    .B1(net2622),
    .Y(_07237_));
 sky130_fd_sc_hd__nor2_1 _26550_ (.A(_07236_),
    .B(_07237_),
    .Y(_07238_));
 sky130_fd_sc_hd__inv_1 _26551_ (.A(\inst$top.soc.cpu.gprf.mem[24][26] ),
    .Y(_07239_));
 sky130_fd_sc_hd__o21ai_0 _26552_ (.A1(_07239_),
    .A2(_20236_),
    .B1(net2451),
    .Y(_07240_));
 sky130_fd_sc_hd__a211oi_1 _26553_ (.A1(\inst$top.soc.cpu.gprf.mem[25][26] ),
    .A2(net1950),
    .B1(_07238_),
    .C1(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__a211oi_1 _26554_ (.A1(_07232_),
    .A2(_07235_),
    .B1(_06038_),
    .C1(_07241_),
    .Y(_07242_));
 sky130_fd_sc_hd__a221oi_1 _26555_ (.A1(net2499),
    .A2(_07227_),
    .B1(net1934),
    .B2(_07231_),
    .C1(_07242_),
    .Y(_07243_));
 sky130_fd_sc_hd__a32oi_1 _26556_ (.A1(_07213_),
    .A2(_07218_),
    .A3(_07223_),
    .B1(_07243_),
    .B2(net2592),
    .Y(_00018_));
 sky130_fd_sc_hd__nor2_1 _26557_ (.A(\inst$top.soc.cpu.gprf.mem[15][27] ),
    .B(net2479),
    .Y(_07244_));
 sky130_fd_sc_hd__o21ai_0 _26558_ (.A1(net2668),
    .A2(\inst$top.soc.cpu.gprf.mem[14][27] ),
    .B1(net2634),
    .Y(_07245_));
 sky130_fd_sc_hd__a221oi_1 _26559_ (.A1(net2520),
    .A2(\inst$top.soc.cpu.gprf.mem[12][27] ),
    .B1(net1960),
    .B2(\inst$top.soc.cpu.gprf.mem[13][27] ),
    .C1(net2456),
    .Y(_07246_));
 sky130_fd_sc_hd__o21ai_0 _26560_ (.A1(_07244_),
    .A2(_07245_),
    .B1(_07246_),
    .Y(_07247_));
 sky130_fd_sc_hd__nor2_1 _26561_ (.A(\inst$top.soc.cpu.gprf.mem[11][27] ),
    .B(net2480),
    .Y(_07248_));
 sky130_fd_sc_hd__o21ai_0 _26562_ (.A1(net2675),
    .A2(\inst$top.soc.cpu.gprf.mem[10][27] ),
    .B1(net2634),
    .Y(_07249_));
 sky130_fd_sc_hd__a221oi_1 _26563_ (.A1(net2527),
    .A2(\inst$top.soc.cpu.gprf.mem[8][27] ),
    .B1(net1967),
    .B2(\inst$top.soc.cpu.gprf.mem[9][27] ),
    .C1(net2611),
    .Y(_07250_));
 sky130_fd_sc_hd__o21ai_0 _26564_ (.A1(_07248_),
    .A2(_07249_),
    .B1(_07250_),
    .Y(_07251_));
 sky130_fd_sc_hd__nand3_1 _26565_ (.A(_07247_),
    .B(_07251_),
    .C(net2601),
    .Y(_07252_));
 sky130_fd_sc_hd__nor2_1 _26566_ (.A(\inst$top.soc.cpu.gprf.mem[7][27] ),
    .B(net2479),
    .Y(_07253_));
 sky130_fd_sc_hd__o21ai_0 _26567_ (.A1(net2668),
    .A2(\inst$top.soc.cpu.gprf.mem[6][27] ),
    .B1(net2633),
    .Y(_07254_));
 sky130_fd_sc_hd__a22oi_1 _26568_ (.A1(net2520),
    .A2(\inst$top.soc.cpu.gprf.mem[4][27] ),
    .B1(net1960),
    .B2(\inst$top.soc.cpu.gprf.mem[5][27] ),
    .Y(_07255_));
 sky130_fd_sc_hd__o21ai_0 _26569_ (.A1(_07253_),
    .A2(_07254_),
    .B1(_07255_),
    .Y(_07256_));
 sky130_fd_sc_hd__nand2_1 _26570_ (.A(_07256_),
    .B(net1937),
    .Y(_07257_));
 sky130_fd_sc_hd__nor2_1 _26571_ (.A(\inst$top.soc.cpu.gprf.mem[3][27] ),
    .B(net2479),
    .Y(_07258_));
 sky130_fd_sc_hd__o21ai_0 _26572_ (.A1(net2668),
    .A2(\inst$top.soc.cpu.gprf.mem[2][27] ),
    .B1(net2634),
    .Y(_07259_));
 sky130_fd_sc_hd__a22oi_1 _26573_ (.A1(net2520),
    .A2(\inst$top.soc.cpu.gprf.mem[0][27] ),
    .B1(net1960),
    .B2(\inst$top.soc.cpu.gprf.mem[1][27] ),
    .Y(_07260_));
 sky130_fd_sc_hd__o21ai_0 _26574_ (.A1(_07258_),
    .A2(_07259_),
    .B1(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__a21oi_1 _26575_ (.A1(_07261_),
    .A2(net2500),
    .B1(net2593),
    .Y(_07262_));
 sky130_fd_sc_hd__nor2_1 _26576_ (.A(\inst$top.soc.cpu.gprf.mem[23][27] ),
    .B(net2479),
    .Y(_07263_));
 sky130_fd_sc_hd__o21ai_0 _26577_ (.A1(net2668),
    .A2(\inst$top.soc.cpu.gprf.mem[22][27] ),
    .B1(net2633),
    .Y(_07264_));
 sky130_fd_sc_hd__a22oi_1 _26578_ (.A1(net2520),
    .A2(\inst$top.soc.cpu.gprf.mem[20][27] ),
    .B1(net1960),
    .B2(\inst$top.soc.cpu.gprf.mem[21][27] ),
    .Y(_07265_));
 sky130_fd_sc_hd__o21ai_0 _26579_ (.A1(_07263_),
    .A2(_07264_),
    .B1(_07265_),
    .Y(_07266_));
 sky130_fd_sc_hd__nor2_1 _26580_ (.A(\inst$top.soc.cpu.gprf.mem[19][27] ),
    .B(net2479),
    .Y(_07267_));
 sky130_fd_sc_hd__o21ai_0 _26581_ (.A1(net2668),
    .A2(\inst$top.soc.cpu.gprf.mem[18][27] ),
    .B1(net2633),
    .Y(_07268_));
 sky130_fd_sc_hd__a22oi_1 _26582_ (.A1(net2520),
    .A2(\inst$top.soc.cpu.gprf.mem[16][27] ),
    .B1(net1960),
    .B2(\inst$top.soc.cpu.gprf.mem[17][27] ),
    .Y(_07269_));
 sky130_fd_sc_hd__o21ai_0 _26583_ (.A1(_07267_),
    .A2(_07268_),
    .B1(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__a221oi_1 _26584_ (.A1(_07266_),
    .A2(net1937),
    .B1(net2500),
    .B2(_07270_),
    .C1(net2447),
    .Y(_07271_));
 sky130_fd_sc_hd__nor2_1 _26585_ (.A(\inst$top.soc.cpu.gprf.mem[31][27] ),
    .B(net2480),
    .Y(_07272_));
 sky130_fd_sc_hd__o21ai_0 _26586_ (.A1(net2675),
    .A2(\inst$top.soc.cpu.gprf.mem[30][27] ),
    .B1(net2634),
    .Y(_07273_));
 sky130_fd_sc_hd__a221oi_1 _26587_ (.A1(net2520),
    .A2(\inst$top.soc.cpu.gprf.mem[28][27] ),
    .B1(net1960),
    .B2(\inst$top.soc.cpu.gprf.mem[29][27] ),
    .C1(net2456),
    .Y(_07274_));
 sky130_fd_sc_hd__o21ai_0 _26588_ (.A1(_07272_),
    .A2(_07273_),
    .B1(_07274_),
    .Y(_07275_));
 sky130_fd_sc_hd__nor2_1 _26589_ (.A(\inst$top.soc.cpu.gprf.mem[27][27] ),
    .B(net2479),
    .Y(_07276_));
 sky130_fd_sc_hd__o21ai_0 _26590_ (.A1(net2668),
    .A2(\inst$top.soc.cpu.gprf.mem[26][27] ),
    .B1(net2633),
    .Y(_07277_));
 sky130_fd_sc_hd__a221oi_1 _26591_ (.A1(net2527),
    .A2(\inst$top.soc.cpu.gprf.mem[24][27] ),
    .B1(net1967),
    .B2(\inst$top.soc.cpu.gprf.mem[25][27] ),
    .C1(net2611),
    .Y(_07278_));
 sky130_fd_sc_hd__o21ai_0 _26592_ (.A1(_07276_),
    .A2(_07277_),
    .B1(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__nand3_1 _26593_ (.A(_07275_),
    .B(_07279_),
    .C(net2601),
    .Y(_07280_));
 sky130_fd_sc_hd__a32oi_1 _26594_ (.A1(_07252_),
    .A2(_07257_),
    .A3(_07262_),
    .B1(_07271_),
    .B2(_07280_),
    .Y(_00019_));
 sky130_fd_sc_hd__nor2_1 _26595_ (.A(\inst$top.soc.cpu.gprf.mem[11][28] ),
    .B(net2481),
    .Y(_07281_));
 sky130_fd_sc_hd__o21ai_0 _26596_ (.A1(net2676),
    .A2(\inst$top.soc.cpu.gprf.mem[10][28] ),
    .B1(net2636),
    .Y(_07282_));
 sky130_fd_sc_hd__a221oi_1 _26597_ (.A1(net2528),
    .A2(\inst$top.soc.cpu.gprf.mem[8][28] ),
    .B1(net1968),
    .B2(\inst$top.soc.cpu.gprf.mem[9][28] ),
    .C1(net2611),
    .Y(_07283_));
 sky130_fd_sc_hd__o21ai_0 _26598_ (.A1(_07281_),
    .A2(_07282_),
    .B1(_07283_),
    .Y(_07284_));
 sky130_fd_sc_hd__nor2_1 _26599_ (.A(\inst$top.soc.cpu.gprf.mem[15][28] ),
    .B(net2482),
    .Y(_07285_));
 sky130_fd_sc_hd__o21ai_0 _26600_ (.A1(net2668),
    .A2(\inst$top.soc.cpu.gprf.mem[14][28] ),
    .B1(net2635),
    .Y(_07286_));
 sky130_fd_sc_hd__a221oi_1 _26601_ (.A1(net2520),
    .A2(\inst$top.soc.cpu.gprf.mem[12][28] ),
    .B1(net1961),
    .B2(\inst$top.soc.cpu.gprf.mem[13][28] ),
    .C1(net2456),
    .Y(_07287_));
 sky130_fd_sc_hd__o21ai_0 _26602_ (.A1(_07285_),
    .A2(_07286_),
    .B1(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__nand3_1 _26603_ (.A(_07284_),
    .B(_07288_),
    .C(net2603),
    .Y(_07289_));
 sky130_fd_sc_hd__nor2_1 _26604_ (.A(\inst$top.soc.cpu.gprf.mem[7][28] ),
    .B(net2481),
    .Y(_07290_));
 sky130_fd_sc_hd__o21ai_0 _26605_ (.A1(net2669),
    .A2(\inst$top.soc.cpu.gprf.mem[6][28] ),
    .B1(net2635),
    .Y(_07291_));
 sky130_fd_sc_hd__a22oi_1 _26606_ (.A1(net2521),
    .A2(\inst$top.soc.cpu.gprf.mem[4][28] ),
    .B1(net1961),
    .B2(\inst$top.soc.cpu.gprf.mem[5][28] ),
    .Y(_07292_));
 sky130_fd_sc_hd__o21ai_0 _26607_ (.A1(_07290_),
    .A2(_07291_),
    .B1(_07292_),
    .Y(_07293_));
 sky130_fd_sc_hd__nand2_1 _26608_ (.A(_07293_),
    .B(net1937),
    .Y(_07294_));
 sky130_fd_sc_hd__nor2_1 _26609_ (.A(\inst$top.soc.cpu.gprf.mem[3][28] ),
    .B(net2481),
    .Y(_07295_));
 sky130_fd_sc_hd__o21ai_0 _26610_ (.A1(net2669),
    .A2(\inst$top.soc.cpu.gprf.mem[2][28] ),
    .B1(net2636),
    .Y(_07296_));
 sky130_fd_sc_hd__a22oi_1 _26611_ (.A1(net2521),
    .A2(\inst$top.soc.cpu.gprf.mem[0][28] ),
    .B1(net1961),
    .B2(\inst$top.soc.cpu.gprf.mem[1][28] ),
    .Y(_07297_));
 sky130_fd_sc_hd__o21ai_0 _26612_ (.A1(_07295_),
    .A2(_07296_),
    .B1(_07297_),
    .Y(_07298_));
 sky130_fd_sc_hd__a21oi_1 _26613_ (.A1(_07298_),
    .A2(net2500),
    .B1(net2593),
    .Y(_07299_));
 sky130_fd_sc_hd__nor2_1 _26614_ (.A(\inst$top.soc.cpu.gprf.mem[19][28] ),
    .B(net2484),
    .Y(_07300_));
 sky130_fd_sc_hd__o21ai_0 _26615_ (.A1(net2676),
    .A2(\inst$top.soc.cpu.gprf.mem[18][28] ),
    .B1(net2639),
    .Y(_07301_));
 sky130_fd_sc_hd__a22oi_1 _26616_ (.A1(net2528),
    .A2(\inst$top.soc.cpu.gprf.mem[16][28] ),
    .B1(net1968),
    .B2(\inst$top.soc.cpu.gprf.mem[17][28] ),
    .Y(_07302_));
 sky130_fd_sc_hd__o21ai_0 _26617_ (.A1(_07300_),
    .A2(_07301_),
    .B1(_07302_),
    .Y(_07303_));
 sky130_fd_sc_hd__nor2_1 _26618_ (.A(\inst$top.soc.cpu.gprf.mem[23][28] ),
    .B(net2481),
    .Y(_07304_));
 sky130_fd_sc_hd__o21ai_0 _26619_ (.A1(net2676),
    .A2(\inst$top.soc.cpu.gprf.mem[22][28] ),
    .B1(net2639),
    .Y(_07305_));
 sky130_fd_sc_hd__a22oi_1 _26620_ (.A1(net2528),
    .A2(\inst$top.soc.cpu.gprf.mem[20][28] ),
    .B1(net1968),
    .B2(\inst$top.soc.cpu.gprf.mem[21][28] ),
    .Y(_07306_));
 sky130_fd_sc_hd__o21ai_0 _26621_ (.A1(_07304_),
    .A2(_07305_),
    .B1(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__a221oi_1 _26622_ (.A1(_07303_),
    .A2(net2501),
    .B1(net1938),
    .B2(_07307_),
    .C1(net2448),
    .Y(_07308_));
 sky130_fd_sc_hd__nor2_1 _26623_ (.A(\inst$top.soc.cpu.gprf.mem[31][28] ),
    .B(net2481),
    .Y(_07309_));
 sky130_fd_sc_hd__o21ai_0 _26624_ (.A1(net2676),
    .A2(\inst$top.soc.cpu.gprf.mem[30][28] ),
    .B1(net2636),
    .Y(_07310_));
 sky130_fd_sc_hd__a221oi_1 _26625_ (.A1(net2528),
    .A2(\inst$top.soc.cpu.gprf.mem[28][28] ),
    .B1(net1968),
    .B2(\inst$top.soc.cpu.gprf.mem[29][28] ),
    .C1(net2456),
    .Y(_07311_));
 sky130_fd_sc_hd__o21ai_0 _26626_ (.A1(_07309_),
    .A2(_07310_),
    .B1(_07311_),
    .Y(_07312_));
 sky130_fd_sc_hd__nor2_1 _26627_ (.A(\inst$top.soc.cpu.gprf.mem[27][28] ),
    .B(net2481),
    .Y(_07313_));
 sky130_fd_sc_hd__o21ai_0 _26628_ (.A1(net2675),
    .A2(\inst$top.soc.cpu.gprf.mem[26][28] ),
    .B1(net2635),
    .Y(_07314_));
 sky130_fd_sc_hd__a221oi_1 _26629_ (.A1(net2528),
    .A2(\inst$top.soc.cpu.gprf.mem[24][28] ),
    .B1(net1968),
    .B2(\inst$top.soc.cpu.gprf.mem[25][28] ),
    .C1(net2611),
    .Y(_07315_));
 sky130_fd_sc_hd__o21ai_0 _26630_ (.A1(_07313_),
    .A2(_07314_),
    .B1(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__nand3_1 _26631_ (.A(_07312_),
    .B(_07316_),
    .C(net2603),
    .Y(_07317_));
 sky130_fd_sc_hd__a32oi_1 _26632_ (.A1(_07289_),
    .A2(_07294_),
    .A3(_07299_),
    .B1(_07308_),
    .B2(_07317_),
    .Y(_00020_));
 sky130_fd_sc_hd__nor2_1 _26633_ (.A(\inst$top.soc.cpu.gprf.mem[15][29] ),
    .B(net2488),
    .Y(_07318_));
 sky130_fd_sc_hd__o21ai_0 _26634_ (.A1(net2673),
    .A2(\inst$top.soc.cpu.gprf.mem[14][29] ),
    .B1(net2643),
    .Y(_07319_));
 sky130_fd_sc_hd__a221oi_1 _26635_ (.A1(net2525),
    .A2(\inst$top.soc.cpu.gprf.mem[12][29] ),
    .B1(net1964),
    .B2(\inst$top.soc.cpu.gprf.mem[13][29] ),
    .C1(net2456),
    .Y(_07320_));
 sky130_fd_sc_hd__o21ai_0 _26636_ (.A1(_07318_),
    .A2(_07319_),
    .B1(_07320_),
    .Y(_07321_));
 sky130_fd_sc_hd__nor2_1 _26637_ (.A(\inst$top.soc.cpu.gprf.mem[11][29] ),
    .B(net2488),
    .Y(_07322_));
 sky130_fd_sc_hd__o21ai_0 _26638_ (.A1(net2672),
    .A2(\inst$top.soc.cpu.gprf.mem[10][29] ),
    .B1(net2643),
    .Y(_07323_));
 sky130_fd_sc_hd__a221oi_1 _26639_ (.A1(net2524),
    .A2(\inst$top.soc.cpu.gprf.mem[8][29] ),
    .B1(net1965),
    .B2(\inst$top.soc.cpu.gprf.mem[9][29] ),
    .C1(net2613),
    .Y(_07324_));
 sky130_fd_sc_hd__o21ai_0 _26640_ (.A1(_07322_),
    .A2(_07323_),
    .B1(_07324_),
    .Y(_07325_));
 sky130_fd_sc_hd__nand3_1 _26641_ (.A(_07321_),
    .B(_07325_),
    .C(net2602),
    .Y(_07326_));
 sky130_fd_sc_hd__nor2_1 _26642_ (.A(\inst$top.soc.cpu.gprf.mem[7][29] ),
    .B(net2488),
    .Y(_07327_));
 sky130_fd_sc_hd__o21ai_0 _26643_ (.A1(net2673),
    .A2(\inst$top.soc.cpu.gprf.mem[6][29] ),
    .B1(net2643),
    .Y(_07328_));
 sky130_fd_sc_hd__a22oi_1 _26644_ (.A1(net2525),
    .A2(\inst$top.soc.cpu.gprf.mem[4][29] ),
    .B1(net1965),
    .B2(\inst$top.soc.cpu.gprf.mem[5][29] ),
    .Y(_07329_));
 sky130_fd_sc_hd__o21ai_0 _26645_ (.A1(_07327_),
    .A2(_07328_),
    .B1(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__nand2_1 _26646_ (.A(_07330_),
    .B(net1937),
    .Y(_07331_));
 sky130_fd_sc_hd__nor2_1 _26647_ (.A(\inst$top.soc.cpu.gprf.mem[3][29] ),
    .B(net2476),
    .Y(_07332_));
 sky130_fd_sc_hd__o21ai_0 _26648_ (.A1(net2670),
    .A2(\inst$top.soc.cpu.gprf.mem[2][29] ),
    .B1(net2629),
    .Y(_07333_));
 sky130_fd_sc_hd__a22oi_1 _26649_ (.A1(net2522),
    .A2(\inst$top.soc.cpu.gprf.mem[0][29] ),
    .B1(net1962),
    .B2(\inst$top.soc.cpu.gprf.mem[1][29] ),
    .Y(_07334_));
 sky130_fd_sc_hd__o21ai_0 _26650_ (.A1(_07332_),
    .A2(_07333_),
    .B1(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__a21oi_1 _26651_ (.A1(_07335_),
    .A2(net2500),
    .B1(net2594),
    .Y(_07336_));
 sky130_fd_sc_hd__nor2_1 _26652_ (.A(\inst$top.soc.cpu.gprf.mem[23][29] ),
    .B(net2476),
    .Y(_07337_));
 sky130_fd_sc_hd__o21ai_0 _26653_ (.A1(net2670),
    .A2(\inst$top.soc.cpu.gprf.mem[22][29] ),
    .B1(net2629),
    .Y(_07338_));
 sky130_fd_sc_hd__a22oi_1 _26654_ (.A1(net2522),
    .A2(\inst$top.soc.cpu.gprf.mem[20][29] ),
    .B1(net1962),
    .B2(\inst$top.soc.cpu.gprf.mem[21][29] ),
    .Y(_07339_));
 sky130_fd_sc_hd__o21ai_0 _26655_ (.A1(_07337_),
    .A2(_07338_),
    .B1(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__nor2_1 _26656_ (.A(\inst$top.soc.cpu.gprf.mem[19][29] ),
    .B(net2488),
    .Y(_07341_));
 sky130_fd_sc_hd__o21ai_0 _26657_ (.A1(net2670),
    .A2(\inst$top.soc.cpu.gprf.mem[18][29] ),
    .B1(net2643),
    .Y(_07342_));
 sky130_fd_sc_hd__a22oi_1 _26658_ (.A1(net2525),
    .A2(\inst$top.soc.cpu.gprf.mem[16][29] ),
    .B1(net1965),
    .B2(\inst$top.soc.cpu.gprf.mem[17][29] ),
    .Y(_07343_));
 sky130_fd_sc_hd__o21ai_0 _26659_ (.A1(_07341_),
    .A2(_07342_),
    .B1(_07343_),
    .Y(_07344_));
 sky130_fd_sc_hd__a221oi_1 _26660_ (.A1(_07340_),
    .A2(net1937),
    .B1(net2503),
    .B2(_07344_),
    .C1(net2447),
    .Y(_07345_));
 sky130_fd_sc_hd__nor2_1 _26661_ (.A(\inst$top.soc.cpu.gprf.mem[31][29] ),
    .B(net2476),
    .Y(_07346_));
 sky130_fd_sc_hd__o21ai_0 _26662_ (.A1(net2671),
    .A2(\inst$top.soc.cpu.gprf.mem[30][29] ),
    .B1(net2630),
    .Y(_07347_));
 sky130_fd_sc_hd__a221oi_1 _26663_ (.A1(net2522),
    .A2(\inst$top.soc.cpu.gprf.mem[28][29] ),
    .B1(net1963),
    .B2(\inst$top.soc.cpu.gprf.mem[29][29] ),
    .C1(net2454),
    .Y(_07348_));
 sky130_fd_sc_hd__o21ai_0 _26664_ (.A1(_07346_),
    .A2(_07347_),
    .B1(_07348_),
    .Y(_07349_));
 sky130_fd_sc_hd__nor2_1 _26665_ (.A(\inst$top.soc.cpu.gprf.mem[27][29] ),
    .B(net2488),
    .Y(_07350_));
 sky130_fd_sc_hd__o21ai_0 _26666_ (.A1(net2670),
    .A2(\inst$top.soc.cpu.gprf.mem[26][29] ),
    .B1(net2643),
    .Y(_07351_));
 sky130_fd_sc_hd__a221oi_1 _26667_ (.A1(net2522),
    .A2(\inst$top.soc.cpu.gprf.mem[24][29] ),
    .B1(net1962),
    .B2(\inst$top.soc.cpu.gprf.mem[25][29] ),
    .C1(net2615),
    .Y(_07352_));
 sky130_fd_sc_hd__o21ai_0 _26668_ (.A1(_07350_),
    .A2(_07351_),
    .B1(_07352_),
    .Y(_07353_));
 sky130_fd_sc_hd__nand3_1 _26669_ (.A(_07349_),
    .B(_07353_),
    .C(net2602),
    .Y(_07354_));
 sky130_fd_sc_hd__a32oi_1 _26670_ (.A1(_07326_),
    .A2(_07331_),
    .A3(_07336_),
    .B1(_07345_),
    .B2(_07354_),
    .Y(_00021_));
 sky130_fd_sc_hd__nor2_1 _26671_ (.A(\inst$top.soc.cpu.gprf.mem[11][30] ),
    .B(net2477),
    .Y(_07355_));
 sky130_fd_sc_hd__o21ai_0 _26672_ (.A1(net2662),
    .A2(\inst$top.soc.cpu.gprf.mem[10][30] ),
    .B1(net2631),
    .Y(_07356_));
 sky130_fd_sc_hd__a221oi_1 _26673_ (.A1(net2513),
    .A2(\inst$top.soc.cpu.gprf.mem[8][30] ),
    .B1(net1951),
    .B2(\inst$top.soc.cpu.gprf.mem[9][30] ),
    .C1(net2609),
    .Y(_07357_));
 sky130_fd_sc_hd__o21ai_0 _26674_ (.A1(_07355_),
    .A2(_07356_),
    .B1(_07357_),
    .Y(_07358_));
 sky130_fd_sc_hd__nor2_1 _26675_ (.A(\inst$top.soc.cpu.gprf.mem[15][30] ),
    .B(net2471),
    .Y(_07359_));
 sky130_fd_sc_hd__o21ai_0 _26676_ (.A1(net2659),
    .A2(\inst$top.soc.cpu.gprf.mem[14][30] ),
    .B1(net2625),
    .Y(_07360_));
 sky130_fd_sc_hd__a221oi_1 _26677_ (.A1(net2513),
    .A2(\inst$top.soc.cpu.gprf.mem[12][30] ),
    .B1(net1952),
    .B2(\inst$top.soc.cpu.gprf.mem[13][30] ),
    .C1(net2455),
    .Y(_07361_));
 sky130_fd_sc_hd__o21ai_0 _26678_ (.A1(_07359_),
    .A2(_07360_),
    .B1(_07361_),
    .Y(_07362_));
 sky130_fd_sc_hd__nand3_1 _26679_ (.A(_07358_),
    .B(_07362_),
    .C(net2598),
    .Y(_07363_));
 sky130_fd_sc_hd__nor2_1 _26680_ (.A(\inst$top.soc.cpu.gprf.mem[7][30] ),
    .B(net2473),
    .Y(_07364_));
 sky130_fd_sc_hd__o21ai_0 _26681_ (.A1(net2661),
    .A2(\inst$top.soc.cpu.gprf.mem[6][30] ),
    .B1(net2628),
    .Y(_07365_));
 sky130_fd_sc_hd__a22oi_1 _26682_ (.A1(net2514),
    .A2(\inst$top.soc.cpu.gprf.mem[4][30] ),
    .B1(net1953),
    .B2(\inst$top.soc.cpu.gprf.mem[5][30] ),
    .Y(_07366_));
 sky130_fd_sc_hd__o21ai_0 _26683_ (.A1(_07364_),
    .A2(_07365_),
    .B1(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__nand2_1 _26684_ (.A(_07367_),
    .B(net1934),
    .Y(_07368_));
 sky130_fd_sc_hd__nor2_1 _26685_ (.A(\inst$top.soc.cpu.gprf.mem[3][30] ),
    .B(net2473),
    .Y(_07369_));
 sky130_fd_sc_hd__o21ai_0 _26686_ (.A1(net2661),
    .A2(\inst$top.soc.cpu.gprf.mem[2][30] ),
    .B1(net2627),
    .Y(_07370_));
 sky130_fd_sc_hd__a22oi_1 _26687_ (.A1(net2515),
    .A2(\inst$top.soc.cpu.gprf.mem[0][30] ),
    .B1(net1954),
    .B2(\inst$top.soc.cpu.gprf.mem[1][30] ),
    .Y(_07371_));
 sky130_fd_sc_hd__o21ai_0 _26688_ (.A1(_07369_),
    .A2(_07370_),
    .B1(_07371_),
    .Y(_07372_));
 sky130_fd_sc_hd__a21oi_1 _26689_ (.A1(_07372_),
    .A2(net2499),
    .B1(net2592),
    .Y(_07373_));
 sky130_fd_sc_hd__nor2_1 _26690_ (.A(\inst$top.soc.cpu.gprf.mem[23][30] ),
    .B(net2473),
    .Y(_07374_));
 sky130_fd_sc_hd__o21ai_0 _26691_ (.A1(net2662),
    .A2(\inst$top.soc.cpu.gprf.mem[22][30] ),
    .B1(net2627),
    .Y(_07375_));
 sky130_fd_sc_hd__a22oi_1 _26692_ (.A1(net2515),
    .A2(\inst$top.soc.cpu.gprf.mem[20][30] ),
    .B1(net1954),
    .B2(\inst$top.soc.cpu.gprf.mem[21][30] ),
    .Y(_07376_));
 sky130_fd_sc_hd__o21ai_0 _26693_ (.A1(_07374_),
    .A2(_07375_),
    .B1(_07376_),
    .Y(_07377_));
 sky130_fd_sc_hd__nor2_1 _26694_ (.A(\inst$top.soc.cpu.gprf.mem[19][30] ),
    .B(net2473),
    .Y(_07378_));
 sky130_fd_sc_hd__o21ai_0 _26695_ (.A1(net2662),
    .A2(\inst$top.soc.cpu.gprf.mem[18][30] ),
    .B1(net2627),
    .Y(_07379_));
 sky130_fd_sc_hd__a22oi_1 _26696_ (.A1(net2515),
    .A2(\inst$top.soc.cpu.gprf.mem[16][30] ),
    .B1(net1954),
    .B2(\inst$top.soc.cpu.gprf.mem[17][30] ),
    .Y(_07380_));
 sky130_fd_sc_hd__o21ai_0 _26697_ (.A1(_07378_),
    .A2(_07379_),
    .B1(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__a221oi_1 _26698_ (.A1(_07377_),
    .A2(net1934),
    .B1(net2499),
    .B2(_07381_),
    .C1(net2446),
    .Y(_07382_));
 sky130_fd_sc_hd__nor2_1 _26699_ (.A(\inst$top.soc.cpu.gprf.mem[31][30] ),
    .B(net2468),
    .Y(_07383_));
 sky130_fd_sc_hd__o21ai_0 _26700_ (.A1(net2658),
    .A2(\inst$top.soc.cpu.gprf.mem[30][30] ),
    .B1(net2623),
    .Y(_07384_));
 sky130_fd_sc_hd__a221oi_1 _26701_ (.A1(net2511),
    .A2(\inst$top.soc.cpu.gprf.mem[28][30] ),
    .B1(net1950),
    .B2(\inst$top.soc.cpu.gprf.mem[29][30] ),
    .C1(net2453),
    .Y(_07385_));
 sky130_fd_sc_hd__o21ai_0 _26702_ (.A1(_07383_),
    .A2(_07384_),
    .B1(_07385_),
    .Y(_07386_));
 sky130_fd_sc_hd__nor2_1 _26703_ (.A(\inst$top.soc.cpu.gprf.mem[27][30] ),
    .B(net2468),
    .Y(_07387_));
 sky130_fd_sc_hd__o21ai_0 _26704_ (.A1(net2657),
    .A2(\inst$top.soc.cpu.gprf.mem[26][30] ),
    .B1(net2622),
    .Y(_07388_));
 sky130_fd_sc_hd__a221oi_1 _26705_ (.A1(net2512),
    .A2(\inst$top.soc.cpu.gprf.mem[24][30] ),
    .B1(net1952),
    .B2(\inst$top.soc.cpu.gprf.mem[25][30] ),
    .C1(net2609),
    .Y(_07389_));
 sky130_fd_sc_hd__o21ai_0 _26706_ (.A1(_07387_),
    .A2(_07388_),
    .B1(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__nand3_1 _26707_ (.A(_07386_),
    .B(_07390_),
    .C(net2599),
    .Y(_07391_));
 sky130_fd_sc_hd__a32oi_1 _26708_ (.A1(_07363_),
    .A2(_07368_),
    .A3(_07373_),
    .B1(_07382_),
    .B2(_07391_),
    .Y(_00023_));
 sky130_fd_sc_hd__nor2_1 _26709_ (.A(\inst$top.soc.cpu.gprf.mem[31][31] ),
    .B(net2487),
    .Y(_07392_));
 sky130_fd_sc_hd__o21ai_0 _26710_ (.A1(net2672),
    .A2(\inst$top.soc.cpu.gprf.mem[30][31] ),
    .B1(net2645),
    .Y(_07393_));
 sky130_fd_sc_hd__a221oi_1 _26711_ (.A1(net2524),
    .A2(\inst$top.soc.cpu.gprf.mem[28][31] ),
    .B1(net1964),
    .B2(\inst$top.soc.cpu.gprf.mem[29][31] ),
    .C1(net2456),
    .Y(_07394_));
 sky130_fd_sc_hd__o21ai_0 _26712_ (.A1(_07392_),
    .A2(_07393_),
    .B1(_07394_),
    .Y(_07395_));
 sky130_fd_sc_hd__nor2_1 _26713_ (.A(\inst$top.soc.cpu.gprf.mem[27][31] ),
    .B(net2487),
    .Y(_07396_));
 sky130_fd_sc_hd__o21ai_0 _26714_ (.A1(net2672),
    .A2(\inst$top.soc.cpu.gprf.mem[26][31] ),
    .B1(net2642),
    .Y(_07397_));
 sky130_fd_sc_hd__a221oi_1 _26715_ (.A1(net2524),
    .A2(\inst$top.soc.cpu.gprf.mem[24][31] ),
    .B1(net1964),
    .B2(\inst$top.soc.cpu.gprf.mem[25][31] ),
    .C1(net2613),
    .Y(_07398_));
 sky130_fd_sc_hd__o21ai_0 _26716_ (.A1(_07396_),
    .A2(_07397_),
    .B1(_07398_),
    .Y(_07399_));
 sky130_fd_sc_hd__nand3_1 _26717_ (.A(_07395_),
    .B(_07399_),
    .C(net2601),
    .Y(_07400_));
 sky130_fd_sc_hd__nor2_1 _26718_ (.A(\inst$top.soc.cpu.gprf.mem[19][31] ),
    .B(net2487),
    .Y(_07401_));
 sky130_fd_sc_hd__o21ai_0 _26719_ (.A1(net2672),
    .A2(\inst$top.soc.cpu.gprf.mem[18][31] ),
    .B1(net2642),
    .Y(_07402_));
 sky130_fd_sc_hd__a22oi_1 _26720_ (.A1(net2524),
    .A2(\inst$top.soc.cpu.gprf.mem[16][31] ),
    .B1(net1964),
    .B2(\inst$top.soc.cpu.gprf.mem[17][31] ),
    .Y(_07403_));
 sky130_fd_sc_hd__o21ai_0 _26721_ (.A1(_07401_),
    .A2(_07402_),
    .B1(_07403_),
    .Y(_07404_));
 sky130_fd_sc_hd__nand2_1 _26722_ (.A(_07404_),
    .B(net2500),
    .Y(_07405_));
 sky130_fd_sc_hd__nor2_1 _26723_ (.A(\inst$top.soc.cpu.gprf.mem[23][31] ),
    .B(net2487),
    .Y(_07406_));
 sky130_fd_sc_hd__o21ai_0 _26724_ (.A1(net2672),
    .A2(\inst$top.soc.cpu.gprf.mem[22][31] ),
    .B1(net2642),
    .Y(_07407_));
 sky130_fd_sc_hd__a22oi_1 _26725_ (.A1(net2524),
    .A2(\inst$top.soc.cpu.gprf.mem[20][31] ),
    .B1(net1964),
    .B2(\inst$top.soc.cpu.gprf.mem[21][31] ),
    .Y(_07408_));
 sky130_fd_sc_hd__o21ai_0 _26726_ (.A1(_07406_),
    .A2(_07407_),
    .B1(_07408_),
    .Y(_07409_));
 sky130_fd_sc_hd__a21oi_1 _26727_ (.A1(_07409_),
    .A2(net1937),
    .B1(net2447),
    .Y(_07410_));
 sky130_fd_sc_hd__nor2_1 _26728_ (.A(\inst$top.soc.cpu.gprf.mem[3][31] ),
    .B(net2487),
    .Y(_07411_));
 sky130_fd_sc_hd__o21ai_0 _26729_ (.A1(net2672),
    .A2(\inst$top.soc.cpu.gprf.mem[2][31] ),
    .B1(net2642),
    .Y(_07412_));
 sky130_fd_sc_hd__a22oi_1 _26730_ (.A1(net2524),
    .A2(\inst$top.soc.cpu.gprf.mem[0][31] ),
    .B1(net1964),
    .B2(\inst$top.soc.cpu.gprf.mem[1][31] ),
    .Y(_07413_));
 sky130_fd_sc_hd__o21ai_0 _26731_ (.A1(_07411_),
    .A2(_07412_),
    .B1(_07413_),
    .Y(_07414_));
 sky130_fd_sc_hd__nor2_1 _26732_ (.A(\inst$top.soc.cpu.gprf.mem[7][31] ),
    .B(net2487),
    .Y(_07415_));
 sky130_fd_sc_hd__o21ai_0 _26733_ (.A1(net2672),
    .A2(\inst$top.soc.cpu.gprf.mem[6][31] ),
    .B1(net2642),
    .Y(_07416_));
 sky130_fd_sc_hd__a22oi_1 _26734_ (.A1(net2524),
    .A2(\inst$top.soc.cpu.gprf.mem[4][31] ),
    .B1(net1964),
    .B2(\inst$top.soc.cpu.gprf.mem[5][31] ),
    .Y(_07417_));
 sky130_fd_sc_hd__o21ai_0 _26735_ (.A1(_07415_),
    .A2(_07416_),
    .B1(_07417_),
    .Y(_07418_));
 sky130_fd_sc_hd__a221oi_1 _26736_ (.A1(_07414_),
    .A2(net2500),
    .B1(net1937),
    .B2(_07418_),
    .C1(net2594),
    .Y(_07419_));
 sky130_fd_sc_hd__nor2_1 _26737_ (.A(\inst$top.soc.cpu.gprf.mem[15][31] ),
    .B(net2487),
    .Y(_07420_));
 sky130_fd_sc_hd__o21ai_0 _26738_ (.A1(net2672),
    .A2(\inst$top.soc.cpu.gprf.mem[14][31] ),
    .B1(net2642),
    .Y(_07421_));
 sky130_fd_sc_hd__a221oi_1 _26739_ (.A1(net2524),
    .A2(\inst$top.soc.cpu.gprf.mem[12][31] ),
    .B1(net1964),
    .B2(\inst$top.soc.cpu.gprf.mem[13][31] ),
    .C1(net2454),
    .Y(_07422_));
 sky130_fd_sc_hd__o21ai_0 _26740_ (.A1(_07420_),
    .A2(_07421_),
    .B1(_07422_),
    .Y(_07423_));
 sky130_fd_sc_hd__nor2_1 _26741_ (.A(\inst$top.soc.cpu.gprf.mem[11][31] ),
    .B(net2487),
    .Y(_07424_));
 sky130_fd_sc_hd__o21ai_0 _26742_ (.A1(net2672),
    .A2(\inst$top.soc.cpu.gprf.mem[10][31] ),
    .B1(net2642),
    .Y(_07425_));
 sky130_fd_sc_hd__a221oi_1 _26743_ (.A1(net2524),
    .A2(\inst$top.soc.cpu.gprf.mem[8][31] ),
    .B1(net1964),
    .B2(\inst$top.soc.cpu.gprf.mem[9][31] ),
    .C1(net2615),
    .Y(_07426_));
 sky130_fd_sc_hd__o21ai_0 _26744_ (.A1(_07424_),
    .A2(_07425_),
    .B1(_07426_),
    .Y(_07427_));
 sky130_fd_sc_hd__nand3_1 _26745_ (.A(_07423_),
    .B(_07427_),
    .C(net2602),
    .Y(_07428_));
 sky130_fd_sc_hd__a32oi_1 _26746_ (.A1(_07400_),
    .A2(_07405_),
    .A3(_07410_),
    .B1(_07419_),
    .B2(_07428_),
    .Y(_00024_));
 sky130_fd_sc_hd__nand2_1 _26748_ (.A(net2562),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[24] ),
    .Y(_07430_));
 sky130_fd_sc_hd__inv_2 _26749_ (.A(_07430_),
    .Y(\inst$top.soc.bus__dat_w[24] ));
 sky130_fd_sc_hd__nand2_1 _26751_ (.A(net2565),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[16] ),
    .Y(_07432_));
 sky130_fd_sc_hd__inv_2 _26752_ (.A(_07432_),
    .Y(\inst$top.soc.bus__dat_w[16] ));
 sky130_fd_sc_hd__nand2_1 _26754_ (.A(net2562),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[8] ),
    .Y(_07434_));
 sky130_fd_sc_hd__inv_2 _26755_ (.A(_07434_),
    .Y(\inst$top.soc.bus__dat_w[8] ));
 sky130_fd_sc_hd__nand2_1 _26756_ (.A(net2562),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[0] ),
    .Y(_07435_));
 sky130_fd_sc_hd__inv_2 _26757_ (.A(_07435_),
    .Y(\inst$top.soc.bus__dat_w[0] ));
 sky130_fd_sc_hd__nand2_1 _26758_ (.A(net2564),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[25] ),
    .Y(_07436_));
 sky130_fd_sc_hd__inv_2 _26759_ (.A(_07436_),
    .Y(\inst$top.soc.bus__dat_w[25] ));
 sky130_fd_sc_hd__nand2_1 _26760_ (.A(net2564),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[17] ),
    .Y(_07437_));
 sky130_fd_sc_hd__inv_2 _26761_ (.A(_07437_),
    .Y(\inst$top.soc.bus__dat_w[17] ));
 sky130_fd_sc_hd__nand2_1 _26762_ (.A(net2563),
    .B(net3035),
    .Y(_07438_));
 sky130_fd_sc_hd__inv_2 _26763_ (.A(_07438_),
    .Y(\inst$top.soc.bus__dat_w[9] ));
 sky130_fd_sc_hd__nand2_1 _26764_ (.A(net2563),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[1] ),
    .Y(_07439_));
 sky130_fd_sc_hd__inv_2 _26765_ (.A(_07439_),
    .Y(\inst$top.soc.bus__dat_w[1] ));
 sky130_fd_sc_hd__nand2_1 _26766_ (.A(net2563),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[26] ),
    .Y(_07440_));
 sky130_fd_sc_hd__inv_2 _26767_ (.A(_07440_),
    .Y(\inst$top.soc.bus__dat_w[26] ));
 sky130_fd_sc_hd__nand2_1 _26768_ (.A(net2564),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[18] ),
    .Y(_07441_));
 sky130_fd_sc_hd__inv_2 _26769_ (.A(_07441_),
    .Y(\inst$top.soc.bus__dat_w[18] ));
 sky130_fd_sc_hd__nand2_1 _26770_ (.A(net2562),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[10] ),
    .Y(_07442_));
 sky130_fd_sc_hd__inv_2 _26771_ (.A(_07442_),
    .Y(\inst$top.soc.bus__dat_w[10] ));
 sky130_fd_sc_hd__nand2_1 _26772_ (.A(net2563),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[2] ),
    .Y(_07443_));
 sky130_fd_sc_hd__inv_2 _26773_ (.A(_07443_),
    .Y(\inst$top.soc.bus__dat_w[2] ));
 sky130_fd_sc_hd__nand2_1 _26774_ (.A(net2562),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[27] ),
    .Y(_07444_));
 sky130_fd_sc_hd__inv_2 _26775_ (.A(_07444_),
    .Y(\inst$top.soc.bus__dat_w[27] ));
 sky130_fd_sc_hd__nand2_1 _26776_ (.A(net2564),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[19] ),
    .Y(_07445_));
 sky130_fd_sc_hd__inv_2 _26777_ (.A(_07445_),
    .Y(\inst$top.soc.bus__dat_w[19] ));
 sky130_fd_sc_hd__nand2_1 _26778_ (.A(net2563),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[11] ),
    .Y(_07446_));
 sky130_fd_sc_hd__inv_2 _26779_ (.A(_07446_),
    .Y(\inst$top.soc.bus__dat_w[11] ));
 sky130_fd_sc_hd__nand2_1 _26780_ (.A(net2562),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[3] ),
    .Y(_07447_));
 sky130_fd_sc_hd__inv_2 _26781_ (.A(_07447_),
    .Y(\inst$top.soc.bus__dat_w[3] ));
 sky130_fd_sc_hd__nand2_1 _26782_ (.A(net2565),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[28] ),
    .Y(_07448_));
 sky130_fd_sc_hd__inv_2 _26783_ (.A(_07448_),
    .Y(\inst$top.soc.bus__dat_w[28] ));
 sky130_fd_sc_hd__nand2_1 _26784_ (.A(net2564),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[20] ),
    .Y(_07449_));
 sky130_fd_sc_hd__inv_2 _26785_ (.A(_07449_),
    .Y(\inst$top.soc.bus__dat_w[20] ));
 sky130_fd_sc_hd__nand2_1 _26786_ (.A(net2562),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[12] ),
    .Y(_07450_));
 sky130_fd_sc_hd__inv_2 _26787_ (.A(_07450_),
    .Y(\inst$top.soc.bus__dat_w[12] ));
 sky130_fd_sc_hd__nand2_1 _26788_ (.A(net2562),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[4] ),
    .Y(_07451_));
 sky130_fd_sc_hd__inv_2 _26789_ (.A(_07451_),
    .Y(\inst$top.soc.bus__dat_w[4] ));
 sky130_fd_sc_hd__nand2_1 _26790_ (.A(net2565),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[29] ),
    .Y(_07452_));
 sky130_fd_sc_hd__inv_2 _26791_ (.A(_07452_),
    .Y(\inst$top.soc.bus__dat_w[29] ));
 sky130_fd_sc_hd__nand2_1 _26792_ (.A(net2564),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[21] ),
    .Y(_07453_));
 sky130_fd_sc_hd__inv_2 _26793_ (.A(_07453_),
    .Y(\inst$top.soc.bus__dat_w[21] ));
 sky130_fd_sc_hd__nand2_1 _26794_ (.A(net2565),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[13] ),
    .Y(_07454_));
 sky130_fd_sc_hd__inv_2 _26795_ (.A(_07454_),
    .Y(\inst$top.soc.bus__dat_w[13] ));
 sky130_fd_sc_hd__nand2_1 _26796_ (.A(net2562),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[5] ),
    .Y(_07455_));
 sky130_fd_sc_hd__inv_2 _26797_ (.A(_07455_),
    .Y(\inst$top.soc.bus__dat_w[5] ));
 sky130_fd_sc_hd__nand2_1 _26798_ (.A(net2563),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[30] ),
    .Y(_07456_));
 sky130_fd_sc_hd__inv_2 _26799_ (.A(_07456_),
    .Y(\inst$top.soc.bus__dat_w[30] ));
 sky130_fd_sc_hd__nand2_1 _26800_ (.A(net2564),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[22] ),
    .Y(_07457_));
 sky130_fd_sc_hd__inv_2 _26801_ (.A(_07457_),
    .Y(\inst$top.soc.bus__dat_w[22] ));
 sky130_fd_sc_hd__nand2_1 _26802_ (.A(net2563),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[14] ),
    .Y(_07458_));
 sky130_fd_sc_hd__inv_2 _26803_ (.A(_07458_),
    .Y(\inst$top.soc.bus__dat_w[14] ));
 sky130_fd_sc_hd__nand2_1 _26804_ (.A(net2563),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[6] ),
    .Y(_07459_));
 sky130_fd_sc_hd__inv_2 _26805_ (.A(_07459_),
    .Y(\inst$top.soc.bus__dat_w[6] ));
 sky130_fd_sc_hd__nand2_1 _26806_ (.A(net2565),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[31] ),
    .Y(_07460_));
 sky130_fd_sc_hd__inv_2 _26807_ (.A(_07460_),
    .Y(\inst$top.soc.bus__dat_w[31] ));
 sky130_fd_sc_hd__nand2_1 _26808_ (.A(net2564),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[23] ),
    .Y(_07461_));
 sky130_fd_sc_hd__inv_2 _26809_ (.A(_07461_),
    .Y(\inst$top.soc.bus__dat_w[23] ));
 sky130_fd_sc_hd__nand2_1 _26810_ (.A(net2563),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[15] ),
    .Y(_07462_));
 sky130_fd_sc_hd__inv_2 _26811_ (.A(_07462_),
    .Y(\inst$top.soc.bus__dat_w[15] ));
 sky130_fd_sc_hd__nand2_1 _26812_ (.A(net2562),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[7] ),
    .Y(_07463_));
 sky130_fd_sc_hd__inv_2 _26813_ (.A(_07463_),
    .Y(\inst$top.soc.bus__dat_w[7] ));
 sky130_fd_sc_hd__inv_2 _26814_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[0] ),
    .Y(_02710_));
 sky130_fd_sc_hd__inv_1 _26815_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[0] ),
    .Y(_07464_));
 sky130_fd_sc_hd__nor2_1 _26816_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[23] ),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[22] ),
    .Y(_07465_));
 sky130_fd_sc_hd__inv_1 _26817_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[21] ),
    .Y(_07466_));
 sky130_fd_sc_hd__inv_1 _26818_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[20] ),
    .Y(_07467_));
 sky130_fd_sc_hd__nand3_1 _26819_ (.A(_07465_),
    .B(_07466_),
    .C(_07467_),
    .Y(_07468_));
 sky130_fd_sc_hd__nor4_1 _26820_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[13] ),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[12] ),
    .C(\inst$top.soc.uart_0._phy.rx.lower.timer[15] ),
    .D(\inst$top.soc.uart_0._phy.rx.lower.timer[14] ),
    .Y(_07469_));
 sky130_fd_sc_hd__inv_1 _26821_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[9] ),
    .Y(_07470_));
 sky130_fd_sc_hd__inv_1 _26822_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[10] ),
    .Y(_07471_));
 sky130_fd_sc_hd__nand3_1 _26823_ (.A(_07469_),
    .B(_07470_),
    .C(_07471_),
    .Y(_07472_));
 sky130_fd_sc_hd__nor4_1 _26824_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[17] ),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[18] ),
    .C(_07468_),
    .D(_07472_),
    .Y(_07473_));
 sky130_fd_sc_hd__inv_1 _26825_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[8] ),
    .Y(_07474_));
 sky130_fd_sc_hd__inv_1 _26826_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[11] ),
    .Y(_07475_));
 sky130_fd_sc_hd__inv_1 _26827_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[16] ),
    .Y(_07476_));
 sky130_fd_sc_hd__inv_1 _26828_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[19] ),
    .Y(_07477_));
 sky130_fd_sc_hd__nand4_1 _26829_ (.A(_07474_),
    .B(_07475_),
    .C(_07476_),
    .D(_07477_),
    .Y(_07478_));
 sky130_fd_sc_hd__nor4_1 _26830_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[5] ),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[4] ),
    .C(\inst$top.soc.uart_0._phy.rx.lower.timer[7] ),
    .D(\inst$top.soc.uart_0._phy.rx.lower.timer[6] ),
    .Y(_07479_));
 sky130_fd_sc_hd__nor2_1 _26831_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[1] ),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[2] ),
    .Y(_07480_));
 sky130_fd_sc_hd__nand2_1 _26832_ (.A(_07479_),
    .B(_07480_),
    .Y(_07481_));
 sky130_fd_sc_hd__nor4_1 _26833_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[0] ),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[3] ),
    .C(_07478_),
    .D(_07481_),
    .Y(_07482_));
 sky130_fd_sc_hd__nand2_1 _26834_ (.A(_07473_),
    .B(_07482_),
    .Y(_07483_));
 sky130_fd_sc_hd__o21bai_1 _26836_ (.A1(_07464_),
    .A2(net1667),
    .B1_N(\inst$top.soc.uart_0._phy.rx.lower.timer[0] ),
    .Y(_07485_));
 sky130_fd_sc_hd__inv_2 _26837_ (.A(_07485_),
    .Y(_02720_));
 sky130_fd_sc_hd__inv_2 _26838_ (.A(\inst$top.soc.spiflash.ctrl.o_data_count[0] ),
    .Y(_02727_));
 sky130_fd_sc_hd__inv_2 _26839_ (.A(\inst$top.soc.spiflash.ctrl.o_data_count[1] ),
    .Y(_02728_));
 sky130_fd_sc_hd__inv_2 _26840_ (.A(\inst$top.soc.spiflash.ctrl.o_addr_count[0] ),
    .Y(_02723_));
 sky130_fd_sc_hd__inv_2 _26841_ (.A(\inst$top.soc.cpu.divider.quotient[31] ),
    .Y(_02850_));
 sky130_fd_sc_hd__nor2_1 _26845_ (.A(\inst$top.soc.cpu.gprf.mem[7][0] ),
    .B(net2348),
    .Y(_07489_));
 sky130_fd_sc_hd__o21ai_0 _26850_ (.A1(net2751),
    .A2(\inst$top.soc.cpu.gprf.mem[6][0] ),
    .B1(net2724),
    .Y(_07494_));
 sky130_fd_sc_hd__nor2_1 _26854_ (.A(net2754),
    .B(\inst$top.soc.cpu.gprf.mem[4][0] ),
    .Y(_07498_));
 sky130_fd_sc_hd__o21ai_0 _26859_ (.A1(\inst$top.soc.cpu.gprf.mem[5][0] ),
    .A2(net2348),
    .B1(net2322),
    .Y(_07503_));
 sky130_fd_sc_hd__o221ai_1 _26862_ (.A1(_07489_),
    .A2(_07494_),
    .B1(_07498_),
    .B2(_07503_),
    .C1(net2703),
    .Y(_07506_));
 sky130_fd_sc_hd__nor2_1 _26865_ (.A(\inst$top.soc.cpu.gprf.mem[3][0] ),
    .B(net2347),
    .Y(_07509_));
 sky130_fd_sc_hd__o21ai_0 _26869_ (.A1(net2767),
    .A2(\inst$top.soc.cpu.gprf.mem[2][0] ),
    .B1(net2724),
    .Y(_07513_));
 sky130_fd_sc_hd__nor2_1 _26871_ (.A(net2767),
    .B(\inst$top.soc.cpu.gprf.mem[0][0] ),
    .Y(_07515_));
 sky130_fd_sc_hd__o21ai_0 _26874_ (.A1(\inst$top.soc.cpu.gprf.mem[1][0] ),
    .A2(net2347),
    .B1(net2322),
    .Y(_07518_));
 sky130_fd_sc_hd__o221ai_1 _26877_ (.A1(_07509_),
    .A2(_07513_),
    .B1(_07515_),
    .B2(_07518_),
    .C1(net2417),
    .Y(_07521_));
 sky130_fd_sc_hd__nand3_1 _26879_ (.A(_07506_),
    .B(_07521_),
    .C(net2432),
    .Y(_07523_));
 sky130_fd_sc_hd__nor2_1 _26881_ (.A(\inst$top.soc.cpu.gprf.mem[11][0] ),
    .B(net2353),
    .Y(_07525_));
 sky130_fd_sc_hd__o21ai_0 _26885_ (.A1(net2754),
    .A2(\inst$top.soc.cpu.gprf.mem[10][0] ),
    .B1(net2718),
    .Y(_07529_));
 sky130_fd_sc_hd__nor2_1 _26888_ (.A(net2754),
    .B(\inst$top.soc.cpu.gprf.mem[8][0] ),
    .Y(_07532_));
 sky130_fd_sc_hd__o21ai_0 _26892_ (.A1(\inst$top.soc.cpu.gprf.mem[9][0] ),
    .A2(net2354),
    .B1(net2315),
    .Y(_07536_));
 sky130_fd_sc_hd__o221ai_1 _26894_ (.A1(_07525_),
    .A2(_07529_),
    .B1(_07532_),
    .B2(_07536_),
    .C1(net2413),
    .Y(_07538_));
 sky130_fd_sc_hd__nor2_1 _26896_ (.A(\inst$top.soc.cpu.gprf.mem[15][0] ),
    .B(net2351),
    .Y(_07540_));
 sky130_fd_sc_hd__o21ai_0 _26900_ (.A1(net2753),
    .A2(\inst$top.soc.cpu.gprf.mem[14][0] ),
    .B1(net2717),
    .Y(_07544_));
 sky130_fd_sc_hd__nor2_1 _26902_ (.A(net2753),
    .B(\inst$top.soc.cpu.gprf.mem[12][0] ),
    .Y(_07546_));
 sky130_fd_sc_hd__o21ai_0 _26906_ (.A1(\inst$top.soc.cpu.gprf.mem[13][0] ),
    .A2(net2351),
    .B1(net2314),
    .Y(_07550_));
 sky130_fd_sc_hd__o221ai_1 _26908_ (.A1(_07540_),
    .A2(_07544_),
    .B1(_07546_),
    .B2(_07550_),
    .C1(net2700),
    .Y(_07552_));
 sky130_fd_sc_hd__nand3_1 _26910_ (.A(_07538_),
    .B(_07552_),
    .C(net2695),
    .Y(_07554_));
 sky130_fd_sc_hd__nor2_1 _26913_ (.A(\inst$top.soc.cpu.gprf.mem[23][0] ),
    .B(net2353),
    .Y(_07557_));
 sky130_fd_sc_hd__o21ai_0 _26916_ (.A1(net2755),
    .A2(\inst$top.soc.cpu.gprf.mem[22][0] ),
    .B1(net2718),
    .Y(_07560_));
 sky130_fd_sc_hd__nor2_1 _26919_ (.A(net2755),
    .B(\inst$top.soc.cpu.gprf.mem[20][0] ),
    .Y(_07563_));
 sky130_fd_sc_hd__o21ai_0 _26922_ (.A1(\inst$top.soc.cpu.gprf.mem[21][0] ),
    .A2(net2353),
    .B1(net2315),
    .Y(_07566_));
 sky130_fd_sc_hd__o221ai_1 _26924_ (.A1(_07557_),
    .A2(_07560_),
    .B1(_07563_),
    .B2(_07566_),
    .C1(net2701),
    .Y(_07568_));
 sky130_fd_sc_hd__nor2_1 _26926_ (.A(\inst$top.soc.cpu.gprf.mem[19][0] ),
    .B(net2353),
    .Y(_07570_));
 sky130_fd_sc_hd__o21ai_0 _26929_ (.A1(net2755),
    .A2(\inst$top.soc.cpu.gprf.mem[18][0] ),
    .B1(net2718),
    .Y(_07573_));
 sky130_fd_sc_hd__nor2_1 _26932_ (.A(net2755),
    .B(\inst$top.soc.cpu.gprf.mem[16][0] ),
    .Y(_07576_));
 sky130_fd_sc_hd__o21ai_0 _26935_ (.A1(\inst$top.soc.cpu.gprf.mem[17][0] ),
    .A2(net2353),
    .B1(net2315),
    .Y(_07579_));
 sky130_fd_sc_hd__o221ai_1 _26937_ (.A1(_07570_),
    .A2(_07573_),
    .B1(_07576_),
    .B2(_07579_),
    .C1(net2413),
    .Y(_07581_));
 sky130_fd_sc_hd__a31oi_1 _26940_ (.A1(_07568_),
    .A2(_07581_),
    .A3(net2430),
    .B1(net2445),
    .Y(_07584_));
 sky130_fd_sc_hd__nor2_1 _26943_ (.A(\inst$top.soc.cpu.gprf.mem[27][0] ),
    .B(net2353),
    .Y(_07587_));
 sky130_fd_sc_hd__o21ai_0 _26946_ (.A1(net2754),
    .A2(\inst$top.soc.cpu.gprf.mem[26][0] ),
    .B1(net2721),
    .Y(_07590_));
 sky130_fd_sc_hd__nor2_1 _26949_ (.A(net2754),
    .B(\inst$top.soc.cpu.gprf.mem[24][0] ),
    .Y(_07593_));
 sky130_fd_sc_hd__o21ai_0 _26954_ (.A1(\inst$top.soc.cpu.gprf.mem[25][0] ),
    .A2(net2353),
    .B1(net2315),
    .Y(_07598_));
 sky130_fd_sc_hd__o221ai_1 _26956_ (.A1(_07587_),
    .A2(_07590_),
    .B1(_07593_),
    .B2(_07598_),
    .C1(net2413),
    .Y(_07600_));
 sky130_fd_sc_hd__nor2_1 _26958_ (.A(\inst$top.soc.cpu.gprf.mem[31][0] ),
    .B(net2348),
    .Y(_07602_));
 sky130_fd_sc_hd__o21ai_0 _26962_ (.A1(net2754),
    .A2(\inst$top.soc.cpu.gprf.mem[30][0] ),
    .B1(net2721),
    .Y(_07606_));
 sky130_fd_sc_hd__nor2_1 _26965_ (.A(net2754),
    .B(\inst$top.soc.cpu.gprf.mem[28][0] ),
    .Y(_07609_));
 sky130_fd_sc_hd__o21ai_0 _26968_ (.A1(\inst$top.soc.cpu.gprf.mem[29][0] ),
    .A2(net2348),
    .B1(net2322),
    .Y(_07612_));
 sky130_fd_sc_hd__o221ai_1 _26970_ (.A1(_07602_),
    .A2(_07606_),
    .B1(_07609_),
    .B2(_07612_),
    .C1(net2701),
    .Y(_07614_));
 sky130_fd_sc_hd__nand3_1 _26972_ (.A(_07600_),
    .B(_07614_),
    .C(net2695),
    .Y(_07616_));
 sky130_fd_sc_hd__a32oi_1 _26973_ (.A1(_07523_),
    .A2(_07554_),
    .A3(net2445),
    .B1(_07584_),
    .B2(_07616_),
    .Y(_00032_));
 sky130_fd_sc_hd__nor2_1 _26976_ (.A(\inst$top.soc.cpu.gprf.mem[31][1] ),
    .B(net2347),
    .Y(_07619_));
 sky130_fd_sc_hd__o21ai_0 _26978_ (.A1(net2752),
    .A2(\inst$top.soc.cpu.gprf.mem[30][1] ),
    .B1(net2717),
    .Y(_07621_));
 sky130_fd_sc_hd__nor2_1 _26979_ (.A(net2752),
    .B(\inst$top.soc.cpu.gprf.mem[28][1] ),
    .Y(_07622_));
 sky130_fd_sc_hd__o21ai_0 _26982_ (.A1(\inst$top.soc.cpu.gprf.mem[29][1] ),
    .A2(net2348),
    .B1(net2314),
    .Y(_07625_));
 sky130_fd_sc_hd__o221ai_1 _26984_ (.A1(_07619_),
    .A2(_07621_),
    .B1(_07622_),
    .B2(_07625_),
    .C1(net2700),
    .Y(_07627_));
 sky130_fd_sc_hd__nor2_1 _26985_ (.A(\inst$top.soc.cpu.gprf.mem[27][1] ),
    .B(net2350),
    .Y(_07628_));
 sky130_fd_sc_hd__o21ai_0 _26987_ (.A1(net2751),
    .A2(\inst$top.soc.cpu.gprf.mem[26][1] ),
    .B1(net2717),
    .Y(_07630_));
 sky130_fd_sc_hd__nor2_1 _26989_ (.A(net2751),
    .B(\inst$top.soc.cpu.gprf.mem[24][1] ),
    .Y(_07632_));
 sky130_fd_sc_hd__o21ai_0 _26992_ (.A1(\inst$top.soc.cpu.gprf.mem[25][1] ),
    .A2(net2350),
    .B1(net2314),
    .Y(_07635_));
 sky130_fd_sc_hd__o221ai_1 _26994_ (.A1(_07628_),
    .A2(_07630_),
    .B1(_07632_),
    .B2(_07635_),
    .C1(net2413),
    .Y(_07637_));
 sky130_fd_sc_hd__nand3_1 _26995_ (.A(_07627_),
    .B(_07637_),
    .C(net2695),
    .Y(_07638_));
 sky130_fd_sc_hd__nor2_1 _26996_ (.A(\inst$top.soc.cpu.gprf.mem[23][1] ),
    .B(net2351),
    .Y(_07639_));
 sky130_fd_sc_hd__o21ai_0 _26999_ (.A1(net2756),
    .A2(\inst$top.soc.cpu.gprf.mem[22][1] ),
    .B1(net2718),
    .Y(_07642_));
 sky130_fd_sc_hd__nor2_1 _27000_ (.A(net2759),
    .B(\inst$top.soc.cpu.gprf.mem[20][1] ),
    .Y(_07643_));
 sky130_fd_sc_hd__o21ai_0 _27002_ (.A1(\inst$top.soc.cpu.gprf.mem[21][1] ),
    .A2(net2351),
    .B1(net2314),
    .Y(_07645_));
 sky130_fd_sc_hd__o221ai_1 _27004_ (.A1(_07639_),
    .A2(_07642_),
    .B1(_07643_),
    .B2(_07645_),
    .C1(net2700),
    .Y(_07647_));
 sky130_fd_sc_hd__nor2_1 _27005_ (.A(\inst$top.soc.cpu.gprf.mem[19][1] ),
    .B(net2351),
    .Y(_07648_));
 sky130_fd_sc_hd__o21ai_0 _27007_ (.A1(net2757),
    .A2(\inst$top.soc.cpu.gprf.mem[18][1] ),
    .B1(net2717),
    .Y(_07650_));
 sky130_fd_sc_hd__nor2_1 _27009_ (.A(net2757),
    .B(\inst$top.soc.cpu.gprf.mem[16][1] ),
    .Y(_07652_));
 sky130_fd_sc_hd__o21ai_0 _27012_ (.A1(\inst$top.soc.cpu.gprf.mem[17][1] ),
    .A2(net2352),
    .B1(net2315),
    .Y(_07655_));
 sky130_fd_sc_hd__o221ai_1 _27013_ (.A1(_07648_),
    .A2(_07650_),
    .B1(_07652_),
    .B2(_07655_),
    .C1(net2413),
    .Y(_07656_));
 sky130_fd_sc_hd__nand3_1 _27015_ (.A(_07647_),
    .B(_07656_),
    .C(net2430),
    .Y(_07658_));
 sky130_fd_sc_hd__nor2_1 _27017_ (.A(\inst$top.soc.cpu.gprf.mem[11][1] ),
    .B(net2352),
    .Y(_07660_));
 sky130_fd_sc_hd__o21ai_0 _27020_ (.A1(net2757),
    .A2(\inst$top.soc.cpu.gprf.mem[10][1] ),
    .B1(net2719),
    .Y(_07663_));
 sky130_fd_sc_hd__nor2_1 _27021_ (.A(net2757),
    .B(\inst$top.soc.cpu.gprf.mem[8][1] ),
    .Y(_07664_));
 sky130_fd_sc_hd__o21ai_0 _27024_ (.A1(\inst$top.soc.cpu.gprf.mem[9][1] ),
    .A2(net2352),
    .B1(net2315),
    .Y(_07667_));
 sky130_fd_sc_hd__o221ai_1 _27026_ (.A1(_07660_),
    .A2(_07663_),
    .B1(_07664_),
    .B2(_07667_),
    .C1(net2413),
    .Y(_07669_));
 sky130_fd_sc_hd__nor2_1 _27027_ (.A(\inst$top.soc.cpu.gprf.mem[15][1] ),
    .B(net2352),
    .Y(_07670_));
 sky130_fd_sc_hd__o21ai_0 _27028_ (.A1(net2753),
    .A2(\inst$top.soc.cpu.gprf.mem[14][1] ),
    .B1(net2718),
    .Y(_07671_));
 sky130_fd_sc_hd__nor2_1 _27029_ (.A(net2753),
    .B(\inst$top.soc.cpu.gprf.mem[12][1] ),
    .Y(_07672_));
 sky130_fd_sc_hd__o21ai_0 _27032_ (.A1(\inst$top.soc.cpu.gprf.mem[13][1] ),
    .A2(net2352),
    .B1(net2315),
    .Y(_07675_));
 sky130_fd_sc_hd__o221ai_1 _27034_ (.A1(_07670_),
    .A2(_07671_),
    .B1(_07672_),
    .B2(_07675_),
    .C1(net2700),
    .Y(_07677_));
 sky130_fd_sc_hd__nor2_1 _27037_ (.A(\inst$top.soc.cpu.gprf.mem[3][1] ),
    .B(net2348),
    .Y(_07680_));
 sky130_fd_sc_hd__o21ai_0 _27038_ (.A1(net2767),
    .A2(\inst$top.soc.cpu.gprf.mem[2][1] ),
    .B1(net2724),
    .Y(_07681_));
 sky130_fd_sc_hd__nor2_1 _27039_ (.A(net2767),
    .B(\inst$top.soc.cpu.gprf.mem[0][1] ),
    .Y(_07682_));
 sky130_fd_sc_hd__o21ai_0 _27040_ (.A1(\inst$top.soc.cpu.gprf.mem[1][1] ),
    .A2(net2347),
    .B1(net2322),
    .Y(_07683_));
 sky130_fd_sc_hd__o22ai_1 _27041_ (.A1(_07680_),
    .A2(_07681_),
    .B1(_07682_),
    .B2(_07683_),
    .Y(_07684_));
 sky130_fd_sc_hd__nor2_1 _27042_ (.A(\inst$top.soc.cpu.gprf.mem[7][1] ),
    .B(net2347),
    .Y(_07685_));
 sky130_fd_sc_hd__o21ai_0 _27043_ (.A1(net2751),
    .A2(\inst$top.soc.cpu.gprf.mem[6][1] ),
    .B1(net2717),
    .Y(_07686_));
 sky130_fd_sc_hd__nor2_1 _27045_ (.A(net2751),
    .B(\inst$top.soc.cpu.gprf.mem[4][1] ),
    .Y(_07688_));
 sky130_fd_sc_hd__o21ai_0 _27046_ (.A1(\inst$top.soc.cpu.gprf.mem[5][1] ),
    .A2(net2347),
    .B1(net2322),
    .Y(_07689_));
 sky130_fd_sc_hd__o221ai_1 _27047_ (.A1(_07685_),
    .A2(_07686_),
    .B1(_07688_),
    .B2(_07689_),
    .C1(net2700),
    .Y(_07690_));
 sky130_fd_sc_hd__o21ai_0 _27048_ (.A1(net2700),
    .A2(_07684_),
    .B1(_07690_),
    .Y(_07691_));
 sky130_fd_sc_hd__nor2_1 _27049_ (.A(net2695),
    .B(_07691_),
    .Y(_07692_));
 sky130_fd_sc_hd__a311oi_1 _27050_ (.A1(net2695),
    .A2(_07669_),
    .A3(_07677_),
    .B1(net2689),
    .C1(_07692_),
    .Y(_07693_));
 sky130_fd_sc_hd__a31oi_1 _27051_ (.A1(net2689),
    .A2(_07638_),
    .A3(_07658_),
    .B1(_07693_),
    .Y(_00043_));
 sky130_fd_sc_hd__nor2_1 _27052_ (.A(\inst$top.soc.cpu.gprf.mem[23][2] ),
    .B(net2350),
    .Y(_07694_));
 sky130_fd_sc_hd__o21ai_0 _27053_ (.A1(net2753),
    .A2(\inst$top.soc.cpu.gprf.mem[22][2] ),
    .B1(net2717),
    .Y(_07695_));
 sky130_fd_sc_hd__nor2_1 _27054_ (.A(net2753),
    .B(\inst$top.soc.cpu.gprf.mem[20][2] ),
    .Y(_07696_));
 sky130_fd_sc_hd__o21ai_0 _27055_ (.A1(\inst$top.soc.cpu.gprf.mem[21][2] ),
    .A2(net2350),
    .B1(net2314),
    .Y(_07697_));
 sky130_fd_sc_hd__o221ai_1 _27057_ (.A1(_07694_),
    .A2(_07695_),
    .B1(_07696_),
    .B2(_07697_),
    .C1(net2700),
    .Y(_07699_));
 sky130_fd_sc_hd__nor2_1 _27058_ (.A(\inst$top.soc.cpu.gprf.mem[19][2] ),
    .B(net2350),
    .Y(_07700_));
 sky130_fd_sc_hd__o21ai_0 _27059_ (.A1(net2753),
    .A2(\inst$top.soc.cpu.gprf.mem[18][2] ),
    .B1(net2717),
    .Y(_07701_));
 sky130_fd_sc_hd__nor2_1 _27060_ (.A(net2753),
    .B(\inst$top.soc.cpu.gprf.mem[16][2] ),
    .Y(_07702_));
 sky130_fd_sc_hd__o21ai_0 _27061_ (.A1(\inst$top.soc.cpu.gprf.mem[17][2] ),
    .A2(net2350),
    .B1(net2314),
    .Y(_07703_));
 sky130_fd_sc_hd__o221ai_1 _27062_ (.A1(_07700_),
    .A2(_07701_),
    .B1(_07702_),
    .B2(_07703_),
    .C1(net2413),
    .Y(_07704_));
 sky130_fd_sc_hd__nand3_1 _27063_ (.A(_07699_),
    .B(_07704_),
    .C(net2430),
    .Y(_07705_));
 sky130_fd_sc_hd__nor2_1 _27064_ (.A(\inst$top.soc.cpu.gprf.mem[31][2] ),
    .B(net2351),
    .Y(_07706_));
 sky130_fd_sc_hd__o21ai_0 _27065_ (.A1(net2751),
    .A2(\inst$top.soc.cpu.gprf.mem[30][2] ),
    .B1(net2717),
    .Y(_07707_));
 sky130_fd_sc_hd__nor2_1 _27066_ (.A(net2752),
    .B(\inst$top.soc.cpu.gprf.mem[28][2] ),
    .Y(_07708_));
 sky130_fd_sc_hd__o21ai_0 _27068_ (.A1(\inst$top.soc.cpu.gprf.mem[29][2] ),
    .A2(net2351),
    .B1(net2314),
    .Y(_07710_));
 sky130_fd_sc_hd__o221ai_1 _27069_ (.A1(_07706_),
    .A2(_07707_),
    .B1(_07708_),
    .B2(_07710_),
    .C1(net2700),
    .Y(_07711_));
 sky130_fd_sc_hd__nor2_1 _27070_ (.A(\inst$top.soc.cpu.gprf.mem[27][2] ),
    .B(net2351),
    .Y(_07712_));
 sky130_fd_sc_hd__o21ai_0 _27072_ (.A1(net2752),
    .A2(\inst$top.soc.cpu.gprf.mem[26][2] ),
    .B1(net2717),
    .Y(_07714_));
 sky130_fd_sc_hd__nor2_1 _27073_ (.A(net2752),
    .B(\inst$top.soc.cpu.gprf.mem[24][2] ),
    .Y(_07715_));
 sky130_fd_sc_hd__o21ai_0 _27074_ (.A1(\inst$top.soc.cpu.gprf.mem[25][2] ),
    .A2(net2351),
    .B1(net2314),
    .Y(_07716_));
 sky130_fd_sc_hd__o221ai_1 _27076_ (.A1(_07712_),
    .A2(_07714_),
    .B1(_07715_),
    .B2(_07716_),
    .C1(net2413),
    .Y(_07718_));
 sky130_fd_sc_hd__nand3_1 _27077_ (.A(_07711_),
    .B(_07718_),
    .C(net2695),
    .Y(_07719_));
 sky130_fd_sc_hd__nor2_1 _27079_ (.A(\inst$top.soc.cpu.gprf.mem[7][2] ),
    .B(net2347),
    .Y(_07721_));
 sky130_fd_sc_hd__o21ai_0 _27080_ (.A1(net2751),
    .A2(\inst$top.soc.cpu.gprf.mem[6][2] ),
    .B1(net2724),
    .Y(_07722_));
 sky130_fd_sc_hd__nor2_1 _27081_ (.A(net2751),
    .B(\inst$top.soc.cpu.gprf.mem[4][2] ),
    .Y(_07723_));
 sky130_fd_sc_hd__o21ai_0 _27082_ (.A1(\inst$top.soc.cpu.gprf.mem[5][2] ),
    .A2(net2347),
    .B1(net2322),
    .Y(_07724_));
 sky130_fd_sc_hd__o221ai_1 _27083_ (.A1(_07721_),
    .A2(_07722_),
    .B1(_07723_),
    .B2(_07724_),
    .C1(net2703),
    .Y(_07725_));
 sky130_fd_sc_hd__nor2_1 _27085_ (.A(\inst$top.soc.cpu.gprf.mem[3][2] ),
    .B(net2347),
    .Y(_07727_));
 sky130_fd_sc_hd__o21ai_0 _27086_ (.A1(net2767),
    .A2(\inst$top.soc.cpu.gprf.mem[2][2] ),
    .B1(net2724),
    .Y(_07728_));
 sky130_fd_sc_hd__nor2_1 _27087_ (.A(net2767),
    .B(\inst$top.soc.cpu.gprf.mem[0][2] ),
    .Y(_07729_));
 sky130_fd_sc_hd__o21ai_0 _27088_ (.A1(\inst$top.soc.cpu.gprf.mem[1][2] ),
    .A2(net2347),
    .B1(net2322),
    .Y(_07730_));
 sky130_fd_sc_hd__o221ai_1 _27089_ (.A1(_07727_),
    .A2(_07728_),
    .B1(_07729_),
    .B2(_07730_),
    .C1(net2417),
    .Y(_07731_));
 sky130_fd_sc_hd__a31oi_1 _27090_ (.A1(_07725_),
    .A2(_07731_),
    .A3(net2432),
    .B1(net2689),
    .Y(_07732_));
 sky130_fd_sc_hd__nor2_1 _27092_ (.A(\inst$top.soc.cpu.gprf.mem[15][2] ),
    .B(net2350),
    .Y(_07734_));
 sky130_fd_sc_hd__o21ai_0 _27095_ (.A1(net2751),
    .A2(\inst$top.soc.cpu.gprf.mem[14][2] ),
    .B1(net2717),
    .Y(_07737_));
 sky130_fd_sc_hd__nor2_1 _27096_ (.A(net2751),
    .B(\inst$top.soc.cpu.gprf.mem[12][2] ),
    .Y(_07738_));
 sky130_fd_sc_hd__o21ai_0 _27099_ (.A1(\inst$top.soc.cpu.gprf.mem[13][2] ),
    .A2(net2350),
    .B1(net2314),
    .Y(_07741_));
 sky130_fd_sc_hd__o22ai_1 _27100_ (.A1(_07734_),
    .A2(_07737_),
    .B1(_07738_),
    .B2(_07741_),
    .Y(_07742_));
 sky130_fd_sc_hd__nor2_1 _27103_ (.A(\inst$top.soc.cpu.gprf.mem[11][2] ),
    .B(net2350),
    .Y(_07745_));
 sky130_fd_sc_hd__o21ai_0 _27105_ (.A1(net2753),
    .A2(\inst$top.soc.cpu.gprf.mem[10][2] ),
    .B1(net2718),
    .Y(_07747_));
 sky130_fd_sc_hd__nor2_1 _27106_ (.A(net2753),
    .B(\inst$top.soc.cpu.gprf.mem[8][2] ),
    .Y(_07748_));
 sky130_fd_sc_hd__o21ai_0 _27107_ (.A1(\inst$top.soc.cpu.gprf.mem[9][2] ),
    .A2(net2350),
    .B1(net2314),
    .Y(_07749_));
 sky130_fd_sc_hd__o22ai_1 _27108_ (.A1(_07745_),
    .A2(_07747_),
    .B1(_07748_),
    .B2(_07749_),
    .Y(_07750_));
 sky130_fd_sc_hd__nor2_1 _27109_ (.A(net2700),
    .B(_07750_),
    .Y(_07751_));
 sky130_fd_sc_hd__nor2_1 _27110_ (.A(net2430),
    .B(_07751_),
    .Y(_07752_));
 sky130_fd_sc_hd__o21ai_0 _27111_ (.A1(net2413),
    .A2(_07742_),
    .B1(_07752_),
    .Y(_07753_));
 sky130_fd_sc_hd__a32oi_1 _27112_ (.A1(_07705_),
    .A2(_07719_),
    .A3(net2689),
    .B1(_07732_),
    .B2(_07753_),
    .Y(_00054_));
 sky130_fd_sc_hd__nor2_1 _27115_ (.A(\inst$top.soc.cpu.gprf.mem[31][3] ),
    .B(net2389),
    .Y(_07756_));
 sky130_fd_sc_hd__o21ai_0 _27118_ (.A1(net2793),
    .A2(\inst$top.soc.cpu.gprf.mem[30][3] ),
    .B1(net2739),
    .Y(_07759_));
 sky130_fd_sc_hd__nor2_1 _27119_ (.A(net2793),
    .B(\inst$top.soc.cpu.gprf.mem[28][3] ),
    .Y(_07760_));
 sky130_fd_sc_hd__o21ai_0 _27122_ (.A1(\inst$top.soc.cpu.gprf.mem[29][3] ),
    .A2(net2389),
    .B1(net2335),
    .Y(_07763_));
 sky130_fd_sc_hd__o22ai_1 _27123_ (.A1(_07756_),
    .A2(_07759_),
    .B1(_07760_),
    .B2(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__nor2_1 _27127_ (.A(\inst$top.soc.cpu.gprf.mem[27][3] ),
    .B(net2389),
    .Y(_07768_));
 sky130_fd_sc_hd__o21ai_0 _27129_ (.A1(net2797),
    .A2(\inst$top.soc.cpu.gprf.mem[26][3] ),
    .B1(net2740),
    .Y(_07770_));
 sky130_fd_sc_hd__nor2_1 _27131_ (.A(net2797),
    .B(\inst$top.soc.cpu.gprf.mem[24][3] ),
    .Y(_07772_));
 sky130_fd_sc_hd__o21ai_0 _27133_ (.A1(\inst$top.soc.cpu.gprf.mem[25][3] ),
    .A2(net2392),
    .B1(net2336),
    .Y(_07774_));
 sky130_fd_sc_hd__o22ai_1 _27134_ (.A1(_07768_),
    .A2(_07770_),
    .B1(_07772_),
    .B2(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__nor2_1 _27135_ (.A(net2711),
    .B(_07775_),
    .Y(_07776_));
 sky130_fd_sc_hd__nor2_1 _27136_ (.A(net2437),
    .B(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__o21ai_0 _27137_ (.A1(net2423),
    .A2(_07764_),
    .B1(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__nor2_1 _27138_ (.A(\inst$top.soc.cpu.gprf.mem[23][3] ),
    .B(net2390),
    .Y(_07779_));
 sky130_fd_sc_hd__o21ai_0 _27141_ (.A1(net2795),
    .A2(\inst$top.soc.cpu.gprf.mem[22][3] ),
    .B1(net2738),
    .Y(_07782_));
 sky130_fd_sc_hd__nor2_1 _27143_ (.A(net2795),
    .B(\inst$top.soc.cpu.gprf.mem[20][3] ),
    .Y(_07784_));
 sky130_fd_sc_hd__o21ai_0 _27146_ (.A1(\inst$top.soc.cpu.gprf.mem[21][3] ),
    .A2(net2390),
    .B1(net2335),
    .Y(_07787_));
 sky130_fd_sc_hd__o221ai_1 _27148_ (.A1(_07779_),
    .A2(_07782_),
    .B1(_07784_),
    .B2(_07787_),
    .C1(net2712),
    .Y(_07789_));
 sky130_fd_sc_hd__nor2_1 _27149_ (.A(\inst$top.soc.cpu.gprf.mem[19][3] ),
    .B(net2390),
    .Y(_07790_));
 sky130_fd_sc_hd__o21ai_0 _27152_ (.A1(net2794),
    .A2(\inst$top.soc.cpu.gprf.mem[18][3] ),
    .B1(net2738),
    .Y(_07793_));
 sky130_fd_sc_hd__nor2_1 _27154_ (.A(net2795),
    .B(\inst$top.soc.cpu.gprf.mem[16][3] ),
    .Y(_07795_));
 sky130_fd_sc_hd__o21ai_0 _27157_ (.A1(\inst$top.soc.cpu.gprf.mem[17][3] ),
    .A2(net2389),
    .B1(net2335),
    .Y(_07798_));
 sky130_fd_sc_hd__o221ai_1 _27158_ (.A1(_07790_),
    .A2(_07793_),
    .B1(_07795_),
    .B2(_07798_),
    .C1(net2423),
    .Y(_07799_));
 sky130_fd_sc_hd__nand3_1 _27160_ (.A(_07789_),
    .B(_07799_),
    .C(net2437),
    .Y(_07801_));
 sky130_fd_sc_hd__nor2_1 _27161_ (.A(\inst$top.soc.cpu.gprf.mem[7][3] ),
    .B(net2388),
    .Y(_07802_));
 sky130_fd_sc_hd__o21ai_0 _27162_ (.A1(net2793),
    .A2(\inst$top.soc.cpu.gprf.mem[6][3] ),
    .B1(net2737),
    .Y(_07803_));
 sky130_fd_sc_hd__nor2_1 _27163_ (.A(net2793),
    .B(\inst$top.soc.cpu.gprf.mem[4][3] ),
    .Y(_07804_));
 sky130_fd_sc_hd__o21ai_0 _27165_ (.A1(\inst$top.soc.cpu.gprf.mem[5][3] ),
    .A2(net2388),
    .B1(net2334),
    .Y(_07806_));
 sky130_fd_sc_hd__o221ai_1 _27166_ (.A1(_07802_),
    .A2(_07803_),
    .B1(_07804_),
    .B2(_07806_),
    .C1(net2710),
    .Y(_07807_));
 sky130_fd_sc_hd__nor2_1 _27167_ (.A(\inst$top.soc.cpu.gprf.mem[3][3] ),
    .B(net2388),
    .Y(_07808_));
 sky130_fd_sc_hd__o21ai_0 _27168_ (.A1(net2797),
    .A2(\inst$top.soc.cpu.gprf.mem[2][3] ),
    .B1(net2740),
    .Y(_07809_));
 sky130_fd_sc_hd__nor2_1 _27169_ (.A(net2797),
    .B(\inst$top.soc.cpu.gprf.mem[0][3] ),
    .Y(_07810_));
 sky130_fd_sc_hd__o21ai_0 _27170_ (.A1(\inst$top.soc.cpu.gprf.mem[1][3] ),
    .A2(net2388),
    .B1(net2334),
    .Y(_07811_));
 sky130_fd_sc_hd__o221ai_1 _27171_ (.A1(_07808_),
    .A2(_07809_),
    .B1(_07810_),
    .B2(_07811_),
    .C1(net2423),
    .Y(_07812_));
 sky130_fd_sc_hd__a31oi_1 _27172_ (.A1(_07807_),
    .A2(_07812_),
    .A3(net2437),
    .B1(net2692),
    .Y(_07813_));
 sky130_fd_sc_hd__nor2_1 _27173_ (.A(\inst$top.soc.cpu.gprf.mem[15][3] ),
    .B(net2388),
    .Y(_07814_));
 sky130_fd_sc_hd__o21ai_0 _27174_ (.A1(net2793),
    .A2(\inst$top.soc.cpu.gprf.mem[14][3] ),
    .B1(net2737),
    .Y(_07815_));
 sky130_fd_sc_hd__nor2_1 _27175_ (.A(net2793),
    .B(\inst$top.soc.cpu.gprf.mem[12][3] ),
    .Y(_07816_));
 sky130_fd_sc_hd__o21ai_0 _27176_ (.A1(\inst$top.soc.cpu.gprf.mem[13][3] ),
    .A2(net2388),
    .B1(net2335),
    .Y(_07817_));
 sky130_fd_sc_hd__o22ai_1 _27177_ (.A1(_07814_),
    .A2(_07815_),
    .B1(_07816_),
    .B2(_07817_),
    .Y(_07818_));
 sky130_fd_sc_hd__nor2_1 _27178_ (.A(\inst$top.soc.cpu.gprf.mem[11][3] ),
    .B(net2388),
    .Y(_07819_));
 sky130_fd_sc_hd__o21ai_0 _27179_ (.A1(net2793),
    .A2(\inst$top.soc.cpu.gprf.mem[10][3] ),
    .B1(net2737),
    .Y(_07820_));
 sky130_fd_sc_hd__nor2_1 _27180_ (.A(net2793),
    .B(\inst$top.soc.cpu.gprf.mem[8][3] ),
    .Y(_07821_));
 sky130_fd_sc_hd__o21ai_0 _27181_ (.A1(\inst$top.soc.cpu.gprf.mem[9][3] ),
    .A2(net2388),
    .B1(net2335),
    .Y(_07822_));
 sky130_fd_sc_hd__o22ai_1 _27182_ (.A1(_07819_),
    .A2(_07820_),
    .B1(_07821_),
    .B2(_07822_),
    .Y(_07823_));
 sky130_fd_sc_hd__nor2_1 _27183_ (.A(net2710),
    .B(_07823_),
    .Y(_07824_));
 sky130_fd_sc_hd__nor2_1 _27184_ (.A(net2437),
    .B(_07824_),
    .Y(_07825_));
 sky130_fd_sc_hd__o21ai_0 _27185_ (.A1(net2423),
    .A2(_07818_),
    .B1(_07825_),
    .Y(_07826_));
 sky130_fd_sc_hd__a32oi_1 _27186_ (.A1(net2691),
    .A2(_07778_),
    .A3(_07801_),
    .B1(_07813_),
    .B2(_07826_),
    .Y(_00057_));
 sky130_fd_sc_hd__nor2_1 _27187_ (.A(\inst$top.soc.cpu.gprf.mem[31][4] ),
    .B(net2355),
    .Y(_07827_));
 sky130_fd_sc_hd__o21ai_0 _27188_ (.A1(net2758),
    .A2(\inst$top.soc.cpu.gprf.mem[30][4] ),
    .B1(net2719),
    .Y(_07828_));
 sky130_fd_sc_hd__nor2_1 _27189_ (.A(net2757),
    .B(\inst$top.soc.cpu.gprf.mem[28][4] ),
    .Y(_07829_));
 sky130_fd_sc_hd__o21ai_0 _27190_ (.A1(\inst$top.soc.cpu.gprf.mem[29][4] ),
    .A2(net2355),
    .B1(net2316),
    .Y(_07830_));
 sky130_fd_sc_hd__o221ai_1 _27191_ (.A1(_07827_),
    .A2(_07828_),
    .B1(_07829_),
    .B2(_07830_),
    .C1(net2701),
    .Y(_07831_));
 sky130_fd_sc_hd__nor2_1 _27192_ (.A(\inst$top.soc.cpu.gprf.mem[27][4] ),
    .B(net2355),
    .Y(_07832_));
 sky130_fd_sc_hd__o21ai_0 _27193_ (.A1(net2757),
    .A2(\inst$top.soc.cpu.gprf.mem[26][4] ),
    .B1(net2719),
    .Y(_07833_));
 sky130_fd_sc_hd__nor2_1 _27194_ (.A(net2757),
    .B(\inst$top.soc.cpu.gprf.mem[24][4] ),
    .Y(_07834_));
 sky130_fd_sc_hd__o21ai_0 _27195_ (.A1(\inst$top.soc.cpu.gprf.mem[25][4] ),
    .A2(net2355),
    .B1(net2316),
    .Y(_07835_));
 sky130_fd_sc_hd__o221ai_1 _27196_ (.A1(_07832_),
    .A2(_07833_),
    .B1(_07834_),
    .B2(_07835_),
    .C1(net2414),
    .Y(_07836_));
 sky130_fd_sc_hd__nand3_1 _27197_ (.A(_07831_),
    .B(_07836_),
    .C(net2695),
    .Y(_07837_));
 sky130_fd_sc_hd__nor2_1 _27198_ (.A(\inst$top.soc.cpu.gprf.mem[23][4] ),
    .B(net2356),
    .Y(_07838_));
 sky130_fd_sc_hd__o21ai_0 _27199_ (.A1(net2759),
    .A2(\inst$top.soc.cpu.gprf.mem[22][4] ),
    .B1(net2719),
    .Y(_07839_));
 sky130_fd_sc_hd__nor2_1 _27200_ (.A(net2758),
    .B(\inst$top.soc.cpu.gprf.mem[20][4] ),
    .Y(_07840_));
 sky130_fd_sc_hd__o21ai_0 _27201_ (.A1(\inst$top.soc.cpu.gprf.mem[21][4] ),
    .A2(net2356),
    .B1(net2316),
    .Y(_07841_));
 sky130_fd_sc_hd__o221ai_1 _27202_ (.A1(_07838_),
    .A2(_07839_),
    .B1(_07840_),
    .B2(_07841_),
    .C1(net2701),
    .Y(_07842_));
 sky130_fd_sc_hd__nor2_1 _27203_ (.A(\inst$top.soc.cpu.gprf.mem[19][4] ),
    .B(net2356),
    .Y(_07843_));
 sky130_fd_sc_hd__o21ai_0 _27204_ (.A1(net2758),
    .A2(\inst$top.soc.cpu.gprf.mem[18][4] ),
    .B1(net2719),
    .Y(_07844_));
 sky130_fd_sc_hd__nor2_1 _27205_ (.A(net2758),
    .B(\inst$top.soc.cpu.gprf.mem[16][4] ),
    .Y(_07845_));
 sky130_fd_sc_hd__o21ai_0 _27206_ (.A1(\inst$top.soc.cpu.gprf.mem[17][4] ),
    .A2(net2356),
    .B1(net2316),
    .Y(_07846_));
 sky130_fd_sc_hd__o221ai_1 _27207_ (.A1(_07843_),
    .A2(_07844_),
    .B1(_07845_),
    .B2(_07846_),
    .C1(net2414),
    .Y(_07847_));
 sky130_fd_sc_hd__nand3_1 _27208_ (.A(_07842_),
    .B(_07847_),
    .C(net2430),
    .Y(_07848_));
 sky130_fd_sc_hd__nor2_1 _27211_ (.A(\inst$top.soc.cpu.gprf.mem[3][4] ),
    .B(net2355),
    .Y(_07851_));
 sky130_fd_sc_hd__o21ai_0 _27213_ (.A1(net2758),
    .A2(\inst$top.soc.cpu.gprf.mem[2][4] ),
    .B1(net2719),
    .Y(_07853_));
 sky130_fd_sc_hd__nor2_1 _27214_ (.A(net2758),
    .B(\inst$top.soc.cpu.gprf.mem[0][4] ),
    .Y(_07854_));
 sky130_fd_sc_hd__o21ai_0 _27216_ (.A1(\inst$top.soc.cpu.gprf.mem[1][4] ),
    .A2(net2355),
    .B1(net2316),
    .Y(_07856_));
 sky130_fd_sc_hd__o22ai_1 _27217_ (.A1(_07851_),
    .A2(_07853_),
    .B1(_07854_),
    .B2(_07856_),
    .Y(_07857_));
 sky130_fd_sc_hd__nor2_1 _27218_ (.A(net2701),
    .B(_07857_),
    .Y(_07858_));
 sky130_fd_sc_hd__nor2_1 _27220_ (.A(\inst$top.soc.cpu.gprf.mem[7][4] ),
    .B(net2355),
    .Y(_07860_));
 sky130_fd_sc_hd__o21ai_0 _27222_ (.A1(net2757),
    .A2(\inst$top.soc.cpu.gprf.mem[6][4] ),
    .B1(net2719),
    .Y(_07862_));
 sky130_fd_sc_hd__nor2_1 _27224_ (.A(net2758),
    .B(\inst$top.soc.cpu.gprf.mem[4][4] ),
    .Y(_07864_));
 sky130_fd_sc_hd__o21ai_0 _27226_ (.A1(\inst$top.soc.cpu.gprf.mem[5][4] ),
    .A2(net2355),
    .B1(net2316),
    .Y(_07866_));
 sky130_fd_sc_hd__o22ai_1 _27227_ (.A1(_07860_),
    .A2(_07862_),
    .B1(_07864_),
    .B2(_07866_),
    .Y(_07867_));
 sky130_fd_sc_hd__o21ai_0 _27229_ (.A1(net2414),
    .A2(_07867_),
    .B1(net2431),
    .Y(_07869_));
 sky130_fd_sc_hd__nor2_1 _27230_ (.A(\inst$top.soc.cpu.gprf.mem[11][4] ),
    .B(net2356),
    .Y(_07870_));
 sky130_fd_sc_hd__o21ai_0 _27232_ (.A1(net2768),
    .A2(\inst$top.soc.cpu.gprf.mem[10][4] ),
    .B1(net2725),
    .Y(_07872_));
 sky130_fd_sc_hd__nor2_1 _27233_ (.A(net2768),
    .B(\inst$top.soc.cpu.gprf.mem[8][4] ),
    .Y(_07873_));
 sky130_fd_sc_hd__o21ai_0 _27234_ (.A1(\inst$top.soc.cpu.gprf.mem[9][4] ),
    .A2(net2356),
    .B1(net2316),
    .Y(_07874_));
 sky130_fd_sc_hd__o221ai_1 _27235_ (.A1(_07870_),
    .A2(_07872_),
    .B1(_07873_),
    .B2(_07874_),
    .C1(net2414),
    .Y(_07875_));
 sky130_fd_sc_hd__nor2_1 _27236_ (.A(\inst$top.soc.cpu.gprf.mem[15][4] ),
    .B(net2356),
    .Y(_07876_));
 sky130_fd_sc_hd__o21ai_0 _27237_ (.A1(net2758),
    .A2(\inst$top.soc.cpu.gprf.mem[14][4] ),
    .B1(net2719),
    .Y(_07877_));
 sky130_fd_sc_hd__nor2_1 _27238_ (.A(net2758),
    .B(\inst$top.soc.cpu.gprf.mem[12][4] ),
    .Y(_07878_));
 sky130_fd_sc_hd__o21ai_0 _27240_ (.A1(\inst$top.soc.cpu.gprf.mem[13][4] ),
    .A2(net2356),
    .B1(net2317),
    .Y(_07880_));
 sky130_fd_sc_hd__o221ai_1 _27241_ (.A1(_07876_),
    .A2(_07877_),
    .B1(_07878_),
    .B2(_07880_),
    .C1(net2702),
    .Y(_07881_));
 sky130_fd_sc_hd__nand3_1 _27242_ (.A(_07875_),
    .B(_07881_),
    .C(net2697),
    .Y(_07882_));
 sky130_fd_sc_hd__o21ai_0 _27243_ (.A1(_07858_),
    .A2(_07869_),
    .B1(_07882_),
    .Y(_07883_));
 sky130_fd_sc_hd__nor2_1 _27244_ (.A(net2689),
    .B(_07883_),
    .Y(_07884_));
 sky130_fd_sc_hd__a31oi_1 _27245_ (.A1(net2689),
    .A2(_07837_),
    .A3(_07848_),
    .B1(_07884_),
    .Y(_00058_));
 sky130_fd_sc_hd__nor2_1 _27246_ (.A(\inst$top.soc.cpu.gprf.mem[31][5] ),
    .B(net2371),
    .Y(_07885_));
 sky130_fd_sc_hd__o21ai_0 _27248_ (.A1(net2776),
    .A2(\inst$top.soc.cpu.gprf.mem[30][5] ),
    .B1(net2730),
    .Y(_07887_));
 sky130_fd_sc_hd__nor2_1 _27249_ (.A(net2775),
    .B(\inst$top.soc.cpu.gprf.mem[28][5] ),
    .Y(_07888_));
 sky130_fd_sc_hd__o21ai_0 _27250_ (.A1(\inst$top.soc.cpu.gprf.mem[29][5] ),
    .A2(net2375),
    .B1(net2326),
    .Y(_07889_));
 sky130_fd_sc_hd__o22ai_1 _27251_ (.A1(_07885_),
    .A2(_07887_),
    .B1(_07888_),
    .B2(_07889_),
    .Y(_07890_));
 sky130_fd_sc_hd__nor2_1 _27252_ (.A(\inst$top.soc.cpu.gprf.mem[27][5] ),
    .B(net2375),
    .Y(_07891_));
 sky130_fd_sc_hd__o21ai_0 _27253_ (.A1(net2775),
    .A2(\inst$top.soc.cpu.gprf.mem[26][5] ),
    .B1(net2730),
    .Y(_07892_));
 sky130_fd_sc_hd__nor2_1 _27254_ (.A(net2776),
    .B(\inst$top.soc.cpu.gprf.mem[24][5] ),
    .Y(_07893_));
 sky130_fd_sc_hd__o21ai_0 _27255_ (.A1(\inst$top.soc.cpu.gprf.mem[25][5] ),
    .A2(net2371),
    .B1(net2328),
    .Y(_07894_));
 sky130_fd_sc_hd__o22ai_1 _27256_ (.A1(_07891_),
    .A2(_07892_),
    .B1(_07893_),
    .B2(_07894_),
    .Y(_07895_));
 sky130_fd_sc_hd__nor2_1 _27257_ (.A(net2705),
    .B(_07895_),
    .Y(_07896_));
 sky130_fd_sc_hd__nor2_1 _27258_ (.A(net2434),
    .B(_07896_),
    .Y(_07897_));
 sky130_fd_sc_hd__o21ai_0 _27259_ (.A1(net2419),
    .A2(_07890_),
    .B1(_07897_),
    .Y(_07898_));
 sky130_fd_sc_hd__nor2_1 _27260_ (.A(\inst$top.soc.cpu.gprf.mem[23][5] ),
    .B(net2374),
    .Y(_07899_));
 sky130_fd_sc_hd__o21ai_0 _27261_ (.A1(net2778),
    .A2(\inst$top.soc.cpu.gprf.mem[22][5] ),
    .B1(net2729),
    .Y(_07900_));
 sky130_fd_sc_hd__nor2_1 _27262_ (.A(net2778),
    .B(\inst$top.soc.cpu.gprf.mem[20][5] ),
    .Y(_07901_));
 sky130_fd_sc_hd__o21ai_0 _27263_ (.A1(\inst$top.soc.cpu.gprf.mem[21][5] ),
    .A2(net2374),
    .B1(net2327),
    .Y(_07902_));
 sky130_fd_sc_hd__o221ai_1 _27264_ (.A1(_07899_),
    .A2(_07900_),
    .B1(_07901_),
    .B2(_07902_),
    .C1(net2706),
    .Y(_07903_));
 sky130_fd_sc_hd__nor2_1 _27266_ (.A(\inst$top.soc.cpu.gprf.mem[19][5] ),
    .B(net2374),
    .Y(_07905_));
 sky130_fd_sc_hd__o21ai_0 _27267_ (.A1(net2778),
    .A2(\inst$top.soc.cpu.gprf.mem[18][5] ),
    .B1(net2730),
    .Y(_07906_));
 sky130_fd_sc_hd__nor2_1 _27268_ (.A(net2778),
    .B(\inst$top.soc.cpu.gprf.mem[16][5] ),
    .Y(_07907_));
 sky130_fd_sc_hd__o21ai_0 _27269_ (.A1(\inst$top.soc.cpu.gprf.mem[17][5] ),
    .A2(net2374),
    .B1(net2327),
    .Y(_07908_));
 sky130_fd_sc_hd__o221ai_1 _27271_ (.A1(_07905_),
    .A2(_07906_),
    .B1(_07907_),
    .B2(_07908_),
    .C1(net2419),
    .Y(_07910_));
 sky130_fd_sc_hd__nand3_1 _27272_ (.A(_07903_),
    .B(_07910_),
    .C(net2434),
    .Y(_07911_));
 sky130_fd_sc_hd__nor2_1 _27273_ (.A(\inst$top.soc.cpu.gprf.mem[7][5] ),
    .B(net2371),
    .Y(_07912_));
 sky130_fd_sc_hd__o21ai_0 _27275_ (.A1(net2775),
    .A2(\inst$top.soc.cpu.gprf.mem[6][5] ),
    .B1(net2728),
    .Y(_07914_));
 sky130_fd_sc_hd__nor2_1 _27276_ (.A(net2775),
    .B(\inst$top.soc.cpu.gprf.mem[4][5] ),
    .Y(_07915_));
 sky130_fd_sc_hd__o21ai_0 _27277_ (.A1(\inst$top.soc.cpu.gprf.mem[5][5] ),
    .A2(net2371),
    .B1(net2326),
    .Y(_07916_));
 sky130_fd_sc_hd__o221ai_1 _27278_ (.A1(_07912_),
    .A2(_07914_),
    .B1(_07915_),
    .B2(_07916_),
    .C1(net2705),
    .Y(_07917_));
 sky130_fd_sc_hd__nor2_1 _27279_ (.A(\inst$top.soc.cpu.gprf.mem[3][5] ),
    .B(net2371),
    .Y(_07918_));
 sky130_fd_sc_hd__o21ai_0 _27281_ (.A1(net2775),
    .A2(\inst$top.soc.cpu.gprf.mem[2][5] ),
    .B1(net2730),
    .Y(_07920_));
 sky130_fd_sc_hd__nor2_1 _27282_ (.A(net2775),
    .B(\inst$top.soc.cpu.gprf.mem[0][5] ),
    .Y(_07921_));
 sky130_fd_sc_hd__o21ai_0 _27283_ (.A1(\inst$top.soc.cpu.gprf.mem[1][5] ),
    .A2(net2371),
    .B1(net2326),
    .Y(_07922_));
 sky130_fd_sc_hd__o221ai_1 _27284_ (.A1(_07918_),
    .A2(_07920_),
    .B1(_07921_),
    .B2(_07922_),
    .C1(net2419),
    .Y(_07923_));
 sky130_fd_sc_hd__a31oi_1 _27285_ (.A1(_07917_),
    .A2(_07923_),
    .A3(net2433),
    .B1(net2691),
    .Y(_07924_));
 sky130_fd_sc_hd__nor2_1 _27286_ (.A(\inst$top.soc.cpu.gprf.mem[15][5] ),
    .B(net2371),
    .Y(_07925_));
 sky130_fd_sc_hd__o21ai_0 _27287_ (.A1(net2775),
    .A2(\inst$top.soc.cpu.gprf.mem[14][5] ),
    .B1(net2728),
    .Y(_07926_));
 sky130_fd_sc_hd__nor2_1 _27288_ (.A(net2775),
    .B(\inst$top.soc.cpu.gprf.mem[12][5] ),
    .Y(_07927_));
 sky130_fd_sc_hd__o21ai_0 _27289_ (.A1(\inst$top.soc.cpu.gprf.mem[13][5] ),
    .A2(net2371),
    .B1(net2326),
    .Y(_07928_));
 sky130_fd_sc_hd__o22ai_1 _27290_ (.A1(_07925_),
    .A2(_07926_),
    .B1(_07927_),
    .B2(_07928_),
    .Y(_07929_));
 sky130_fd_sc_hd__nor2_1 _27291_ (.A(\inst$top.soc.cpu.gprf.mem[11][5] ),
    .B(net2371),
    .Y(_07930_));
 sky130_fd_sc_hd__o21ai_0 _27292_ (.A1(net2775),
    .A2(\inst$top.soc.cpu.gprf.mem[10][5] ),
    .B1(net2728),
    .Y(_07931_));
 sky130_fd_sc_hd__nor2_1 _27293_ (.A(net2775),
    .B(\inst$top.soc.cpu.gprf.mem[8][5] ),
    .Y(_07932_));
 sky130_fd_sc_hd__o21ai_0 _27294_ (.A1(\inst$top.soc.cpu.gprf.mem[9][5] ),
    .A2(net2371),
    .B1(net2326),
    .Y(_07933_));
 sky130_fd_sc_hd__o22ai_1 _27295_ (.A1(_07930_),
    .A2(_07931_),
    .B1(_07932_),
    .B2(_07933_),
    .Y(_07934_));
 sky130_fd_sc_hd__nor2_1 _27296_ (.A(net2705),
    .B(_07934_),
    .Y(_07935_));
 sky130_fd_sc_hd__nor2_1 _27297_ (.A(net2433),
    .B(_07935_),
    .Y(_07936_));
 sky130_fd_sc_hd__o21ai_0 _27298_ (.A1(net2419),
    .A2(_07929_),
    .B1(_07936_),
    .Y(_07937_));
 sky130_fd_sc_hd__a32oi_1 _27299_ (.A1(net2691),
    .A2(_07898_),
    .A3(_07911_),
    .B1(_07924_),
    .B2(_07937_),
    .Y(_00059_));
 sky130_fd_sc_hd__nor2_1 _27300_ (.A(\inst$top.soc.cpu.gprf.mem[31][6] ),
    .B(net2366),
    .Y(_07938_));
 sky130_fd_sc_hd__o21ai_0 _27301_ (.A1(net2776),
    .A2(\inst$top.soc.cpu.gprf.mem[30][6] ),
    .B1(net2728),
    .Y(_07939_));
 sky130_fd_sc_hd__nor2_1 _27302_ (.A(net2776),
    .B(\inst$top.soc.cpu.gprf.mem[28][6] ),
    .Y(_07940_));
 sky130_fd_sc_hd__o21ai_0 _27303_ (.A1(\inst$top.soc.cpu.gprf.mem[29][6] ),
    .A2(net2366),
    .B1(net2323),
    .Y(_07941_));
 sky130_fd_sc_hd__o22ai_1 _27304_ (.A1(_07938_),
    .A2(_07939_),
    .B1(_07940_),
    .B2(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__nor2_1 _27305_ (.A(\inst$top.soc.cpu.gprf.mem[27][6] ),
    .B(net2372),
    .Y(_07943_));
 sky130_fd_sc_hd__o21ai_0 _27306_ (.A1(net2774),
    .A2(\inst$top.soc.cpu.gprf.mem[26][6] ),
    .B1(net2728),
    .Y(_07944_));
 sky130_fd_sc_hd__nor2_1 _27307_ (.A(net2774),
    .B(\inst$top.soc.cpu.gprf.mem[24][6] ),
    .Y(_07945_));
 sky130_fd_sc_hd__o21ai_0 _27308_ (.A1(\inst$top.soc.cpu.gprf.mem[25][6] ),
    .A2(net2372),
    .B1(net2326),
    .Y(_07946_));
 sky130_fd_sc_hd__o22ai_1 _27309_ (.A1(_07943_),
    .A2(_07944_),
    .B1(_07945_),
    .B2(_07946_),
    .Y(_07947_));
 sky130_fd_sc_hd__nor2_1 _27310_ (.A(net2705),
    .B(_07947_),
    .Y(_07948_));
 sky130_fd_sc_hd__nor2_1 _27311_ (.A(net2434),
    .B(_07948_),
    .Y(_07949_));
 sky130_fd_sc_hd__o21ai_0 _27312_ (.A1(net2419),
    .A2(_07942_),
    .B1(_07949_),
    .Y(_07950_));
 sky130_fd_sc_hd__nor2_1 _27314_ (.A(\inst$top.soc.cpu.gprf.mem[23][6] ),
    .B(net2372),
    .Y(_07952_));
 sky130_fd_sc_hd__o21ai_0 _27315_ (.A1(net2776),
    .A2(\inst$top.soc.cpu.gprf.mem[22][6] ),
    .B1(net2728),
    .Y(_07953_));
 sky130_fd_sc_hd__nor2_1 _27316_ (.A(net2776),
    .B(\inst$top.soc.cpu.gprf.mem[20][6] ),
    .Y(_07954_));
 sky130_fd_sc_hd__o21ai_0 _27317_ (.A1(\inst$top.soc.cpu.gprf.mem[21][6] ),
    .A2(net2372),
    .B1(net2326),
    .Y(_07955_));
 sky130_fd_sc_hd__o221ai_1 _27318_ (.A1(_07952_),
    .A2(_07953_),
    .B1(_07954_),
    .B2(_07955_),
    .C1(net2705),
    .Y(_07956_));
 sky130_fd_sc_hd__nor2_1 _27319_ (.A(\inst$top.soc.cpu.gprf.mem[19][6] ),
    .B(net2372),
    .Y(_07957_));
 sky130_fd_sc_hd__o21ai_0 _27320_ (.A1(net2774),
    .A2(\inst$top.soc.cpu.gprf.mem[18][6] ),
    .B1(net2728),
    .Y(_07958_));
 sky130_fd_sc_hd__nor2_1 _27321_ (.A(net2774),
    .B(\inst$top.soc.cpu.gprf.mem[16][6] ),
    .Y(_07959_));
 sky130_fd_sc_hd__o21ai_0 _27323_ (.A1(\inst$top.soc.cpu.gprf.mem[17][6] ),
    .A2(net2372),
    .B1(net2326),
    .Y(_07961_));
 sky130_fd_sc_hd__o221ai_1 _27324_ (.A1(_07957_),
    .A2(_07958_),
    .B1(_07959_),
    .B2(_07961_),
    .C1(net2419),
    .Y(_07962_));
 sky130_fd_sc_hd__nand3_1 _27325_ (.A(_07956_),
    .B(_07962_),
    .C(net2434),
    .Y(_07963_));
 sky130_fd_sc_hd__nor2_1 _27327_ (.A(\inst$top.soc.cpu.gprf.mem[7][6] ),
    .B(net2366),
    .Y(_07965_));
 sky130_fd_sc_hd__o21ai_0 _27329_ (.A1(net2774),
    .A2(\inst$top.soc.cpu.gprf.mem[6][6] ),
    .B1(net2728),
    .Y(_07967_));
 sky130_fd_sc_hd__nor2_1 _27331_ (.A(net2769),
    .B(\inst$top.soc.cpu.gprf.mem[4][6] ),
    .Y(_07969_));
 sky130_fd_sc_hd__o21ai_0 _27332_ (.A1(\inst$top.soc.cpu.gprf.mem[5][6] ),
    .A2(net2366),
    .B1(net2323),
    .Y(_07970_));
 sky130_fd_sc_hd__o221ai_1 _27333_ (.A1(_07965_),
    .A2(_07967_),
    .B1(_07969_),
    .B2(_07970_),
    .C1(net2704),
    .Y(_07971_));
 sky130_fd_sc_hd__nor2_1 _27334_ (.A(\inst$top.soc.cpu.gprf.mem[3][6] ),
    .B(net2366),
    .Y(_07972_));
 sky130_fd_sc_hd__o21ai_0 _27335_ (.A1(net2769),
    .A2(\inst$top.soc.cpu.gprf.mem[2][6] ),
    .B1(net2727),
    .Y(_07973_));
 sky130_fd_sc_hd__nor2_1 _27336_ (.A(net2774),
    .B(\inst$top.soc.cpu.gprf.mem[0][6] ),
    .Y(_07974_));
 sky130_fd_sc_hd__o21ai_0 _27337_ (.A1(\inst$top.soc.cpu.gprf.mem[1][6] ),
    .A2(net2366),
    .B1(net2323),
    .Y(_07975_));
 sky130_fd_sc_hd__o221ai_1 _27338_ (.A1(_07972_),
    .A2(_07973_),
    .B1(_07974_),
    .B2(_07975_),
    .C1(net2418),
    .Y(_07976_));
 sky130_fd_sc_hd__a31oi_1 _27340_ (.A1(_07971_),
    .A2(_07976_),
    .A3(net2433),
    .B1(net2694),
    .Y(_07978_));
 sky130_fd_sc_hd__nor2_1 _27341_ (.A(\inst$top.soc.cpu.gprf.mem[15][6] ),
    .B(net2372),
    .Y(_07979_));
 sky130_fd_sc_hd__o21ai_0 _27342_ (.A1(net2774),
    .A2(\inst$top.soc.cpu.gprf.mem[14][6] ),
    .B1(net2728),
    .Y(_07980_));
 sky130_fd_sc_hd__nor2_1 _27343_ (.A(net2774),
    .B(\inst$top.soc.cpu.gprf.mem[12][6] ),
    .Y(_07981_));
 sky130_fd_sc_hd__o21ai_0 _27344_ (.A1(\inst$top.soc.cpu.gprf.mem[13][6] ),
    .A2(net2372),
    .B1(net2326),
    .Y(_07982_));
 sky130_fd_sc_hd__o221ai_1 _27346_ (.A1(_07979_),
    .A2(_07980_),
    .B1(_07981_),
    .B2(_07982_),
    .C1(net2705),
    .Y(_07984_));
 sky130_fd_sc_hd__nor2_1 _27347_ (.A(\inst$top.soc.cpu.gprf.mem[11][6] ),
    .B(net2372),
    .Y(_07985_));
 sky130_fd_sc_hd__o21ai_0 _27348_ (.A1(net2774),
    .A2(\inst$top.soc.cpu.gprf.mem[10][6] ),
    .B1(net2728),
    .Y(_07986_));
 sky130_fd_sc_hd__nor2_1 _27349_ (.A(net2774),
    .B(\inst$top.soc.cpu.gprf.mem[8][6] ),
    .Y(_07987_));
 sky130_fd_sc_hd__o21ai_0 _27350_ (.A1(\inst$top.soc.cpu.gprf.mem[9][6] ),
    .A2(net2372),
    .B1(net2326),
    .Y(_07988_));
 sky130_fd_sc_hd__o221ai_1 _27351_ (.A1(_07985_),
    .A2(_07986_),
    .B1(_07987_),
    .B2(_07988_),
    .C1(net2419),
    .Y(_07989_));
 sky130_fd_sc_hd__nand3_1 _27352_ (.A(_07984_),
    .B(_07989_),
    .C(net2697),
    .Y(_07990_));
 sky130_fd_sc_hd__a32oi_1 _27353_ (.A1(net2694),
    .A2(_07950_),
    .A3(_07963_),
    .B1(_07978_),
    .B2(_07990_),
    .Y(_00060_));
 sky130_fd_sc_hd__nor2_1 _27354_ (.A(\inst$top.soc.cpu.gprf.mem[23][7] ),
    .B(net2393),
    .Y(_07991_));
 sky130_fd_sc_hd__o21ai_0 _27355_ (.A1(net2798),
    .A2(\inst$top.soc.cpu.gprf.mem[22][7] ),
    .B1(net2740),
    .Y(_07992_));
 sky130_fd_sc_hd__nor2_1 _27356_ (.A(net2798),
    .B(\inst$top.soc.cpu.gprf.mem[20][7] ),
    .Y(_07993_));
 sky130_fd_sc_hd__o21ai_0 _27357_ (.A1(\inst$top.soc.cpu.gprf.mem[21][7] ),
    .A2(net2393),
    .B1(net2338),
    .Y(_07994_));
 sky130_fd_sc_hd__o221ai_1 _27358_ (.A1(_07991_),
    .A2(_07992_),
    .B1(_07993_),
    .B2(_07994_),
    .C1(net2711),
    .Y(_07995_));
 sky130_fd_sc_hd__nor2_1 _27359_ (.A(\inst$top.soc.cpu.gprf.mem[19][7] ),
    .B(net2393),
    .Y(_07996_));
 sky130_fd_sc_hd__o21ai_0 _27360_ (.A1(net2798),
    .A2(\inst$top.soc.cpu.gprf.mem[18][7] ),
    .B1(net2740),
    .Y(_07997_));
 sky130_fd_sc_hd__nor2_1 _27361_ (.A(net2798),
    .B(\inst$top.soc.cpu.gprf.mem[16][7] ),
    .Y(_07998_));
 sky130_fd_sc_hd__o21ai_0 _27362_ (.A1(\inst$top.soc.cpu.gprf.mem[17][7] ),
    .A2(net2393),
    .B1(net2336),
    .Y(_07999_));
 sky130_fd_sc_hd__o221ai_1 _27363_ (.A1(_07996_),
    .A2(_07997_),
    .B1(_07998_),
    .B2(_07999_),
    .C1(net2424),
    .Y(_08000_));
 sky130_fd_sc_hd__nand3_1 _27364_ (.A(_07995_),
    .B(_08000_),
    .C(net2438),
    .Y(_08001_));
 sky130_fd_sc_hd__nor2_1 _27365_ (.A(\inst$top.soc.cpu.gprf.mem[31][7] ),
    .B(net2392),
    .Y(_08002_));
 sky130_fd_sc_hd__o21ai_0 _27367_ (.A1(net2799),
    .A2(\inst$top.soc.cpu.gprf.mem[30][7] ),
    .B1(net2740),
    .Y(_08004_));
 sky130_fd_sc_hd__nor2_1 _27368_ (.A(net2797),
    .B(\inst$top.soc.cpu.gprf.mem[28][7] ),
    .Y(_08005_));
 sky130_fd_sc_hd__o21ai_0 _27369_ (.A1(\inst$top.soc.cpu.gprf.mem[29][7] ),
    .A2(net2392),
    .B1(net2336),
    .Y(_08006_));
 sky130_fd_sc_hd__o221ai_1 _27370_ (.A1(_08002_),
    .A2(_08004_),
    .B1(_08005_),
    .B2(_08006_),
    .C1(net2711),
    .Y(_08007_));
 sky130_fd_sc_hd__nor2_1 _27371_ (.A(\inst$top.soc.cpu.gprf.mem[27][7] ),
    .B(net2393),
    .Y(_08008_));
 sky130_fd_sc_hd__o21ai_0 _27372_ (.A1(net2798),
    .A2(\inst$top.soc.cpu.gprf.mem[26][7] ),
    .B1(net2742),
    .Y(_08009_));
 sky130_fd_sc_hd__nor2_1 _27373_ (.A(net2798),
    .B(\inst$top.soc.cpu.gprf.mem[24][7] ),
    .Y(_08010_));
 sky130_fd_sc_hd__o21ai_0 _27374_ (.A1(\inst$top.soc.cpu.gprf.mem[25][7] ),
    .A2(net2393),
    .B1(net2336),
    .Y(_08011_));
 sky130_fd_sc_hd__o221ai_1 _27375_ (.A1(_08008_),
    .A2(_08009_),
    .B1(_08010_),
    .B2(_08011_),
    .C1(net2424),
    .Y(_08012_));
 sky130_fd_sc_hd__nand3_1 _27376_ (.A(_08007_),
    .B(_08012_),
    .C(net2698),
    .Y(_08013_));
 sky130_fd_sc_hd__nor2_1 _27377_ (.A(\inst$top.soc.cpu.gprf.mem[7][7] ),
    .B(net2392),
    .Y(_08014_));
 sky130_fd_sc_hd__o21ai_0 _27378_ (.A1(net2797),
    .A2(\inst$top.soc.cpu.gprf.mem[6][7] ),
    .B1(net2740),
    .Y(_08015_));
 sky130_fd_sc_hd__nor2_1 _27379_ (.A(net2797),
    .B(\inst$top.soc.cpu.gprf.mem[4][7] ),
    .Y(_08016_));
 sky130_fd_sc_hd__o21ai_0 _27380_ (.A1(\inst$top.soc.cpu.gprf.mem[5][7] ),
    .A2(net2392),
    .B1(net2336),
    .Y(_08017_));
 sky130_fd_sc_hd__o221ai_1 _27381_ (.A1(_08014_),
    .A2(_08015_),
    .B1(_08016_),
    .B2(_08017_),
    .C1(net2711),
    .Y(_08018_));
 sky130_fd_sc_hd__nor2_1 _27382_ (.A(\inst$top.soc.cpu.gprf.mem[3][7] ),
    .B(net2392),
    .Y(_08019_));
 sky130_fd_sc_hd__o21ai_0 _27383_ (.A1(net2797),
    .A2(\inst$top.soc.cpu.gprf.mem[2][7] ),
    .B1(net2740),
    .Y(_08020_));
 sky130_fd_sc_hd__nor2_1 _27385_ (.A(net2797),
    .B(\inst$top.soc.cpu.gprf.mem[0][7] ),
    .Y(_08022_));
 sky130_fd_sc_hd__o21ai_0 _27386_ (.A1(\inst$top.soc.cpu.gprf.mem[1][7] ),
    .A2(net2392),
    .B1(net2336),
    .Y(_08023_));
 sky130_fd_sc_hd__o221ai_1 _27387_ (.A1(_08019_),
    .A2(_08020_),
    .B1(_08022_),
    .B2(_08023_),
    .C1(net2424),
    .Y(_08024_));
 sky130_fd_sc_hd__a31oi_1 _27388_ (.A1(_08018_),
    .A2(_08024_),
    .A3(net2438),
    .B1(net2692),
    .Y(_08025_));
 sky130_fd_sc_hd__nor2_1 _27389_ (.A(\inst$top.soc.cpu.gprf.mem[15][7] ),
    .B(net2393),
    .Y(_08026_));
 sky130_fd_sc_hd__o21ai_0 _27390_ (.A1(net2798),
    .A2(\inst$top.soc.cpu.gprf.mem[14][7] ),
    .B1(net2740),
    .Y(_08027_));
 sky130_fd_sc_hd__nor2_1 _27391_ (.A(net2798),
    .B(\inst$top.soc.cpu.gprf.mem[12][7] ),
    .Y(_08028_));
 sky130_fd_sc_hd__o21ai_0 _27392_ (.A1(\inst$top.soc.cpu.gprf.mem[13][7] ),
    .A2(net2393),
    .B1(net2338),
    .Y(_08029_));
 sky130_fd_sc_hd__o22ai_1 _27393_ (.A1(_08026_),
    .A2(_08027_),
    .B1(_08028_),
    .B2(_08029_),
    .Y(_08030_));
 sky130_fd_sc_hd__nor2_1 _27395_ (.A(\inst$top.soc.cpu.gprf.mem[11][7] ),
    .B(net2393),
    .Y(_08032_));
 sky130_fd_sc_hd__o21ai_0 _27396_ (.A1(net2798),
    .A2(\inst$top.soc.cpu.gprf.mem[10][7] ),
    .B1(net2742),
    .Y(_08033_));
 sky130_fd_sc_hd__nor2_1 _27397_ (.A(net2798),
    .B(\inst$top.soc.cpu.gprf.mem[8][7] ),
    .Y(_08034_));
 sky130_fd_sc_hd__o21ai_0 _27398_ (.A1(\inst$top.soc.cpu.gprf.mem[9][7] ),
    .A2(net2393),
    .B1(net2338),
    .Y(_08035_));
 sky130_fd_sc_hd__o22ai_1 _27399_ (.A1(_08032_),
    .A2(_08033_),
    .B1(_08034_),
    .B2(_08035_),
    .Y(_08036_));
 sky130_fd_sc_hd__nor2_1 _27400_ (.A(net2711),
    .B(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__nor2_1 _27401_ (.A(net2438),
    .B(_08037_),
    .Y(_08038_));
 sky130_fd_sc_hd__o21ai_0 _27402_ (.A1(net2424),
    .A2(_08030_),
    .B1(_08038_),
    .Y(_08039_));
 sky130_fd_sc_hd__a32oi_1 _27403_ (.A1(_08001_),
    .A2(_08013_),
    .A3(net2691),
    .B1(_08025_),
    .B2(_08039_),
    .Y(_00061_));
 sky130_fd_sc_hd__nor2_1 _27404_ (.A(\inst$top.soc.cpu.gprf.mem[7][8] ),
    .B(net2359),
    .Y(_08040_));
 sky130_fd_sc_hd__o21ai_0 _27405_ (.A1(net2771),
    .A2(\inst$top.soc.cpu.gprf.mem[6][8] ),
    .B1(net2726),
    .Y(_08041_));
 sky130_fd_sc_hd__nor2_1 _27406_ (.A(net2771),
    .B(\inst$top.soc.cpu.gprf.mem[4][8] ),
    .Y(_08042_));
 sky130_fd_sc_hd__o21ai_0 _27407_ (.A1(\inst$top.soc.cpu.gprf.mem[5][8] ),
    .A2(net2359),
    .B1(net2317),
    .Y(_08043_));
 sky130_fd_sc_hd__o221ai_1 _27408_ (.A1(_08040_),
    .A2(_08041_),
    .B1(_08042_),
    .B2(_08043_),
    .C1(net2704),
    .Y(_08044_));
 sky130_fd_sc_hd__nor2_1 _27409_ (.A(\inst$top.soc.cpu.gprf.mem[3][8] ),
    .B(net2368),
    .Y(_08045_));
 sky130_fd_sc_hd__o21ai_0 _27410_ (.A1(net2771),
    .A2(\inst$top.soc.cpu.gprf.mem[2][8] ),
    .B1(net2726),
    .Y(_08046_));
 sky130_fd_sc_hd__nor2_1 _27411_ (.A(net2771),
    .B(\inst$top.soc.cpu.gprf.mem[0][8] ),
    .Y(_08047_));
 sky130_fd_sc_hd__o21ai_0 _27412_ (.A1(\inst$top.soc.cpu.gprf.mem[1][8] ),
    .A2(net2368),
    .B1(net2324),
    .Y(_08048_));
 sky130_fd_sc_hd__o221ai_1 _27413_ (.A1(_08045_),
    .A2(_08046_),
    .B1(_08047_),
    .B2(_08048_),
    .C1(net2418),
    .Y(_08049_));
 sky130_fd_sc_hd__nand3_1 _27414_ (.A(_08044_),
    .B(_08049_),
    .C(net2433),
    .Y(_08050_));
 sky130_fd_sc_hd__nor2_1 _27415_ (.A(\inst$top.soc.cpu.gprf.mem[11][8] ),
    .B(net2365),
    .Y(_08051_));
 sky130_fd_sc_hd__o21ai_0 _27416_ (.A1(net2770),
    .A2(\inst$top.soc.cpu.gprf.mem[10][8] ),
    .B1(net2725),
    .Y(_08052_));
 sky130_fd_sc_hd__nor2_1 _27417_ (.A(net2768),
    .B(\inst$top.soc.cpu.gprf.mem[8][8] ),
    .Y(_08053_));
 sky130_fd_sc_hd__o21ai_0 _27418_ (.A1(\inst$top.soc.cpu.gprf.mem[9][8] ),
    .A2(net2365),
    .B1(net2323),
    .Y(_08054_));
 sky130_fd_sc_hd__o221ai_1 _27419_ (.A1(_08051_),
    .A2(_08052_),
    .B1(_08053_),
    .B2(_08054_),
    .C1(net2418),
    .Y(_08055_));
 sky130_fd_sc_hd__nor2_1 _27421_ (.A(\inst$top.soc.cpu.gprf.mem[15][8] ),
    .B(net2357),
    .Y(_08057_));
 sky130_fd_sc_hd__o21ai_0 _27423_ (.A1(net2770),
    .A2(\inst$top.soc.cpu.gprf.mem[14][8] ),
    .B1(net2725),
    .Y(_08059_));
 sky130_fd_sc_hd__nor2_1 _27424_ (.A(net2768),
    .B(\inst$top.soc.cpu.gprf.mem[12][8] ),
    .Y(_08060_));
 sky130_fd_sc_hd__o21ai_0 _27425_ (.A1(\inst$top.soc.cpu.gprf.mem[13][8] ),
    .A2(net2356),
    .B1(net2316),
    .Y(_08061_));
 sky130_fd_sc_hd__o221ai_1 _27426_ (.A1(_08057_),
    .A2(_08059_),
    .B1(_08060_),
    .B2(_08061_),
    .C1(net2704),
    .Y(_08062_));
 sky130_fd_sc_hd__nand3_1 _27427_ (.A(_08055_),
    .B(_08062_),
    .C(net2697),
    .Y(_08063_));
 sky130_fd_sc_hd__nor2_1 _27428_ (.A(\inst$top.soc.cpu.gprf.mem[31][8] ),
    .B(net2359),
    .Y(_08064_));
 sky130_fd_sc_hd__o21ai_0 _27429_ (.A1(net2771),
    .A2(\inst$top.soc.cpu.gprf.mem[30][8] ),
    .B1(net2726),
    .Y(_08065_));
 sky130_fd_sc_hd__nor2_1 _27430_ (.A(net2761),
    .B(\inst$top.soc.cpu.gprf.mem[28][8] ),
    .Y(_08066_));
 sky130_fd_sc_hd__o21ai_0 _27431_ (.A1(\inst$top.soc.cpu.gprf.mem[29][8] ),
    .A2(net2359),
    .B1(net2317),
    .Y(_08067_));
 sky130_fd_sc_hd__o221ai_1 _27432_ (.A1(_08064_),
    .A2(_08065_),
    .B1(_08066_),
    .B2(_08067_),
    .C1(net2701),
    .Y(_08068_));
 sky130_fd_sc_hd__nor2_1 _27433_ (.A(\inst$top.soc.cpu.gprf.mem[27][8] ),
    .B(net2359),
    .Y(_08069_));
 sky130_fd_sc_hd__o21ai_0 _27434_ (.A1(net2771),
    .A2(\inst$top.soc.cpu.gprf.mem[26][8] ),
    .B1(net2726),
    .Y(_08070_));
 sky130_fd_sc_hd__nor2_1 _27435_ (.A(net2773),
    .B(\inst$top.soc.cpu.gprf.mem[24][8] ),
    .Y(_08071_));
 sky130_fd_sc_hd__o21ai_0 _27437_ (.A1(\inst$top.soc.cpu.gprf.mem[25][8] ),
    .A2(net2368),
    .B1(net2324),
    .Y(_08073_));
 sky130_fd_sc_hd__o221ai_1 _27439_ (.A1(_08069_),
    .A2(_08070_),
    .B1(_08071_),
    .B2(_08073_),
    .C1(net2420),
    .Y(_08075_));
 sky130_fd_sc_hd__a31oi_1 _27441_ (.A1(_08068_),
    .A2(_08075_),
    .A3(net2697),
    .B1(net2442),
    .Y(_08077_));
 sky130_fd_sc_hd__nor2_1 _27442_ (.A(\inst$top.soc.cpu.gprf.mem[23][8] ),
    .B(net2368),
    .Y(_08078_));
 sky130_fd_sc_hd__o21ai_0 _27444_ (.A1(net2773),
    .A2(\inst$top.soc.cpu.gprf.mem[22][8] ),
    .B1(net2726),
    .Y(_08080_));
 sky130_fd_sc_hd__nor2_1 _27445_ (.A(net2771),
    .B(\inst$top.soc.cpu.gprf.mem[20][8] ),
    .Y(_08081_));
 sky130_fd_sc_hd__o21ai_0 _27447_ (.A1(\inst$top.soc.cpu.gprf.mem[21][8] ),
    .A2(net2368),
    .B1(net2324),
    .Y(_08083_));
 sky130_fd_sc_hd__o221ai_1 _27448_ (.A1(_08078_),
    .A2(_08080_),
    .B1(_08081_),
    .B2(_08083_),
    .C1(net2706),
    .Y(_08084_));
 sky130_fd_sc_hd__nor2_1 _27449_ (.A(\inst$top.soc.cpu.gprf.mem[19][8] ),
    .B(net2368),
    .Y(_08085_));
 sky130_fd_sc_hd__o21ai_0 _27450_ (.A1(net2771),
    .A2(\inst$top.soc.cpu.gprf.mem[18][8] ),
    .B1(net2726),
    .Y(_08086_));
 sky130_fd_sc_hd__nor2_1 _27451_ (.A(net2771),
    .B(\inst$top.soc.cpu.gprf.mem[16][8] ),
    .Y(_08087_));
 sky130_fd_sc_hd__o21ai_0 _27453_ (.A1(\inst$top.soc.cpu.gprf.mem[17][8] ),
    .A2(net2368),
    .B1(net2324),
    .Y(_08089_));
 sky130_fd_sc_hd__o221ai_1 _27454_ (.A1(_08085_),
    .A2(_08086_),
    .B1(_08087_),
    .B2(_08089_),
    .C1(net2418),
    .Y(_08090_));
 sky130_fd_sc_hd__nand3_1 _27456_ (.A(_08084_),
    .B(_08090_),
    .C(net2433),
    .Y(_08092_));
 sky130_fd_sc_hd__a32oi_1 _27457_ (.A1(_08050_),
    .A2(_08063_),
    .A3(net2442),
    .B1(_08077_),
    .B2(_08092_),
    .Y(_00062_));
 sky130_fd_sc_hd__nor2_1 _27458_ (.A(\inst$top.soc.cpu.gprf.mem[31][9] ),
    .B(net2373),
    .Y(_08093_));
 sky130_fd_sc_hd__o21ai_0 _27459_ (.A1(net2779),
    .A2(\inst$top.soc.cpu.gprf.mem[30][9] ),
    .B1(net2730),
    .Y(_08094_));
 sky130_fd_sc_hd__nor2_1 _27461_ (.A(net2779),
    .B(\inst$top.soc.cpu.gprf.mem[28][9] ),
    .Y(_08096_));
 sky130_fd_sc_hd__o21ai_0 _27462_ (.A1(\inst$top.soc.cpu.gprf.mem[29][9] ),
    .A2(net2373),
    .B1(net2327),
    .Y(_08097_));
 sky130_fd_sc_hd__o22ai_1 _27463_ (.A1(_08093_),
    .A2(_08094_),
    .B1(_08096_),
    .B2(_08097_),
    .Y(_08098_));
 sky130_fd_sc_hd__nor2_1 _27464_ (.A(\inst$top.soc.cpu.gprf.mem[27][9] ),
    .B(net2373),
    .Y(_08099_));
 sky130_fd_sc_hd__o21ai_0 _27465_ (.A1(net2778),
    .A2(\inst$top.soc.cpu.gprf.mem[26][9] ),
    .B1(net2729),
    .Y(_08100_));
 sky130_fd_sc_hd__nor2_1 _27466_ (.A(net2778),
    .B(\inst$top.soc.cpu.gprf.mem[24][9] ),
    .Y(_08101_));
 sky130_fd_sc_hd__o21ai_0 _27468_ (.A1(\inst$top.soc.cpu.gprf.mem[25][9] ),
    .A2(net2374),
    .B1(net2327),
    .Y(_08103_));
 sky130_fd_sc_hd__o22ai_1 _27469_ (.A1(_08099_),
    .A2(_08100_),
    .B1(_08101_),
    .B2(_08103_),
    .Y(_08104_));
 sky130_fd_sc_hd__nor2_1 _27470_ (.A(net2706),
    .B(_08104_),
    .Y(_08105_));
 sky130_fd_sc_hd__nor2_1 _27471_ (.A(net2433),
    .B(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__o21ai_0 _27472_ (.A1(net2419),
    .A2(_08098_),
    .B1(_08106_),
    .Y(_08107_));
 sky130_fd_sc_hd__nor2_1 _27473_ (.A(\inst$top.soc.cpu.gprf.mem[23][9] ),
    .B(net2374),
    .Y(_08108_));
 sky130_fd_sc_hd__o21ai_0 _27474_ (.A1(net2778),
    .A2(\inst$top.soc.cpu.gprf.mem[22][9] ),
    .B1(net2729),
    .Y(_08109_));
 sky130_fd_sc_hd__nor2_1 _27475_ (.A(net2778),
    .B(\inst$top.soc.cpu.gprf.mem[20][9] ),
    .Y(_08110_));
 sky130_fd_sc_hd__o21ai_0 _27476_ (.A1(\inst$top.soc.cpu.gprf.mem[21][9] ),
    .A2(net2374),
    .B1(net2327),
    .Y(_08111_));
 sky130_fd_sc_hd__o221ai_1 _27477_ (.A1(_08108_),
    .A2(_08109_),
    .B1(_08110_),
    .B2(_08111_),
    .C1(net2706),
    .Y(_08112_));
 sky130_fd_sc_hd__nor2_1 _27478_ (.A(\inst$top.soc.cpu.gprf.mem[19][9] ),
    .B(net2382),
    .Y(_08113_));
 sky130_fd_sc_hd__o21ai_0 _27479_ (.A1(net2778),
    .A2(\inst$top.soc.cpu.gprf.mem[18][9] ),
    .B1(net2735),
    .Y(_08114_));
 sky130_fd_sc_hd__nor2_1 _27480_ (.A(net2785),
    .B(\inst$top.soc.cpu.gprf.mem[16][9] ),
    .Y(_08115_));
 sky130_fd_sc_hd__o21ai_0 _27482_ (.A1(\inst$top.soc.cpu.gprf.mem[17][9] ),
    .A2(net2382),
    .B1(net2332),
    .Y(_08117_));
 sky130_fd_sc_hd__o221ai_1 _27483_ (.A1(_08113_),
    .A2(_08114_),
    .B1(_08115_),
    .B2(_08117_),
    .C1(net2419),
    .Y(_08118_));
 sky130_fd_sc_hd__nand3_1 _27484_ (.A(_08112_),
    .B(_08118_),
    .C(net2434),
    .Y(_08119_));
 sky130_fd_sc_hd__nor2_1 _27485_ (.A(\inst$top.soc.cpu.gprf.mem[11][9] ),
    .B(net2375),
    .Y(_08120_));
 sky130_fd_sc_hd__o21ai_0 _27486_ (.A1(net2778),
    .A2(\inst$top.soc.cpu.gprf.mem[10][9] ),
    .B1(net2730),
    .Y(_08121_));
 sky130_fd_sc_hd__nor2_1 _27487_ (.A(net2779),
    .B(\inst$top.soc.cpu.gprf.mem[8][9] ),
    .Y(_08122_));
 sky130_fd_sc_hd__o21ai_0 _27489_ (.A1(\inst$top.soc.cpu.gprf.mem[9][9] ),
    .A2(net2374),
    .B1(net2328),
    .Y(_08124_));
 sky130_fd_sc_hd__o221ai_1 _27491_ (.A1(_08120_),
    .A2(_08121_),
    .B1(_08122_),
    .B2(_08124_),
    .C1(net2420),
    .Y(_08126_));
 sky130_fd_sc_hd__nor2_1 _27492_ (.A(\inst$top.soc.cpu.gprf.mem[15][9] ),
    .B(net2374),
    .Y(_08127_));
 sky130_fd_sc_hd__o21ai_0 _27494_ (.A1(net2796),
    .A2(\inst$top.soc.cpu.gprf.mem[14][9] ),
    .B1(net2738),
    .Y(_08129_));
 sky130_fd_sc_hd__nor2_1 _27495_ (.A(net2796),
    .B(\inst$top.soc.cpu.gprf.mem[12][9] ),
    .Y(_08130_));
 sky130_fd_sc_hd__o21ai_0 _27496_ (.A1(\inst$top.soc.cpu.gprf.mem[13][9] ),
    .A2(net2374),
    .B1(net2327),
    .Y(_08131_));
 sky130_fd_sc_hd__o221ai_1 _27497_ (.A1(_08127_),
    .A2(_08129_),
    .B1(_08130_),
    .B2(_08131_),
    .C1(net2705),
    .Y(_08132_));
 sky130_fd_sc_hd__a31oi_1 _27498_ (.A1(_08126_),
    .A2(_08132_),
    .A3(net2699),
    .B1(net2691),
    .Y(_08133_));
 sky130_fd_sc_hd__nor2_1 _27499_ (.A(\inst$top.soc.cpu.gprf.mem[7][9] ),
    .B(net2373),
    .Y(_08134_));
 sky130_fd_sc_hd__o21ai_0 _27500_ (.A1(net2779),
    .A2(\inst$top.soc.cpu.gprf.mem[6][9] ),
    .B1(net2729),
    .Y(_08135_));
 sky130_fd_sc_hd__nor2_1 _27501_ (.A(net2777),
    .B(\inst$top.soc.cpu.gprf.mem[4][9] ),
    .Y(_08136_));
 sky130_fd_sc_hd__o21ai_0 _27502_ (.A1(\inst$top.soc.cpu.gprf.mem[5][9] ),
    .A2(net2375),
    .B1(net2327),
    .Y(_08137_));
 sky130_fd_sc_hd__o221ai_1 _27503_ (.A1(_08134_),
    .A2(_08135_),
    .B1(_08136_),
    .B2(_08137_),
    .C1(net2706),
    .Y(_08138_));
 sky130_fd_sc_hd__nor2_1 _27504_ (.A(\inst$top.soc.cpu.gprf.mem[3][9] ),
    .B(net2373),
    .Y(_08139_));
 sky130_fd_sc_hd__o21ai_0 _27505_ (.A1(net2777),
    .A2(\inst$top.soc.cpu.gprf.mem[2][9] ),
    .B1(net2729),
    .Y(_08140_));
 sky130_fd_sc_hd__nor2_1 _27507_ (.A(net2779),
    .B(\inst$top.soc.cpu.gprf.mem[0][9] ),
    .Y(_08142_));
 sky130_fd_sc_hd__o21ai_0 _27508_ (.A1(\inst$top.soc.cpu.gprf.mem[1][9] ),
    .A2(net2373),
    .B1(net2327),
    .Y(_08143_));
 sky130_fd_sc_hd__o221ai_1 _27511_ (.A1(_08139_),
    .A2(_08140_),
    .B1(_08142_),
    .B2(_08143_),
    .C1(net2420),
    .Y(_08146_));
 sky130_fd_sc_hd__nand3_1 _27512_ (.A(_08138_),
    .B(_08146_),
    .C(net2434),
    .Y(_08147_));
 sky130_fd_sc_hd__a32oi_1 _27513_ (.A1(net2694),
    .A2(_08107_),
    .A3(_08119_),
    .B1(_08133_),
    .B2(_08147_),
    .Y(_00063_));
 sky130_fd_sc_hd__nor2_1 _27514_ (.A(\inst$top.soc.cpu.gprf.mem[11][10] ),
    .B(net2382),
    .Y(_08148_));
 sky130_fd_sc_hd__o21ai_0 _27515_ (.A1(net2785),
    .A2(\inst$top.soc.cpu.gprf.mem[10][10] ),
    .B1(net2735),
    .Y(_08149_));
 sky130_fd_sc_hd__nor2_1 _27516_ (.A(net2786),
    .B(\inst$top.soc.cpu.gprf.mem[8][10] ),
    .Y(_08150_));
 sky130_fd_sc_hd__o21ai_0 _27517_ (.A1(\inst$top.soc.cpu.gprf.mem[9][10] ),
    .A2(net2382),
    .B1(net2332),
    .Y(_08151_));
 sky130_fd_sc_hd__o22ai_1 _27518_ (.A1(_08148_),
    .A2(_08149_),
    .B1(_08150_),
    .B2(_08151_),
    .Y(_08152_));
 sky130_fd_sc_hd__nor2_1 _27520_ (.A(\inst$top.soc.cpu.gprf.mem[15][10] ),
    .B(net2382),
    .Y(_08154_));
 sky130_fd_sc_hd__o21ai_0 _27521_ (.A1(net2785),
    .A2(\inst$top.soc.cpu.gprf.mem[14][10] ),
    .B1(net2735),
    .Y(_08155_));
 sky130_fd_sc_hd__nor2_1 _27522_ (.A(net2785),
    .B(\inst$top.soc.cpu.gprf.mem[12][10] ),
    .Y(_08156_));
 sky130_fd_sc_hd__o21ai_0 _27523_ (.A1(\inst$top.soc.cpu.gprf.mem[13][10] ),
    .A2(net2382),
    .B1(net2332),
    .Y(_08157_));
 sky130_fd_sc_hd__o22ai_1 _27524_ (.A1(_08154_),
    .A2(_08155_),
    .B1(_08156_),
    .B2(_08157_),
    .Y(_08158_));
 sky130_fd_sc_hd__nor2_1 _27525_ (.A(net2422),
    .B(_08158_),
    .Y(_08159_));
 sky130_fd_sc_hd__nor2_1 _27526_ (.A(net2436),
    .B(_08159_),
    .Y(_08160_));
 sky130_fd_sc_hd__o21ai_0 _27527_ (.A1(net2708),
    .A2(_08152_),
    .B1(_08160_),
    .Y(_08161_));
 sky130_fd_sc_hd__nor2_1 _27528_ (.A(\inst$top.soc.cpu.gprf.mem[7][10] ),
    .B(net2380),
    .Y(_08162_));
 sky130_fd_sc_hd__o21ai_0 _27529_ (.A1(net2781),
    .A2(\inst$top.soc.cpu.gprf.mem[6][10] ),
    .B1(net2733),
    .Y(_08163_));
 sky130_fd_sc_hd__nor2_1 _27530_ (.A(net2785),
    .B(\inst$top.soc.cpu.gprf.mem[4][10] ),
    .Y(_08164_));
 sky130_fd_sc_hd__o21ai_0 _27531_ (.A1(\inst$top.soc.cpu.gprf.mem[5][10] ),
    .A2(net2376),
    .B1(net2329),
    .Y(_08165_));
 sky130_fd_sc_hd__o221ai_1 _27532_ (.A1(_08162_),
    .A2(_08163_),
    .B1(_08164_),
    .B2(_08165_),
    .C1(net2707),
    .Y(_08166_));
 sky130_fd_sc_hd__nor2_1 _27533_ (.A(\inst$top.soc.cpu.gprf.mem[3][10] ),
    .B(net2376),
    .Y(_08167_));
 sky130_fd_sc_hd__o21ai_0 _27534_ (.A1(net2785),
    .A2(\inst$top.soc.cpu.gprf.mem[2][10] ),
    .B1(net2735),
    .Y(_08168_));
 sky130_fd_sc_hd__nor2_1 _27535_ (.A(net2785),
    .B(\inst$top.soc.cpu.gprf.mem[0][10] ),
    .Y(_08169_));
 sky130_fd_sc_hd__o21ai_0 _27536_ (.A1(\inst$top.soc.cpu.gprf.mem[1][10] ),
    .A2(net2376),
    .B1(net2332),
    .Y(_08170_));
 sky130_fd_sc_hd__o221ai_1 _27537_ (.A1(_08167_),
    .A2(_08168_),
    .B1(_08169_),
    .B2(_08170_),
    .C1(net2421),
    .Y(_08171_));
 sky130_fd_sc_hd__nand3_1 _27538_ (.A(_08166_),
    .B(_08171_),
    .C(net2435),
    .Y(_08172_));
 sky130_fd_sc_hd__nor2_1 _27539_ (.A(\inst$top.soc.cpu.gprf.mem[31][10] ),
    .B(net2376),
    .Y(_08173_));
 sky130_fd_sc_hd__o21ai_0 _27540_ (.A1(net2781),
    .A2(\inst$top.soc.cpu.gprf.mem[30][10] ),
    .B1(net2733),
    .Y(_08174_));
 sky130_fd_sc_hd__nor2_1 _27541_ (.A(net2781),
    .B(\inst$top.soc.cpu.gprf.mem[28][10] ),
    .Y(_08175_));
 sky130_fd_sc_hd__o21ai_0 _27542_ (.A1(\inst$top.soc.cpu.gprf.mem[29][10] ),
    .A2(net2376),
    .B1(net2329),
    .Y(_08176_));
 sky130_fd_sc_hd__o221ai_1 _27543_ (.A1(_08173_),
    .A2(_08174_),
    .B1(_08175_),
    .B2(_08176_),
    .C1(net2707),
    .Y(_08177_));
 sky130_fd_sc_hd__nor2_1 _27544_ (.A(\inst$top.soc.cpu.gprf.mem[27][10] ),
    .B(net2376),
    .Y(_08178_));
 sky130_fd_sc_hd__o21ai_0 _27545_ (.A1(net2785),
    .A2(\inst$top.soc.cpu.gprf.mem[26][10] ),
    .B1(net2735),
    .Y(_08179_));
 sky130_fd_sc_hd__nor2_1 _27546_ (.A(net2785),
    .B(\inst$top.soc.cpu.gprf.mem[24][10] ),
    .Y(_08180_));
 sky130_fd_sc_hd__o21ai_0 _27547_ (.A1(\inst$top.soc.cpu.gprf.mem[25][10] ),
    .A2(net2376),
    .B1(net2332),
    .Y(_08181_));
 sky130_fd_sc_hd__o221ai_1 _27548_ (.A1(_08178_),
    .A2(_08179_),
    .B1(_08180_),
    .B2(_08181_),
    .C1(net2422),
    .Y(_08182_));
 sky130_fd_sc_hd__a31oi_1 _27549_ (.A1(_08177_),
    .A2(_08182_),
    .A3(net2699),
    .B1(net2442),
    .Y(_08183_));
 sky130_fd_sc_hd__nor2_1 _27550_ (.A(\inst$top.soc.cpu.gprf.mem[23][10] ),
    .B(net2376),
    .Y(_08184_));
 sky130_fd_sc_hd__o21ai_0 _27551_ (.A1(net2784),
    .A2(\inst$top.soc.cpu.gprf.mem[22][10] ),
    .B1(net2731),
    .Y(_08185_));
 sky130_fd_sc_hd__nor2_1 _27552_ (.A(net2781),
    .B(\inst$top.soc.cpu.gprf.mem[20][10] ),
    .Y(_08186_));
 sky130_fd_sc_hd__o21ai_0 _27553_ (.A1(\inst$top.soc.cpu.gprf.mem[21][10] ),
    .A2(net2376),
    .B1(net2329),
    .Y(_08187_));
 sky130_fd_sc_hd__o221ai_1 _27554_ (.A1(_08184_),
    .A2(_08185_),
    .B1(_08186_),
    .B2(_08187_),
    .C1(net2707),
    .Y(_08188_));
 sky130_fd_sc_hd__nor2_1 _27556_ (.A(\inst$top.soc.cpu.gprf.mem[19][10] ),
    .B(net2380),
    .Y(_08190_));
 sky130_fd_sc_hd__o21ai_0 _27557_ (.A1(net2781),
    .A2(\inst$top.soc.cpu.gprf.mem[18][10] ),
    .B1(net2731),
    .Y(_08191_));
 sky130_fd_sc_hd__nor2_1 _27558_ (.A(net2784),
    .B(\inst$top.soc.cpu.gprf.mem[16][10] ),
    .Y(_08192_));
 sky130_fd_sc_hd__o21ai_0 _27559_ (.A1(\inst$top.soc.cpu.gprf.mem[17][10] ),
    .A2(net2377),
    .B1(net2329),
    .Y(_08193_));
 sky130_fd_sc_hd__o221ai_1 _27560_ (.A1(_08190_),
    .A2(_08191_),
    .B1(_08192_),
    .B2(_08193_),
    .C1(net2421),
    .Y(_08194_));
 sky130_fd_sc_hd__nand3_1 _27561_ (.A(_08188_),
    .B(_08194_),
    .C(net2435),
    .Y(_08195_));
 sky130_fd_sc_hd__a32oi_1 _27562_ (.A1(net2442),
    .A2(_08161_),
    .A3(_08172_),
    .B1(_08183_),
    .B2(_08195_),
    .Y(_00033_));
 sky130_fd_sc_hd__nor2_1 _27563_ (.A(\inst$top.soc.cpu.gprf.mem[23][11] ),
    .B(net2363),
    .Y(_08196_));
 sky130_fd_sc_hd__o21ai_0 _27564_ (.A1(net2766),
    .A2(\inst$top.soc.cpu.gprf.mem[22][11] ),
    .B1(net2723),
    .Y(_08197_));
 sky130_fd_sc_hd__nor2_1 _27565_ (.A(net2766),
    .B(\inst$top.soc.cpu.gprf.mem[20][11] ),
    .Y(_08198_));
 sky130_fd_sc_hd__o21ai_0 _27566_ (.A1(\inst$top.soc.cpu.gprf.mem[21][11] ),
    .A2(net2363),
    .B1(net2320),
    .Y(_08199_));
 sky130_fd_sc_hd__o221ai_1 _27567_ (.A1(_08196_),
    .A2(_08197_),
    .B1(_08198_),
    .B2(_08199_),
    .C1(net2703),
    .Y(_08200_));
 sky130_fd_sc_hd__nor2_1 _27568_ (.A(\inst$top.soc.cpu.gprf.mem[19][11] ),
    .B(net2363),
    .Y(_08201_));
 sky130_fd_sc_hd__o21ai_0 _27569_ (.A1(net2783),
    .A2(\inst$top.soc.cpu.gprf.mem[18][11] ),
    .B1(net2732),
    .Y(_08202_));
 sky130_fd_sc_hd__nor2_1 _27570_ (.A(net2783),
    .B(\inst$top.soc.cpu.gprf.mem[16][11] ),
    .Y(_08203_));
 sky130_fd_sc_hd__o21ai_0 _27571_ (.A1(\inst$top.soc.cpu.gprf.mem[17][11] ),
    .A2(net2363),
    .B1(net2320),
    .Y(_08204_));
 sky130_fd_sc_hd__o221ai_1 _27572_ (.A1(_08201_),
    .A2(_08202_),
    .B1(_08203_),
    .B2(_08204_),
    .C1(net2415),
    .Y(_08205_));
 sky130_fd_sc_hd__nand3_1 _27573_ (.A(_08200_),
    .B(_08205_),
    .C(net2431),
    .Y(_08206_));
 sky130_fd_sc_hd__nor2_1 _27574_ (.A(\inst$top.soc.cpu.gprf.mem[31][11] ),
    .B(net2377),
    .Y(_08207_));
 sky130_fd_sc_hd__o21ai_0 _27575_ (.A1(net2781),
    .A2(\inst$top.soc.cpu.gprf.mem[30][11] ),
    .B1(net2731),
    .Y(_08208_));
 sky130_fd_sc_hd__nor2_1 _27576_ (.A(net2780),
    .B(\inst$top.soc.cpu.gprf.mem[28][11] ),
    .Y(_08209_));
 sky130_fd_sc_hd__o21ai_0 _27577_ (.A1(\inst$top.soc.cpu.gprf.mem[29][11] ),
    .A2(net2377),
    .B1(net2329),
    .Y(_08210_));
 sky130_fd_sc_hd__o221ai_1 _27578_ (.A1(_08207_),
    .A2(_08208_),
    .B1(_08209_),
    .B2(_08210_),
    .C1(net2707),
    .Y(_08211_));
 sky130_fd_sc_hd__nor2_1 _27579_ (.A(\inst$top.soc.cpu.gprf.mem[27][11] ),
    .B(net2363),
    .Y(_08212_));
 sky130_fd_sc_hd__o21ai_0 _27580_ (.A1(net2781),
    .A2(\inst$top.soc.cpu.gprf.mem[26][11] ),
    .B1(net2731),
    .Y(_08213_));
 sky130_fd_sc_hd__nor2_1 _27581_ (.A(net2764),
    .B(\inst$top.soc.cpu.gprf.mem[24][11] ),
    .Y(_08214_));
 sky130_fd_sc_hd__o21ai_0 _27582_ (.A1(\inst$top.soc.cpu.gprf.mem[25][11] ),
    .A2(net2361),
    .B1(net2319),
    .Y(_08215_));
 sky130_fd_sc_hd__o221ai_1 _27583_ (.A1(_08212_),
    .A2(_08213_),
    .B1(_08214_),
    .B2(_08215_),
    .C1(net2415),
    .Y(_08216_));
 sky130_fd_sc_hd__nand3_1 _27584_ (.A(_08211_),
    .B(_08216_),
    .C(net2697),
    .Y(_08217_));
 sky130_fd_sc_hd__nor2_1 _27585_ (.A(\inst$top.soc.cpu.gprf.mem[7][11] ),
    .B(net2364),
    .Y(_08218_));
 sky130_fd_sc_hd__o21ai_0 _27586_ (.A1(net2783),
    .A2(\inst$top.soc.cpu.gprf.mem[6][11] ),
    .B1(net2732),
    .Y(_08219_));
 sky130_fd_sc_hd__nor2_1 _27587_ (.A(net2783),
    .B(\inst$top.soc.cpu.gprf.mem[4][11] ),
    .Y(_08220_));
 sky130_fd_sc_hd__o21ai_0 _27588_ (.A1(\inst$top.soc.cpu.gprf.mem[5][11] ),
    .A2(net2364),
    .B1(net2320),
    .Y(_08221_));
 sky130_fd_sc_hd__o221ai_1 _27589_ (.A1(_08218_),
    .A2(_08219_),
    .B1(_08220_),
    .B2(_08221_),
    .C1(net2707),
    .Y(_08222_));
 sky130_fd_sc_hd__nor2_1 _27590_ (.A(\inst$top.soc.cpu.gprf.mem[3][11] ),
    .B(net2363),
    .Y(_08223_));
 sky130_fd_sc_hd__o21ai_0 _27591_ (.A1(net2766),
    .A2(\inst$top.soc.cpu.gprf.mem[2][11] ),
    .B1(net2723),
    .Y(_08224_));
 sky130_fd_sc_hd__nor2_1 _27592_ (.A(net2766),
    .B(\inst$top.soc.cpu.gprf.mem[0][11] ),
    .Y(_08225_));
 sky130_fd_sc_hd__o21ai_0 _27593_ (.A1(\inst$top.soc.cpu.gprf.mem[1][11] ),
    .A2(net2363),
    .B1(net2320),
    .Y(_08226_));
 sky130_fd_sc_hd__o221ai_1 _27594_ (.A1(_08223_),
    .A2(_08224_),
    .B1(_08225_),
    .B2(_08226_),
    .C1(net2415),
    .Y(_08227_));
 sky130_fd_sc_hd__a31oi_1 _27595_ (.A1(_08222_),
    .A2(_08227_),
    .A3(net2431),
    .B1(net2694),
    .Y(_08228_));
 sky130_fd_sc_hd__nor2_1 _27596_ (.A(\inst$top.soc.cpu.gprf.mem[15][11] ),
    .B(net2361),
    .Y(_08229_));
 sky130_fd_sc_hd__o21ai_0 _27597_ (.A1(net2780),
    .A2(\inst$top.soc.cpu.gprf.mem[14][11] ),
    .B1(net2731),
    .Y(_08230_));
 sky130_fd_sc_hd__nor2_1 _27598_ (.A(net2780),
    .B(\inst$top.soc.cpu.gprf.mem[12][11] ),
    .Y(_08231_));
 sky130_fd_sc_hd__o21ai_0 _27599_ (.A1(\inst$top.soc.cpu.gprf.mem[13][11] ),
    .A2(net2361),
    .B1(net2319),
    .Y(_08232_));
 sky130_fd_sc_hd__o22ai_1 _27600_ (.A1(_08229_),
    .A2(_08230_),
    .B1(_08231_),
    .B2(_08232_),
    .Y(_08233_));
 sky130_fd_sc_hd__nor2_1 _27601_ (.A(\inst$top.soc.cpu.gprf.mem[11][11] ),
    .B(net2377),
    .Y(_08234_));
 sky130_fd_sc_hd__o21ai_0 _27602_ (.A1(net2780),
    .A2(\inst$top.soc.cpu.gprf.mem[10][11] ),
    .B1(net2731),
    .Y(_08235_));
 sky130_fd_sc_hd__nor2_1 _27603_ (.A(net2780),
    .B(\inst$top.soc.cpu.gprf.mem[8][11] ),
    .Y(_08236_));
 sky130_fd_sc_hd__o21ai_0 _27604_ (.A1(\inst$top.soc.cpu.gprf.mem[9][11] ),
    .A2(net2377),
    .B1(net2329),
    .Y(_08237_));
 sky130_fd_sc_hd__o22ai_1 _27605_ (.A1(_08234_),
    .A2(_08235_),
    .B1(_08236_),
    .B2(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__nor2_1 _27606_ (.A(net2709),
    .B(_08238_),
    .Y(_08239_));
 sky130_fd_sc_hd__nor2_1 _27607_ (.A(net2435),
    .B(_08239_),
    .Y(_08240_));
 sky130_fd_sc_hd__o21ai_0 _27608_ (.A1(net2415),
    .A2(_08233_),
    .B1(_08240_),
    .Y(_08241_));
 sky130_fd_sc_hd__a32oi_1 _27609_ (.A1(_08206_),
    .A2(_08217_),
    .A3(net2694),
    .B1(_08228_),
    .B2(_08241_),
    .Y(_00034_));
 sky130_fd_sc_hd__nor2_1 _27610_ (.A(\inst$top.soc.cpu.gprf.mem[7][12] ),
    .B(net2408),
    .Y(_08242_));
 sky130_fd_sc_hd__o21ai_0 _27611_ (.A1(net2817),
    .A2(\inst$top.soc.cpu.gprf.mem[6][12] ),
    .B1(net2748),
    .Y(_08243_));
 sky130_fd_sc_hd__nor2_1 _27612_ (.A(net2815),
    .B(\inst$top.soc.cpu.gprf.mem[4][12] ),
    .Y(_08244_));
 sky130_fd_sc_hd__o21ai_0 _27613_ (.A1(\inst$top.soc.cpu.gprf.mem[5][12] ),
    .A2(net2408),
    .B1(net2344),
    .Y(_08245_));
 sky130_fd_sc_hd__o221ai_1 _27614_ (.A1(_08242_),
    .A2(_08243_),
    .B1(_08244_),
    .B2(_08245_),
    .C1(net2715),
    .Y(_08246_));
 sky130_fd_sc_hd__nor2_1 _27615_ (.A(\inst$top.soc.cpu.gprf.mem[3][12] ),
    .B(net2408),
    .Y(_08247_));
 sky130_fd_sc_hd__o21ai_0 _27616_ (.A1(net2817),
    .A2(\inst$top.soc.cpu.gprf.mem[2][12] ),
    .B1(net2748),
    .Y(_08248_));
 sky130_fd_sc_hd__nor2_1 _27617_ (.A(net2815),
    .B(\inst$top.soc.cpu.gprf.mem[0][12] ),
    .Y(_08249_));
 sky130_fd_sc_hd__o21ai_0 _27618_ (.A1(\inst$top.soc.cpu.gprf.mem[1][12] ),
    .A2(net2408),
    .B1(net2344),
    .Y(_08250_));
 sky130_fd_sc_hd__o221ai_1 _27619_ (.A1(_08247_),
    .A2(_08248_),
    .B1(_08249_),
    .B2(_08250_),
    .C1(net2427),
    .Y(_08251_));
 sky130_fd_sc_hd__nand3_1 _27620_ (.A(_08246_),
    .B(_08251_),
    .C(net2440),
    .Y(_08252_));
 sky130_fd_sc_hd__nor2_1 _27621_ (.A(\inst$top.soc.cpu.gprf.mem[11][12] ),
    .B(net2408),
    .Y(_08253_));
 sky130_fd_sc_hd__o21ai_0 _27622_ (.A1(net2817),
    .A2(\inst$top.soc.cpu.gprf.mem[10][12] ),
    .B1(net2748),
    .Y(_08254_));
 sky130_fd_sc_hd__nor2_1 _27623_ (.A(net2815),
    .B(\inst$top.soc.cpu.gprf.mem[8][12] ),
    .Y(_08255_));
 sky130_fd_sc_hd__o21ai_0 _27625_ (.A1(\inst$top.soc.cpu.gprf.mem[9][12] ),
    .A2(net2408),
    .B1(net2344),
    .Y(_08257_));
 sky130_fd_sc_hd__o22ai_1 _27626_ (.A1(_08253_),
    .A2(_08254_),
    .B1(_08255_),
    .B2(_08257_),
    .Y(_08258_));
 sky130_fd_sc_hd__nor2_1 _27627_ (.A(\inst$top.soc.cpu.gprf.mem[15][12] ),
    .B(net2409),
    .Y(_08259_));
 sky130_fd_sc_hd__o21ai_0 _27628_ (.A1(net2816),
    .A2(\inst$top.soc.cpu.gprf.mem[14][12] ),
    .B1(net2748),
    .Y(_08260_));
 sky130_fd_sc_hd__nor2_1 _27629_ (.A(net2816),
    .B(\inst$top.soc.cpu.gprf.mem[12][12] ),
    .Y(_08261_));
 sky130_fd_sc_hd__o21ai_0 _27630_ (.A1(\inst$top.soc.cpu.gprf.mem[13][12] ),
    .A2(net2409),
    .B1(net2345),
    .Y(_08262_));
 sky130_fd_sc_hd__o22ai_1 _27631_ (.A1(_08259_),
    .A2(_08260_),
    .B1(_08261_),
    .B2(_08262_),
    .Y(_08263_));
 sky130_fd_sc_hd__nor2_1 _27632_ (.A(net2428),
    .B(_08263_),
    .Y(_08264_));
 sky130_fd_sc_hd__nor2_1 _27633_ (.A(net2440),
    .B(_08264_),
    .Y(_08265_));
 sky130_fd_sc_hd__o21ai_0 _27634_ (.A1(net2715),
    .A2(_08258_),
    .B1(_08265_),
    .Y(_08266_));
 sky130_fd_sc_hd__nor2_1 _27635_ (.A(\inst$top.soc.cpu.gprf.mem[31][12] ),
    .B(net2408),
    .Y(_08267_));
 sky130_fd_sc_hd__o21ai_0 _27636_ (.A1(net2815),
    .A2(\inst$top.soc.cpu.gprf.mem[30][12] ),
    .B1(net2748),
    .Y(_08268_));
 sky130_fd_sc_hd__nor2_1 _27637_ (.A(net2815),
    .B(\inst$top.soc.cpu.gprf.mem[28][12] ),
    .Y(_08269_));
 sky130_fd_sc_hd__o21ai_0 _27638_ (.A1(\inst$top.soc.cpu.gprf.mem[29][12] ),
    .A2(net2408),
    .B1(net2344),
    .Y(_08270_));
 sky130_fd_sc_hd__o22ai_1 _27639_ (.A1(_08267_),
    .A2(_08268_),
    .B1(_08269_),
    .B2(_08270_),
    .Y(_08271_));
 sky130_fd_sc_hd__nor2_1 _27640_ (.A(net2427),
    .B(_08271_),
    .Y(_08272_));
 sky130_fd_sc_hd__nor2_1 _27641_ (.A(\inst$top.soc.cpu.gprf.mem[27][12] ),
    .B(net2408),
    .Y(_08273_));
 sky130_fd_sc_hd__o21ai_0 _27642_ (.A1(net2815),
    .A2(\inst$top.soc.cpu.gprf.mem[26][12] ),
    .B1(net2748),
    .Y(_08274_));
 sky130_fd_sc_hd__nor2_1 _27643_ (.A(net2815),
    .B(\inst$top.soc.cpu.gprf.mem[24][12] ),
    .Y(_08275_));
 sky130_fd_sc_hd__o21ai_0 _27644_ (.A1(\inst$top.soc.cpu.gprf.mem[25][12] ),
    .A2(net2408),
    .B1(net2344),
    .Y(_08276_));
 sky130_fd_sc_hd__o22ai_1 _27645_ (.A1(_08273_),
    .A2(_08274_),
    .B1(_08275_),
    .B2(_08276_),
    .Y(_08277_));
 sky130_fd_sc_hd__o21ai_0 _27646_ (.A1(net2715),
    .A2(_08277_),
    .B1(net2699),
    .Y(_08278_));
 sky130_fd_sc_hd__nor2_1 _27647_ (.A(\inst$top.soc.cpu.gprf.mem[23][12] ),
    .B(net2410),
    .Y(_08279_));
 sky130_fd_sc_hd__o21ai_0 _27648_ (.A1(net2816),
    .A2(\inst$top.soc.cpu.gprf.mem[22][12] ),
    .B1(net2749),
    .Y(_08280_));
 sky130_fd_sc_hd__nor2_1 _27649_ (.A(net2816),
    .B(\inst$top.soc.cpu.gprf.mem[20][12] ),
    .Y(_08281_));
 sky130_fd_sc_hd__o21ai_0 _27650_ (.A1(\inst$top.soc.cpu.gprf.mem[21][12] ),
    .A2(net2410),
    .B1(net2344),
    .Y(_08282_));
 sky130_fd_sc_hd__o221ai_1 _27651_ (.A1(_08279_),
    .A2(_08280_),
    .B1(_08281_),
    .B2(_08282_),
    .C1(net2715),
    .Y(_08283_));
 sky130_fd_sc_hd__nor2_1 _27652_ (.A(\inst$top.soc.cpu.gprf.mem[19][12] ),
    .B(net2410),
    .Y(_08284_));
 sky130_fd_sc_hd__o21ai_0 _27653_ (.A1(net2815),
    .A2(\inst$top.soc.cpu.gprf.mem[18][12] ),
    .B1(net2748),
    .Y(_08285_));
 sky130_fd_sc_hd__nor2_1 _27654_ (.A(net2815),
    .B(\inst$top.soc.cpu.gprf.mem[16][12] ),
    .Y(_08286_));
 sky130_fd_sc_hd__o21ai_0 _27655_ (.A1(\inst$top.soc.cpu.gprf.mem[17][12] ),
    .A2(net2410),
    .B1(net2344),
    .Y(_08287_));
 sky130_fd_sc_hd__o221ai_1 _27656_ (.A1(_08284_),
    .A2(_08285_),
    .B1(_08286_),
    .B2(_08287_),
    .C1(net2428),
    .Y(_08288_));
 sky130_fd_sc_hd__nand3_1 _27657_ (.A(_08283_),
    .B(_08288_),
    .C(net2440),
    .Y(_08289_));
 sky130_fd_sc_hd__o21ai_0 _27658_ (.A1(_08272_),
    .A2(_08278_),
    .B1(_08289_),
    .Y(_08290_));
 sky130_fd_sc_hd__nor2_1 _27659_ (.A(net2443),
    .B(_08290_),
    .Y(_08291_));
 sky130_fd_sc_hd__a31oi_1 _27660_ (.A1(net2443),
    .A2(_08252_),
    .A3(_08266_),
    .B1(_08291_),
    .Y(_00035_));
 sky130_fd_sc_hd__nor2_1 _27661_ (.A(\inst$top.soc.cpu.gprf.mem[7][13] ),
    .B(net2366),
    .Y(_08292_));
 sky130_fd_sc_hd__o21ai_0 _27662_ (.A1(net2769),
    .A2(\inst$top.soc.cpu.gprf.mem[6][13] ),
    .B1(net2725),
    .Y(_08293_));
 sky130_fd_sc_hd__nor2_1 _27663_ (.A(net2769),
    .B(\inst$top.soc.cpu.gprf.mem[4][13] ),
    .Y(_08294_));
 sky130_fd_sc_hd__o21ai_0 _27664_ (.A1(\inst$top.soc.cpu.gprf.mem[5][13] ),
    .A2(net2366),
    .B1(net2323),
    .Y(_08295_));
 sky130_fd_sc_hd__o221ai_1 _27665_ (.A1(_08292_),
    .A2(_08293_),
    .B1(_08294_),
    .B2(_08295_),
    .C1(net2704),
    .Y(_08296_));
 sky130_fd_sc_hd__nor2_1 _27666_ (.A(\inst$top.soc.cpu.gprf.mem[3][13] ),
    .B(net2365),
    .Y(_08297_));
 sky130_fd_sc_hd__o21ai_0 _27667_ (.A1(net2769),
    .A2(\inst$top.soc.cpu.gprf.mem[2][13] ),
    .B1(net2725),
    .Y(_08298_));
 sky130_fd_sc_hd__nor2_1 _27668_ (.A(net2768),
    .B(\inst$top.soc.cpu.gprf.mem[0][13] ),
    .Y(_08299_));
 sky130_fd_sc_hd__o21ai_0 _27669_ (.A1(\inst$top.soc.cpu.gprf.mem[1][13] ),
    .A2(net2365),
    .B1(net2323),
    .Y(_08300_));
 sky130_fd_sc_hd__o221ai_1 _27670_ (.A1(_08297_),
    .A2(_08298_),
    .B1(_08299_),
    .B2(_08300_),
    .C1(net2418),
    .Y(_08301_));
 sky130_fd_sc_hd__nand3_1 _27671_ (.A(_08296_),
    .B(_08301_),
    .C(net2433),
    .Y(_08302_));
 sky130_fd_sc_hd__nor2_1 _27672_ (.A(\inst$top.soc.cpu.gprf.mem[11][13] ),
    .B(net2365),
    .Y(_08303_));
 sky130_fd_sc_hd__o21ai_0 _27673_ (.A1(net2768),
    .A2(\inst$top.soc.cpu.gprf.mem[10][13] ),
    .B1(net2725),
    .Y(_08304_));
 sky130_fd_sc_hd__nor2_1 _27674_ (.A(net2768),
    .B(\inst$top.soc.cpu.gprf.mem[8][13] ),
    .Y(_08305_));
 sky130_fd_sc_hd__o21ai_0 _27675_ (.A1(\inst$top.soc.cpu.gprf.mem[9][13] ),
    .A2(net2365),
    .B1(net2323),
    .Y(_08306_));
 sky130_fd_sc_hd__o221ai_1 _27676_ (.A1(_08303_),
    .A2(_08304_),
    .B1(_08305_),
    .B2(_08306_),
    .C1(net2418),
    .Y(_08307_));
 sky130_fd_sc_hd__nor2_1 _27677_ (.A(\inst$top.soc.cpu.gprf.mem[15][13] ),
    .B(net2365),
    .Y(_08308_));
 sky130_fd_sc_hd__o21ai_0 _27678_ (.A1(net2768),
    .A2(\inst$top.soc.cpu.gprf.mem[14][13] ),
    .B1(net2725),
    .Y(_08309_));
 sky130_fd_sc_hd__nor2_1 _27679_ (.A(net2768),
    .B(\inst$top.soc.cpu.gprf.mem[12][13] ),
    .Y(_08310_));
 sky130_fd_sc_hd__o21ai_0 _27680_ (.A1(\inst$top.soc.cpu.gprf.mem[13][13] ),
    .A2(net2365),
    .B1(net2323),
    .Y(_08311_));
 sky130_fd_sc_hd__o221ai_1 _27681_ (.A1(_08308_),
    .A2(_08309_),
    .B1(_08310_),
    .B2(_08311_),
    .C1(net2704),
    .Y(_08312_));
 sky130_fd_sc_hd__nand3_1 _27682_ (.A(_08307_),
    .B(_08312_),
    .C(net2697),
    .Y(_08313_));
 sky130_fd_sc_hd__nor2_1 _27683_ (.A(\inst$top.soc.cpu.gprf.mem[31][13] ),
    .B(net2367),
    .Y(_08314_));
 sky130_fd_sc_hd__o21ai_0 _27684_ (.A1(net2769),
    .A2(\inst$top.soc.cpu.gprf.mem[30][13] ),
    .B1(net2727),
    .Y(_08315_));
 sky130_fd_sc_hd__nor2_1 _27685_ (.A(net2769),
    .B(\inst$top.soc.cpu.gprf.mem[28][13] ),
    .Y(_08316_));
 sky130_fd_sc_hd__o21ai_0 _27686_ (.A1(\inst$top.soc.cpu.gprf.mem[29][13] ),
    .A2(net2367),
    .B1(net2325),
    .Y(_08317_));
 sky130_fd_sc_hd__o221ai_1 _27687_ (.A1(_08314_),
    .A2(_08315_),
    .B1(_08316_),
    .B2(_08317_),
    .C1(net2704),
    .Y(_08318_));
 sky130_fd_sc_hd__nor2_1 _27688_ (.A(\inst$top.soc.cpu.gprf.mem[27][13] ),
    .B(net2366),
    .Y(_08319_));
 sky130_fd_sc_hd__o21ai_0 _27689_ (.A1(net2769),
    .A2(\inst$top.soc.cpu.gprf.mem[26][13] ),
    .B1(net2725),
    .Y(_08320_));
 sky130_fd_sc_hd__nor2_1 _27690_ (.A(net2769),
    .B(\inst$top.soc.cpu.gprf.mem[24][13] ),
    .Y(_08321_));
 sky130_fd_sc_hd__o21ai_0 _27692_ (.A1(\inst$top.soc.cpu.gprf.mem[25][13] ),
    .A2(net2366),
    .B1(net2325),
    .Y(_08323_));
 sky130_fd_sc_hd__o221ai_1 _27693_ (.A1(_08319_),
    .A2(_08320_),
    .B1(_08321_),
    .B2(_08323_),
    .C1(net2418),
    .Y(_08324_));
 sky130_fd_sc_hd__a31oi_1 _27694_ (.A1(_08318_),
    .A2(_08324_),
    .A3(net2697),
    .B1(net2442),
    .Y(_08325_));
 sky130_fd_sc_hd__nor2_1 _27695_ (.A(\inst$top.soc.cpu.gprf.mem[23][13] ),
    .B(net2365),
    .Y(_08326_));
 sky130_fd_sc_hd__o21ai_0 _27696_ (.A1(net2770),
    .A2(\inst$top.soc.cpu.gprf.mem[22][13] ),
    .B1(net2725),
    .Y(_08327_));
 sky130_fd_sc_hd__nor2_1 _27697_ (.A(net2769),
    .B(\inst$top.soc.cpu.gprf.mem[20][13] ),
    .Y(_08328_));
 sky130_fd_sc_hd__o21ai_0 _27698_ (.A1(\inst$top.soc.cpu.gprf.mem[21][13] ),
    .A2(net2367),
    .B1(net2323),
    .Y(_08329_));
 sky130_fd_sc_hd__o221ai_1 _27699_ (.A1(_08326_),
    .A2(_08327_),
    .B1(_08328_),
    .B2(_08329_),
    .C1(net2704),
    .Y(_08330_));
 sky130_fd_sc_hd__nor2_1 _27700_ (.A(\inst$top.soc.cpu.gprf.mem[19][13] ),
    .B(net2367),
    .Y(_08331_));
 sky130_fd_sc_hd__o21ai_0 _27701_ (.A1(net2768),
    .A2(\inst$top.soc.cpu.gprf.mem[18][13] ),
    .B1(net2725),
    .Y(_08332_));
 sky130_fd_sc_hd__nor2_1 _27702_ (.A(net2770),
    .B(\inst$top.soc.cpu.gprf.mem[16][13] ),
    .Y(_08333_));
 sky130_fd_sc_hd__o21ai_0 _27703_ (.A1(\inst$top.soc.cpu.gprf.mem[17][13] ),
    .A2(net2365),
    .B1(net2323),
    .Y(_08334_));
 sky130_fd_sc_hd__o221ai_1 _27704_ (.A1(_08331_),
    .A2(_08332_),
    .B1(_08333_),
    .B2(_08334_),
    .C1(net2418),
    .Y(_08335_));
 sky130_fd_sc_hd__nand3_1 _27705_ (.A(_08330_),
    .B(_08335_),
    .C(net2433),
    .Y(_08336_));
 sky130_fd_sc_hd__a32oi_1 _27706_ (.A1(_08302_),
    .A2(_08313_),
    .A3(net2442),
    .B1(_08325_),
    .B2(_08336_),
    .Y(_00036_));
 sky130_fd_sc_hd__nor2_1 _27707_ (.A(\inst$top.soc.cpu.gprf.mem[31][14] ),
    .B(net2395),
    .Y(_08337_));
 sky130_fd_sc_hd__o21ai_0 _27708_ (.A1(net2797),
    .A2(\inst$top.soc.cpu.gprf.mem[30][14] ),
    .B1(net2741),
    .Y(_08338_));
 sky130_fd_sc_hd__nor2_1 _27709_ (.A(net2800),
    .B(\inst$top.soc.cpu.gprf.mem[28][14] ),
    .Y(_08339_));
 sky130_fd_sc_hd__o21ai_0 _27710_ (.A1(\inst$top.soc.cpu.gprf.mem[29][14] ),
    .A2(net2392),
    .B1(net2336),
    .Y(_08340_));
 sky130_fd_sc_hd__o22ai_1 _27711_ (.A1(_08337_),
    .A2(_08338_),
    .B1(_08339_),
    .B2(_08340_),
    .Y(_08341_));
 sky130_fd_sc_hd__nor2_1 _27712_ (.A(\inst$top.soc.cpu.gprf.mem[27][14] ),
    .B(net2395),
    .Y(_08342_));
 sky130_fd_sc_hd__o21ai_0 _27713_ (.A1(net2801),
    .A2(\inst$top.soc.cpu.gprf.mem[26][14] ),
    .B1(net2741),
    .Y(_08343_));
 sky130_fd_sc_hd__nor2_1 _27714_ (.A(net2801),
    .B(\inst$top.soc.cpu.gprf.mem[24][14] ),
    .Y(_08344_));
 sky130_fd_sc_hd__o21ai_0 _27715_ (.A1(\inst$top.soc.cpu.gprf.mem[25][14] ),
    .A2(net2395),
    .B1(net2337),
    .Y(_08345_));
 sky130_fd_sc_hd__o22ai_1 _27716_ (.A1(_08342_),
    .A2(_08343_),
    .B1(_08344_),
    .B2(_08345_),
    .Y(_08346_));
 sky130_fd_sc_hd__nor2_1 _27717_ (.A(net2712),
    .B(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__nor2_1 _27718_ (.A(net2438),
    .B(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__o21ai_0 _27719_ (.A1(net2424),
    .A2(_08341_),
    .B1(_08348_),
    .Y(_08349_));
 sky130_fd_sc_hd__nor2_1 _27720_ (.A(\inst$top.soc.cpu.gprf.mem[23][14] ),
    .B(net2394),
    .Y(_08350_));
 sky130_fd_sc_hd__o21ai_0 _27721_ (.A1(net2799),
    .A2(\inst$top.soc.cpu.gprf.mem[22][14] ),
    .B1(net2742),
    .Y(_08351_));
 sky130_fd_sc_hd__nor2_1 _27722_ (.A(net2799),
    .B(\inst$top.soc.cpu.gprf.mem[20][14] ),
    .Y(_08352_));
 sky130_fd_sc_hd__o21ai_0 _27723_ (.A1(\inst$top.soc.cpu.gprf.mem[21][14] ),
    .A2(net2394),
    .B1(net2338),
    .Y(_08353_));
 sky130_fd_sc_hd__o221ai_1 _27724_ (.A1(_08350_),
    .A2(_08351_),
    .B1(_08352_),
    .B2(_08353_),
    .C1(net2711),
    .Y(_08354_));
 sky130_fd_sc_hd__nor2_1 _27725_ (.A(\inst$top.soc.cpu.gprf.mem[19][14] ),
    .B(net2396),
    .Y(_08355_));
 sky130_fd_sc_hd__o21ai_0 _27726_ (.A1(net2802),
    .A2(\inst$top.soc.cpu.gprf.mem[18][14] ),
    .B1(net2741),
    .Y(_08356_));
 sky130_fd_sc_hd__nor2_1 _27727_ (.A(net2802),
    .B(\inst$top.soc.cpu.gprf.mem[16][14] ),
    .Y(_08357_));
 sky130_fd_sc_hd__o21ai_0 _27728_ (.A1(\inst$top.soc.cpu.gprf.mem[17][14] ),
    .A2(net2396),
    .B1(net2337),
    .Y(_08358_));
 sky130_fd_sc_hd__o221ai_1 _27729_ (.A1(_08355_),
    .A2(_08356_),
    .B1(_08357_),
    .B2(_08358_),
    .C1(net2424),
    .Y(_08359_));
 sky130_fd_sc_hd__nand3_1 _27730_ (.A(_08354_),
    .B(_08359_),
    .C(net2438),
    .Y(_08360_));
 sky130_fd_sc_hd__nor2_1 _27731_ (.A(\inst$top.soc.cpu.gprf.mem[7][14] ),
    .B(net2392),
    .Y(_08361_));
 sky130_fd_sc_hd__o21ai_0 _27732_ (.A1(net2800),
    .A2(\inst$top.soc.cpu.gprf.mem[6][14] ),
    .B1(net2740),
    .Y(_08362_));
 sky130_fd_sc_hd__nor2_1 _27733_ (.A(net2800),
    .B(\inst$top.soc.cpu.gprf.mem[4][14] ),
    .Y(_08363_));
 sky130_fd_sc_hd__o21ai_0 _27734_ (.A1(\inst$top.soc.cpu.gprf.mem[5][14] ),
    .A2(net2392),
    .B1(net2336),
    .Y(_08364_));
 sky130_fd_sc_hd__o221ai_1 _27735_ (.A1(_08361_),
    .A2(_08362_),
    .B1(_08363_),
    .B2(_08364_),
    .C1(net2711),
    .Y(_08365_));
 sky130_fd_sc_hd__nor2_1 _27737_ (.A(\inst$top.soc.cpu.gprf.mem[3][14] ),
    .B(net2395),
    .Y(_08367_));
 sky130_fd_sc_hd__o21ai_0 _27738_ (.A1(net2801),
    .A2(\inst$top.soc.cpu.gprf.mem[2][14] ),
    .B1(net2741),
    .Y(_08368_));
 sky130_fd_sc_hd__nor2_1 _27739_ (.A(net2801),
    .B(\inst$top.soc.cpu.gprf.mem[0][14] ),
    .Y(_08369_));
 sky130_fd_sc_hd__o21ai_0 _27740_ (.A1(\inst$top.soc.cpu.gprf.mem[1][14] ),
    .A2(net2394),
    .B1(net2336),
    .Y(_08370_));
 sky130_fd_sc_hd__o221ai_1 _27741_ (.A1(_08367_),
    .A2(_08368_),
    .B1(_08369_),
    .B2(_08370_),
    .C1(net2424),
    .Y(_08371_));
 sky130_fd_sc_hd__a31oi_1 _27742_ (.A1(_08365_),
    .A2(_08371_),
    .A3(net2438),
    .B1(net2692),
    .Y(_08372_));
 sky130_fd_sc_hd__nor2_1 _27743_ (.A(\inst$top.soc.cpu.gprf.mem[15][14] ),
    .B(net2394),
    .Y(_08373_));
 sky130_fd_sc_hd__o21ai_0 _27744_ (.A1(net2799),
    .A2(\inst$top.soc.cpu.gprf.mem[14][14] ),
    .B1(net2740),
    .Y(_08374_));
 sky130_fd_sc_hd__nor2_1 _27745_ (.A(net2799),
    .B(\inst$top.soc.cpu.gprf.mem[12][14] ),
    .Y(_08375_));
 sky130_fd_sc_hd__o21ai_0 _27746_ (.A1(\inst$top.soc.cpu.gprf.mem[13][14] ),
    .A2(net2394),
    .B1(net2336),
    .Y(_08376_));
 sky130_fd_sc_hd__o22ai_1 _27747_ (.A1(_08373_),
    .A2(_08374_),
    .B1(_08375_),
    .B2(_08376_),
    .Y(_08377_));
 sky130_fd_sc_hd__nor2_1 _27748_ (.A(\inst$top.soc.cpu.gprf.mem[11][14] ),
    .B(net2396),
    .Y(_08378_));
 sky130_fd_sc_hd__o21ai_0 _27749_ (.A1(net2802),
    .A2(\inst$top.soc.cpu.gprf.mem[10][14] ),
    .B1(net2741),
    .Y(_08379_));
 sky130_fd_sc_hd__nor2_1 _27750_ (.A(net2802),
    .B(\inst$top.soc.cpu.gprf.mem[8][14] ),
    .Y(_08380_));
 sky130_fd_sc_hd__o21ai_0 _27751_ (.A1(\inst$top.soc.cpu.gprf.mem[9][14] ),
    .A2(net2396),
    .B1(net2337),
    .Y(_08381_));
 sky130_fd_sc_hd__o22ai_1 _27752_ (.A1(_08378_),
    .A2(_08379_),
    .B1(_08380_),
    .B2(_08381_),
    .Y(_08382_));
 sky130_fd_sc_hd__nor2_1 _27753_ (.A(net2712),
    .B(_08382_),
    .Y(_08383_));
 sky130_fd_sc_hd__nor2_1 _27754_ (.A(net2438),
    .B(_08383_),
    .Y(_08384_));
 sky130_fd_sc_hd__o21ai_0 _27755_ (.A1(net2424),
    .A2(_08377_),
    .B1(_08384_),
    .Y(_08385_));
 sky130_fd_sc_hd__a32oi_1 _27756_ (.A1(net2692),
    .A2(_08349_),
    .A3(_08360_),
    .B1(_08372_),
    .B2(_08385_),
    .Y(_00037_));
 sky130_fd_sc_hd__nor2_1 _27757_ (.A(\inst$top.soc.cpu.gprf.mem[31][15] ),
    .B(net2396),
    .Y(_08386_));
 sky130_fd_sc_hd__o21ai_0 _27758_ (.A1(net2802),
    .A2(\inst$top.soc.cpu.gprf.mem[30][15] ),
    .B1(net2742),
    .Y(_08387_));
 sky130_fd_sc_hd__nor2_1 _27759_ (.A(net2803),
    .B(\inst$top.soc.cpu.gprf.mem[28][15] ),
    .Y(_08388_));
 sky130_fd_sc_hd__o21ai_0 _27760_ (.A1(\inst$top.soc.cpu.gprf.mem[29][15] ),
    .A2(net2397),
    .B1(net2337),
    .Y(_08389_));
 sky130_fd_sc_hd__o22ai_1 _27761_ (.A1(_08386_),
    .A2(_08387_),
    .B1(_08388_),
    .B2(_08389_),
    .Y(_08390_));
 sky130_fd_sc_hd__nor2_1 _27762_ (.A(\inst$top.soc.cpu.gprf.mem[27][15] ),
    .B(net2395),
    .Y(_08391_));
 sky130_fd_sc_hd__o21ai_0 _27763_ (.A1(net2801),
    .A2(\inst$top.soc.cpu.gprf.mem[26][15] ),
    .B1(net2741),
    .Y(_08392_));
 sky130_fd_sc_hd__nor2_1 _27764_ (.A(net2803),
    .B(\inst$top.soc.cpu.gprf.mem[24][15] ),
    .Y(_08393_));
 sky130_fd_sc_hd__o21ai_0 _27765_ (.A1(\inst$top.soc.cpu.gprf.mem[25][15] ),
    .A2(net2395),
    .B1(net2337),
    .Y(_08394_));
 sky130_fd_sc_hd__o22ai_1 _27766_ (.A1(_08391_),
    .A2(_08392_),
    .B1(_08393_),
    .B2(_08394_),
    .Y(_08395_));
 sky130_fd_sc_hd__nor2_1 _27767_ (.A(net2711),
    .B(_08395_),
    .Y(_08396_));
 sky130_fd_sc_hd__nor2_1 _27768_ (.A(net2438),
    .B(_08396_),
    .Y(_08397_));
 sky130_fd_sc_hd__o21ai_0 _27769_ (.A1(net2424),
    .A2(_08390_),
    .B1(_08397_),
    .Y(_08398_));
 sky130_fd_sc_hd__nor2_1 _27770_ (.A(\inst$top.soc.cpu.gprf.mem[23][15] ),
    .B(net2396),
    .Y(_08399_));
 sky130_fd_sc_hd__o21ai_0 _27771_ (.A1(net2802),
    .A2(\inst$top.soc.cpu.gprf.mem[22][15] ),
    .B1(net2741),
    .Y(_08400_));
 sky130_fd_sc_hd__nor2_1 _27772_ (.A(net2802),
    .B(\inst$top.soc.cpu.gprf.mem[20][15] ),
    .Y(_08401_));
 sky130_fd_sc_hd__o21ai_0 _27773_ (.A1(\inst$top.soc.cpu.gprf.mem[21][15] ),
    .A2(net2396),
    .B1(net2337),
    .Y(_08402_));
 sky130_fd_sc_hd__o221ai_1 _27774_ (.A1(_08399_),
    .A2(_08400_),
    .B1(_08401_),
    .B2(_08402_),
    .C1(net2712),
    .Y(_08403_));
 sky130_fd_sc_hd__nor2_1 _27775_ (.A(\inst$top.soc.cpu.gprf.mem[19][15] ),
    .B(net2396),
    .Y(_08404_));
 sky130_fd_sc_hd__o21ai_0 _27776_ (.A1(net2803),
    .A2(\inst$top.soc.cpu.gprf.mem[18][15] ),
    .B1(net2741),
    .Y(_08405_));
 sky130_fd_sc_hd__nor2_1 _27777_ (.A(net2803),
    .B(\inst$top.soc.cpu.gprf.mem[16][15] ),
    .Y(_08406_));
 sky130_fd_sc_hd__o21ai_0 _27778_ (.A1(\inst$top.soc.cpu.gprf.mem[17][15] ),
    .A2(net2397),
    .B1(net2337),
    .Y(_08407_));
 sky130_fd_sc_hd__o221ai_1 _27779_ (.A1(_08404_),
    .A2(_08405_),
    .B1(_08406_),
    .B2(_08407_),
    .C1(net2424),
    .Y(_08408_));
 sky130_fd_sc_hd__nand3_1 _27780_ (.A(_08403_),
    .B(_08408_),
    .C(net2438),
    .Y(_08409_));
 sky130_fd_sc_hd__nor2_1 _27781_ (.A(\inst$top.soc.cpu.gprf.mem[11][15] ),
    .B(net2396),
    .Y(_08410_));
 sky130_fd_sc_hd__o21ai_0 _27782_ (.A1(net2802),
    .A2(\inst$top.soc.cpu.gprf.mem[10][15] ),
    .B1(net2742),
    .Y(_08411_));
 sky130_fd_sc_hd__nor2_1 _27783_ (.A(net2802),
    .B(\inst$top.soc.cpu.gprf.mem[8][15] ),
    .Y(_08412_));
 sky130_fd_sc_hd__o21ai_0 _27785_ (.A1(\inst$top.soc.cpu.gprf.mem[9][15] ),
    .A2(net2396),
    .B1(net2338),
    .Y(_08414_));
 sky130_fd_sc_hd__o221ai_1 _27786_ (.A1(_08410_),
    .A2(_08411_),
    .B1(_08412_),
    .B2(_08414_),
    .C1(net2425),
    .Y(_08415_));
 sky130_fd_sc_hd__nor2_1 _27787_ (.A(\inst$top.soc.cpu.gprf.mem[15][15] ),
    .B(net2397),
    .Y(_08416_));
 sky130_fd_sc_hd__o21ai_0 _27788_ (.A1(net2803),
    .A2(\inst$top.soc.cpu.gprf.mem[14][15] ),
    .B1(net2742),
    .Y(_08417_));
 sky130_fd_sc_hd__nor2_1 _27789_ (.A(net2803),
    .B(\inst$top.soc.cpu.gprf.mem[12][15] ),
    .Y(_08418_));
 sky130_fd_sc_hd__o21ai_0 _27790_ (.A1(\inst$top.soc.cpu.gprf.mem[13][15] ),
    .A2(net2397),
    .B1(net2338),
    .Y(_08419_));
 sky130_fd_sc_hd__o221ai_1 _27791_ (.A1(_08416_),
    .A2(_08417_),
    .B1(_08418_),
    .B2(_08419_),
    .C1(net2711),
    .Y(_08420_));
 sky130_fd_sc_hd__a31oi_1 _27792_ (.A1(_08415_),
    .A2(_08420_),
    .A3(net2698),
    .B1(net2692),
    .Y(_08421_));
 sky130_fd_sc_hd__nor2_1 _27793_ (.A(\inst$top.soc.cpu.gprf.mem[7][15] ),
    .B(net2395),
    .Y(_08422_));
 sky130_fd_sc_hd__o21ai_0 _27794_ (.A1(net2801),
    .A2(\inst$top.soc.cpu.gprf.mem[6][15] ),
    .B1(net2741),
    .Y(_08423_));
 sky130_fd_sc_hd__nor2_1 _27795_ (.A(net2801),
    .B(\inst$top.soc.cpu.gprf.mem[4][15] ),
    .Y(_08424_));
 sky130_fd_sc_hd__o21ai_0 _27796_ (.A1(\inst$top.soc.cpu.gprf.mem[5][15] ),
    .A2(net2395),
    .B1(net2337),
    .Y(_08425_));
 sky130_fd_sc_hd__o221ai_1 _27797_ (.A1(_08422_),
    .A2(_08423_),
    .B1(_08424_),
    .B2(_08425_),
    .C1(net2712),
    .Y(_08426_));
 sky130_fd_sc_hd__nor2_1 _27798_ (.A(\inst$top.soc.cpu.gprf.mem[3][15] ),
    .B(net2397),
    .Y(_08427_));
 sky130_fd_sc_hd__o21ai_0 _27799_ (.A1(net2801),
    .A2(\inst$top.soc.cpu.gprf.mem[2][15] ),
    .B1(net2741),
    .Y(_08428_));
 sky130_fd_sc_hd__nor2_1 _27800_ (.A(net2803),
    .B(\inst$top.soc.cpu.gprf.mem[0][15] ),
    .Y(_08429_));
 sky130_fd_sc_hd__o21ai_0 _27801_ (.A1(\inst$top.soc.cpu.gprf.mem[1][15] ),
    .A2(net2395),
    .B1(net2337),
    .Y(_08430_));
 sky130_fd_sc_hd__o221ai_1 _27802_ (.A1(_08427_),
    .A2(_08428_),
    .B1(_08429_),
    .B2(_08430_),
    .C1(net2425),
    .Y(_08431_));
 sky130_fd_sc_hd__nand3_1 _27803_ (.A(_08426_),
    .B(_08431_),
    .C(net2438),
    .Y(_08432_));
 sky130_fd_sc_hd__a32oi_1 _27804_ (.A1(net2692),
    .A2(_08398_),
    .A3(_08409_),
    .B1(_08421_),
    .B2(_08432_),
    .Y(_00038_));
 sky130_fd_sc_hd__nor2_1 _27805_ (.A(\inst$top.soc.cpu.gprf.mem[23][16] ),
    .B(net2400),
    .Y(_08433_));
 sky130_fd_sc_hd__o21ai_0 _27806_ (.A1(net2810),
    .A2(\inst$top.soc.cpu.gprf.mem[22][16] ),
    .B1(net2744),
    .Y(_08434_));
 sky130_fd_sc_hd__nor2_1 _27807_ (.A(net2808),
    .B(\inst$top.soc.cpu.gprf.mem[20][16] ),
    .Y(_08435_));
 sky130_fd_sc_hd__o21ai_0 _27808_ (.A1(\inst$top.soc.cpu.gprf.mem[21][16] ),
    .A2(net2400),
    .B1(net2341),
    .Y(_08436_));
 sky130_fd_sc_hd__o221ai_1 _27809_ (.A1(_08433_),
    .A2(_08434_),
    .B1(_08435_),
    .B2(_08436_),
    .C1(net2713),
    .Y(_08437_));
 sky130_fd_sc_hd__nor2_1 _27810_ (.A(\inst$top.soc.cpu.gprf.mem[19][16] ),
    .B(net2400),
    .Y(_08438_));
 sky130_fd_sc_hd__o21ai_0 _27811_ (.A1(net2810),
    .A2(\inst$top.soc.cpu.gprf.mem[18][16] ),
    .B1(net2744),
    .Y(_08439_));
 sky130_fd_sc_hd__nor2_1 _27812_ (.A(net2808),
    .B(\inst$top.soc.cpu.gprf.mem[16][16] ),
    .Y(_08440_));
 sky130_fd_sc_hd__o21ai_0 _27813_ (.A1(\inst$top.soc.cpu.gprf.mem[17][16] ),
    .A2(net2400),
    .B1(net2341),
    .Y(_08441_));
 sky130_fd_sc_hd__o221ai_1 _27814_ (.A1(_08438_),
    .A2(_08439_),
    .B1(_08440_),
    .B2(_08441_),
    .C1(net2426),
    .Y(_08442_));
 sky130_fd_sc_hd__nand3_1 _27815_ (.A(_08437_),
    .B(_08442_),
    .C(net2439),
    .Y(_08443_));
 sky130_fd_sc_hd__nor2_1 _27816_ (.A(\inst$top.soc.cpu.gprf.mem[31][16] ),
    .B(net2400),
    .Y(_08444_));
 sky130_fd_sc_hd__o21ai_0 _27817_ (.A1(net2808),
    .A2(\inst$top.soc.cpu.gprf.mem[30][16] ),
    .B1(net2744),
    .Y(_08445_));
 sky130_fd_sc_hd__nor2_1 _27818_ (.A(net2808),
    .B(\inst$top.soc.cpu.gprf.mem[28][16] ),
    .Y(_08446_));
 sky130_fd_sc_hd__o21ai_0 _27819_ (.A1(\inst$top.soc.cpu.gprf.mem[29][16] ),
    .A2(net2400),
    .B1(net2341),
    .Y(_08447_));
 sky130_fd_sc_hd__o22ai_1 _27820_ (.A1(_08444_),
    .A2(_08445_),
    .B1(_08446_),
    .B2(_08447_),
    .Y(_08448_));
 sky130_fd_sc_hd__nor2_1 _27821_ (.A(\inst$top.soc.cpu.gprf.mem[27][16] ),
    .B(net2400),
    .Y(_08449_));
 sky130_fd_sc_hd__o21ai_0 _27822_ (.A1(net2808),
    .A2(\inst$top.soc.cpu.gprf.mem[26][16] ),
    .B1(net2744),
    .Y(_08450_));
 sky130_fd_sc_hd__nor2_1 _27823_ (.A(net2808),
    .B(\inst$top.soc.cpu.gprf.mem[24][16] ),
    .Y(_08451_));
 sky130_fd_sc_hd__o21ai_0 _27824_ (.A1(\inst$top.soc.cpu.gprf.mem[25][16] ),
    .A2(net2384),
    .B1(net2341),
    .Y(_08452_));
 sky130_fd_sc_hd__o22ai_1 _27825_ (.A1(_08449_),
    .A2(_08450_),
    .B1(_08451_),
    .B2(_08452_),
    .Y(_08453_));
 sky130_fd_sc_hd__nor2_1 _27826_ (.A(net2716),
    .B(_08453_),
    .Y(_08454_));
 sky130_fd_sc_hd__nor2_1 _27827_ (.A(net2439),
    .B(_08454_),
    .Y(_08455_));
 sky130_fd_sc_hd__o21ai_0 _27828_ (.A1(net2426),
    .A2(_08448_),
    .B1(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__nor2_1 _27829_ (.A(\inst$top.soc.cpu.gprf.mem[11][16] ),
    .B(net2401),
    .Y(_08457_));
 sky130_fd_sc_hd__o21ai_0 _27830_ (.A1(net2809),
    .A2(\inst$top.soc.cpu.gprf.mem[10][16] ),
    .B1(net2744),
    .Y(_08458_));
 sky130_fd_sc_hd__nor2_1 _27831_ (.A(net2809),
    .B(\inst$top.soc.cpu.gprf.mem[8][16] ),
    .Y(_08459_));
 sky130_fd_sc_hd__o21ai_0 _27832_ (.A1(\inst$top.soc.cpu.gprf.mem[9][16] ),
    .A2(net2400),
    .B1(net2341),
    .Y(_08460_));
 sky130_fd_sc_hd__o22ai_1 _27833_ (.A1(_08457_),
    .A2(_08458_),
    .B1(_08459_),
    .B2(_08460_),
    .Y(_08461_));
 sky130_fd_sc_hd__nor2_1 _27834_ (.A(net2713),
    .B(_08461_),
    .Y(_08462_));
 sky130_fd_sc_hd__nor2_1 _27835_ (.A(\inst$top.soc.cpu.gprf.mem[15][16] ),
    .B(net2400),
    .Y(_08463_));
 sky130_fd_sc_hd__o21ai_0 _27836_ (.A1(net2808),
    .A2(\inst$top.soc.cpu.gprf.mem[14][16] ),
    .B1(net2744),
    .Y(_08464_));
 sky130_fd_sc_hd__nor2_1 _27837_ (.A(net2808),
    .B(\inst$top.soc.cpu.gprf.mem[12][16] ),
    .Y(_08465_));
 sky130_fd_sc_hd__o21ai_0 _27838_ (.A1(\inst$top.soc.cpu.gprf.mem[13][16] ),
    .A2(net2400),
    .B1(net2341),
    .Y(_08466_));
 sky130_fd_sc_hd__o22ai_1 _27839_ (.A1(_08463_),
    .A2(_08464_),
    .B1(_08465_),
    .B2(_08466_),
    .Y(_08467_));
 sky130_fd_sc_hd__o21ai_0 _27840_ (.A1(net2426),
    .A2(_08467_),
    .B1(net2698),
    .Y(_08468_));
 sky130_fd_sc_hd__nor2_1 _27841_ (.A(\inst$top.soc.cpu.gprf.mem[7][16] ),
    .B(net2401),
    .Y(_08469_));
 sky130_fd_sc_hd__o21ai_0 _27842_ (.A1(net2809),
    .A2(\inst$top.soc.cpu.gprf.mem[6][16] ),
    .B1(net2744),
    .Y(_08470_));
 sky130_fd_sc_hd__nor2_1 _27843_ (.A(net2809),
    .B(\inst$top.soc.cpu.gprf.mem[4][16] ),
    .Y(_08471_));
 sky130_fd_sc_hd__o21ai_0 _27844_ (.A1(\inst$top.soc.cpu.gprf.mem[5][16] ),
    .A2(net2401),
    .B1(net2341),
    .Y(_08472_));
 sky130_fd_sc_hd__o221ai_1 _27845_ (.A1(_08469_),
    .A2(_08470_),
    .B1(_08471_),
    .B2(_08472_),
    .C1(net2713),
    .Y(_08473_));
 sky130_fd_sc_hd__nor2_1 _27846_ (.A(\inst$top.soc.cpu.gprf.mem[3][16] ),
    .B(net2401),
    .Y(_08474_));
 sky130_fd_sc_hd__o21ai_0 _27847_ (.A1(net2808),
    .A2(\inst$top.soc.cpu.gprf.mem[2][16] ),
    .B1(net2744),
    .Y(_08475_));
 sky130_fd_sc_hd__nor2_1 _27848_ (.A(net2808),
    .B(\inst$top.soc.cpu.gprf.mem[0][16] ),
    .Y(_08476_));
 sky130_fd_sc_hd__o21ai_0 _27849_ (.A1(\inst$top.soc.cpu.gprf.mem[1][16] ),
    .A2(net2401),
    .B1(net2341),
    .Y(_08477_));
 sky130_fd_sc_hd__o221ai_1 _27850_ (.A1(_08474_),
    .A2(_08475_),
    .B1(_08476_),
    .B2(_08477_),
    .C1(net2428),
    .Y(_08478_));
 sky130_fd_sc_hd__nand3_1 _27851_ (.A(_08473_),
    .B(_08478_),
    .C(net2439),
    .Y(_08479_));
 sky130_fd_sc_hd__o21ai_0 _27852_ (.A1(_08462_),
    .A2(_08468_),
    .B1(_08479_),
    .Y(_08480_));
 sky130_fd_sc_hd__nor2_1 _27853_ (.A(net2693),
    .B(_08480_),
    .Y(_08481_));
 sky130_fd_sc_hd__a31oi_1 _27854_ (.A1(net2693),
    .A2(_08443_),
    .A3(_08456_),
    .B1(_08481_),
    .Y(_00039_));
 sky130_fd_sc_hd__nor2_1 _27855_ (.A(\inst$top.soc.cpu.gprf.mem[15][17] ),
    .B(net2405),
    .Y(_08482_));
 sky130_fd_sc_hd__o21ai_0 _27856_ (.A1(net2812),
    .A2(\inst$top.soc.cpu.gprf.mem[14][17] ),
    .B1(net2746),
    .Y(_08483_));
 sky130_fd_sc_hd__nor2_1 _27857_ (.A(net2812),
    .B(\inst$top.soc.cpu.gprf.mem[12][17] ),
    .Y(_08484_));
 sky130_fd_sc_hd__o21ai_0 _27858_ (.A1(\inst$top.soc.cpu.gprf.mem[13][17] ),
    .A2(net2405),
    .B1(net2343),
    .Y(_08485_));
 sky130_fd_sc_hd__o221ai_1 _27859_ (.A1(_08482_),
    .A2(_08483_),
    .B1(_08484_),
    .B2(_08485_),
    .C1(net2714),
    .Y(_08486_));
 sky130_fd_sc_hd__nor2_1 _27860_ (.A(\inst$top.soc.cpu.gprf.mem[11][17] ),
    .B(net2406),
    .Y(_08487_));
 sky130_fd_sc_hd__o21ai_0 _27861_ (.A1(net2813),
    .A2(\inst$top.soc.cpu.gprf.mem[10][17] ),
    .B1(net2747),
    .Y(_08488_));
 sky130_fd_sc_hd__nor2_1 _27862_ (.A(net2813),
    .B(\inst$top.soc.cpu.gprf.mem[8][17] ),
    .Y(_08489_));
 sky130_fd_sc_hd__o21ai_0 _27863_ (.A1(\inst$top.soc.cpu.gprf.mem[9][17] ),
    .A2(net2406),
    .B1(net2345),
    .Y(_08490_));
 sky130_fd_sc_hd__o221ai_1 _27864_ (.A1(_08487_),
    .A2(_08488_),
    .B1(_08489_),
    .B2(_08490_),
    .C1(net2427),
    .Y(_08491_));
 sky130_fd_sc_hd__nand3_1 _27865_ (.A(_08486_),
    .B(_08491_),
    .C(net2698),
    .Y(_08492_));
 sky130_fd_sc_hd__nor2_1 _27866_ (.A(\inst$top.soc.cpu.gprf.mem[7][17] ),
    .B(net2404),
    .Y(_08493_));
 sky130_fd_sc_hd__o21ai_0 _27867_ (.A1(net2811),
    .A2(\inst$top.soc.cpu.gprf.mem[6][17] ),
    .B1(net2746),
    .Y(_08494_));
 sky130_fd_sc_hd__nor2_1 _27868_ (.A(net2811),
    .B(\inst$top.soc.cpu.gprf.mem[4][17] ),
    .Y(_08495_));
 sky130_fd_sc_hd__o21ai_0 _27869_ (.A1(\inst$top.soc.cpu.gprf.mem[5][17] ),
    .A2(net2404),
    .B1(net2343),
    .Y(_08496_));
 sky130_fd_sc_hd__o221ai_1 _27870_ (.A1(_08493_),
    .A2(_08494_),
    .B1(_08495_),
    .B2(_08496_),
    .C1(net2714),
    .Y(_08497_));
 sky130_fd_sc_hd__nor2_1 _27871_ (.A(\inst$top.soc.cpu.gprf.mem[3][17] ),
    .B(net2407),
    .Y(_08498_));
 sky130_fd_sc_hd__o21ai_0 _27872_ (.A1(net2814),
    .A2(\inst$top.soc.cpu.gprf.mem[2][17] ),
    .B1(net2746),
    .Y(_08499_));
 sky130_fd_sc_hd__nor2_1 _27873_ (.A(net2811),
    .B(\inst$top.soc.cpu.gprf.mem[0][17] ),
    .Y(_08500_));
 sky130_fd_sc_hd__o21ai_0 _27874_ (.A1(\inst$top.soc.cpu.gprf.mem[1][17] ),
    .A2(net2404),
    .B1(net2343),
    .Y(_08501_));
 sky130_fd_sc_hd__o221ai_1 _27875_ (.A1(_08498_),
    .A2(_08499_),
    .B1(_08500_),
    .B2(_08501_),
    .C1(net2427),
    .Y(_08502_));
 sky130_fd_sc_hd__nand3_1 _27876_ (.A(_08497_),
    .B(_08502_),
    .C(net2440),
    .Y(_08503_));
 sky130_fd_sc_hd__nor2_1 _27877_ (.A(\inst$top.soc.cpu.gprf.mem[31][17] ),
    .B(net2404),
    .Y(_08504_));
 sky130_fd_sc_hd__o21ai_0 _27879_ (.A1(net2813),
    .A2(\inst$top.soc.cpu.gprf.mem[30][17] ),
    .B1(net2749),
    .Y(_08506_));
 sky130_fd_sc_hd__nor2_1 _27880_ (.A(net2815),
    .B(\inst$top.soc.cpu.gprf.mem[28][17] ),
    .Y(_08507_));
 sky130_fd_sc_hd__o21ai_0 _27881_ (.A1(\inst$top.soc.cpu.gprf.mem[29][17] ),
    .A2(net2407),
    .B1(net2344),
    .Y(_08508_));
 sky130_fd_sc_hd__o221ai_1 _27882_ (.A1(_08504_),
    .A2(_08506_),
    .B1(_08507_),
    .B2(_08508_),
    .C1(net2714),
    .Y(_08509_));
 sky130_fd_sc_hd__nor2_1 _27883_ (.A(\inst$top.soc.cpu.gprf.mem[27][17] ),
    .B(net2407),
    .Y(_08510_));
 sky130_fd_sc_hd__o21ai_0 _27885_ (.A1(net2814),
    .A2(\inst$top.soc.cpu.gprf.mem[26][17] ),
    .B1(net2747),
    .Y(_08512_));
 sky130_fd_sc_hd__nor2_1 _27886_ (.A(net2811),
    .B(\inst$top.soc.cpu.gprf.mem[24][17] ),
    .Y(_08513_));
 sky130_fd_sc_hd__o21ai_0 _27887_ (.A1(\inst$top.soc.cpu.gprf.mem[25][17] ),
    .A2(net2407),
    .B1(net2343),
    .Y(_08514_));
 sky130_fd_sc_hd__o221ai_1 _27888_ (.A1(_08510_),
    .A2(_08512_),
    .B1(_08513_),
    .B2(_08514_),
    .C1(net2427),
    .Y(_08515_));
 sky130_fd_sc_hd__a31oi_1 _27889_ (.A1(_08509_),
    .A2(_08515_),
    .A3(net2699),
    .B1(net2443),
    .Y(_08516_));
 sky130_fd_sc_hd__nor2_1 _27890_ (.A(\inst$top.soc.cpu.gprf.mem[23][17] ),
    .B(net2409),
    .Y(_08517_));
 sky130_fd_sc_hd__o21ai_0 _27891_ (.A1(net2816),
    .A2(\inst$top.soc.cpu.gprf.mem[22][17] ),
    .B1(net2748),
    .Y(_08518_));
 sky130_fd_sc_hd__nor2_1 _27892_ (.A(net2813),
    .B(\inst$top.soc.cpu.gprf.mem[20][17] ),
    .Y(_08519_));
 sky130_fd_sc_hd__o21ai_0 _27893_ (.A1(\inst$top.soc.cpu.gprf.mem[21][17] ),
    .A2(net2406),
    .B1(net2343),
    .Y(_08520_));
 sky130_fd_sc_hd__o221ai_1 _27894_ (.A1(_08517_),
    .A2(_08518_),
    .B1(_08519_),
    .B2(_08520_),
    .C1(net2715),
    .Y(_08521_));
 sky130_fd_sc_hd__nor2_1 _27895_ (.A(\inst$top.soc.cpu.gprf.mem[19][17] ),
    .B(net2406),
    .Y(_08522_));
 sky130_fd_sc_hd__o21ai_0 _27896_ (.A1(net2813),
    .A2(\inst$top.soc.cpu.gprf.mem[18][17] ),
    .B1(net2746),
    .Y(_08523_));
 sky130_fd_sc_hd__nor2_1 _27897_ (.A(net2813),
    .B(\inst$top.soc.cpu.gprf.mem[16][17] ),
    .Y(_08524_));
 sky130_fd_sc_hd__o21ai_0 _27898_ (.A1(\inst$top.soc.cpu.gprf.mem[17][17] ),
    .A2(net2406),
    .B1(net2345),
    .Y(_08525_));
 sky130_fd_sc_hd__o221ai_1 _27899_ (.A1(_08522_),
    .A2(_08523_),
    .B1(_08524_),
    .B2(_08525_),
    .C1(net2427),
    .Y(_08526_));
 sky130_fd_sc_hd__nand3_1 _27900_ (.A(_08521_),
    .B(_08526_),
    .C(net2440),
    .Y(_08527_));
 sky130_fd_sc_hd__a32oi_1 _27901_ (.A1(_08492_),
    .A2(_08503_),
    .A3(net2443),
    .B1(_08516_),
    .B2(_08527_),
    .Y(_00040_));
 sky130_fd_sc_hd__nor2_1 _27902_ (.A(\inst$top.soc.cpu.gprf.mem[23][18] ),
    .B(net2353),
    .Y(_08528_));
 sky130_fd_sc_hd__o21ai_0 _27903_ (.A1(net2755),
    .A2(\inst$top.soc.cpu.gprf.mem[22][18] ),
    .B1(net2718),
    .Y(_08529_));
 sky130_fd_sc_hd__nor2_1 _27904_ (.A(net2754),
    .B(\inst$top.soc.cpu.gprf.mem[20][18] ),
    .Y(_08530_));
 sky130_fd_sc_hd__o21ai_0 _27905_ (.A1(\inst$top.soc.cpu.gprf.mem[21][18] ),
    .A2(net2354),
    .B1(net2318),
    .Y(_08531_));
 sky130_fd_sc_hd__o221ai_1 _27906_ (.A1(_08528_),
    .A2(_08529_),
    .B1(_08530_),
    .B2(_08531_),
    .C1(net2701),
    .Y(_08532_));
 sky130_fd_sc_hd__nor2_1 _27907_ (.A(\inst$top.soc.cpu.gprf.mem[19][18] ),
    .B(net2364),
    .Y(_08533_));
 sky130_fd_sc_hd__o21ai_0 _27908_ (.A1(net2819),
    .A2(\inst$top.soc.cpu.gprf.mem[18][18] ),
    .B1(net2723),
    .Y(_08534_));
 sky130_fd_sc_hd__nor2_1 _27909_ (.A(net2819),
    .B(\inst$top.soc.cpu.gprf.mem[16][18] ),
    .Y(_08535_));
 sky130_fd_sc_hd__o21ai_0 _27910_ (.A1(\inst$top.soc.cpu.gprf.mem[17][18] ),
    .A2(net2364),
    .B1(net2321),
    .Y(_08536_));
 sky130_fd_sc_hd__o221ai_1 _27911_ (.A1(_08533_),
    .A2(_08534_),
    .B1(_08535_),
    .B2(_08536_),
    .C1(net2415),
    .Y(_08537_));
 sky130_fd_sc_hd__nand3_1 _27912_ (.A(_08532_),
    .B(_08537_),
    .C(net2430),
    .Y(_08538_));
 sky130_fd_sc_hd__nor2_1 _27913_ (.A(\inst$top.soc.cpu.gprf.mem[31][18] ),
    .B(net2354),
    .Y(_08539_));
 sky130_fd_sc_hd__o21ai_0 _27914_ (.A1(net2755),
    .A2(\inst$top.soc.cpu.gprf.mem[30][18] ),
    .B1(net2721),
    .Y(_08540_));
 sky130_fd_sc_hd__nor2_1 _27915_ (.A(net2754),
    .B(\inst$top.soc.cpu.gprf.mem[28][18] ),
    .Y(_08541_));
 sky130_fd_sc_hd__o21ai_0 _27916_ (.A1(\inst$top.soc.cpu.gprf.mem[29][18] ),
    .A2(net2354),
    .B1(net2315),
    .Y(_08542_));
 sky130_fd_sc_hd__o22ai_1 _27917_ (.A1(_08539_),
    .A2(_08540_),
    .B1(_08541_),
    .B2(_08542_),
    .Y(_08543_));
 sky130_fd_sc_hd__nand2_1 _27918_ (.A(net2760),
    .B(\inst$top.soc.cpu.gprf.mem[25][18] ),
    .Y(_08544_));
 sky130_fd_sc_hd__o21ai_0 _27919_ (.A1(net2760),
    .A2(_06930_),
    .B1(_08544_),
    .Y(_08545_));
 sky130_fd_sc_hd__nor2_1 _27920_ (.A(\inst$top.soc.cpu.gprf.mem[27][18] ),
    .B(net2358),
    .Y(_08546_));
 sky130_fd_sc_hd__o21ai_0 _27921_ (.A1(net2760),
    .A2(\inst$top.soc.cpu.gprf.mem[26][18] ),
    .B1(net2720),
    .Y(_08547_));
 sky130_fd_sc_hd__nor2_1 _27922_ (.A(_08546_),
    .B(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__a21oi_1 _27923_ (.A1(net2318),
    .A2(_08545_),
    .B1(_08548_),
    .Y(_08549_));
 sky130_fd_sc_hd__a21oi_1 _27924_ (.A1(_08549_),
    .A2(net2414),
    .B1(net2430),
    .Y(_08550_));
 sky130_fd_sc_hd__o21ai_0 _27925_ (.A1(net2414),
    .A2(_08543_),
    .B1(_08550_),
    .Y(_08551_));
 sky130_fd_sc_hd__nor2_1 _27927_ (.A(\inst$top.soc.cpu.gprf.mem[11][18] ),
    .B(net2362),
    .Y(_08553_));
 sky130_fd_sc_hd__o21ai_0 _27929_ (.A1(net2764),
    .A2(\inst$top.soc.cpu.gprf.mem[10][18] ),
    .B1(net2722),
    .Y(_08555_));
 sky130_fd_sc_hd__nor2_1 _27931_ (.A(net2764),
    .B(\inst$top.soc.cpu.gprf.mem[8][18] ),
    .Y(_08557_));
 sky130_fd_sc_hd__o21ai_0 _27932_ (.A1(\inst$top.soc.cpu.gprf.mem[9][18] ),
    .A2(net2358),
    .B1(net2319),
    .Y(_08558_));
 sky130_fd_sc_hd__o221ai_1 _27933_ (.A1(_08553_),
    .A2(_08555_),
    .B1(_08557_),
    .B2(_08558_),
    .C1(net2416),
    .Y(_08559_));
 sky130_fd_sc_hd__nor2_1 _27934_ (.A(\inst$top.soc.cpu.gprf.mem[15][18] ),
    .B(net2364),
    .Y(_08560_));
 sky130_fd_sc_hd__o21ai_0 _27935_ (.A1(net2763),
    .A2(\inst$top.soc.cpu.gprf.mem[14][18] ),
    .B1(net2722),
    .Y(_08561_));
 sky130_fd_sc_hd__nor2_1 _27936_ (.A(net2763),
    .B(\inst$top.soc.cpu.gprf.mem[12][18] ),
    .Y(_08562_));
 sky130_fd_sc_hd__o21ai_0 _27937_ (.A1(\inst$top.soc.cpu.gprf.mem[13][18] ),
    .A2(net2362),
    .B1(net2319),
    .Y(_08563_));
 sky130_fd_sc_hd__o221ai_1 _27938_ (.A1(_08560_),
    .A2(_08561_),
    .B1(_08562_),
    .B2(_08563_),
    .C1(net2702),
    .Y(_08564_));
 sky130_fd_sc_hd__a31oi_1 _27939_ (.A1(_08559_),
    .A2(_08564_),
    .A3(net2696),
    .B1(net2690),
    .Y(_08565_));
 sky130_fd_sc_hd__nor2_1 _27940_ (.A(\inst$top.soc.cpu.gprf.mem[7][18] ),
    .B(net2358),
    .Y(_08566_));
 sky130_fd_sc_hd__o21ai_0 _27942_ (.A1(net2760),
    .A2(\inst$top.soc.cpu.gprf.mem[6][18] ),
    .B1(net2720),
    .Y(_08568_));
 sky130_fd_sc_hd__nor2_1 _27944_ (.A(net2760),
    .B(\inst$top.soc.cpu.gprf.mem[4][18] ),
    .Y(_08570_));
 sky130_fd_sc_hd__o21ai_0 _27945_ (.A1(\inst$top.soc.cpu.gprf.mem[5][18] ),
    .A2(net2358),
    .B1(net2317),
    .Y(_08571_));
 sky130_fd_sc_hd__o221ai_1 _27946_ (.A1(_08566_),
    .A2(_08568_),
    .B1(_08570_),
    .B2(_08571_),
    .C1(net2702),
    .Y(_08572_));
 sky130_fd_sc_hd__nor2_1 _27947_ (.A(\inst$top.soc.cpu.gprf.mem[3][18] ),
    .B(net2354),
    .Y(_08573_));
 sky130_fd_sc_hd__o21ai_0 _27949_ (.A1(net2761),
    .A2(\inst$top.soc.cpu.gprf.mem[2][18] ),
    .B1(net2720),
    .Y(_08575_));
 sky130_fd_sc_hd__nor2_1 _27950_ (.A(net2760),
    .B(\inst$top.soc.cpu.gprf.mem[0][18] ),
    .Y(_08576_));
 sky130_fd_sc_hd__o21ai_0 _27951_ (.A1(\inst$top.soc.cpu.gprf.mem[1][18] ),
    .A2(net2354),
    .B1(net2318),
    .Y(_08577_));
 sky130_fd_sc_hd__o221ai_1 _27952_ (.A1(_08573_),
    .A2(_08575_),
    .B1(_08576_),
    .B2(_08577_),
    .C1(net2414),
    .Y(_08578_));
 sky130_fd_sc_hd__nand3_1 _27953_ (.A(_08572_),
    .B(_08578_),
    .C(net2430),
    .Y(_08579_));
 sky130_fd_sc_hd__a32oi_1 _27954_ (.A1(net2690),
    .A2(_08538_),
    .A3(_08551_),
    .B1(_08565_),
    .B2(_08579_),
    .Y(_00041_));
 sky130_fd_sc_hd__nor2_1 _27955_ (.A(\inst$top.soc.cpu.gprf.mem[23][19] ),
    .B(net2405),
    .Y(_08580_));
 sky130_fd_sc_hd__o21ai_0 _27956_ (.A1(net2812),
    .A2(\inst$top.soc.cpu.gprf.mem[22][19] ),
    .B1(net2746),
    .Y(_08581_));
 sky130_fd_sc_hd__nor2_1 _27957_ (.A(net2812),
    .B(\inst$top.soc.cpu.gprf.mem[20][19] ),
    .Y(_08582_));
 sky130_fd_sc_hd__o21ai_0 _27958_ (.A1(\inst$top.soc.cpu.gprf.mem[21][19] ),
    .A2(net2405),
    .B1(net2343),
    .Y(_08583_));
 sky130_fd_sc_hd__o221ai_1 _27959_ (.A1(_08580_),
    .A2(_08581_),
    .B1(_08582_),
    .B2(_08583_),
    .C1(net2714),
    .Y(_08584_));
 sky130_fd_sc_hd__nor2_1 _27960_ (.A(\inst$top.soc.cpu.gprf.mem[19][19] ),
    .B(net2405),
    .Y(_08585_));
 sky130_fd_sc_hd__o21ai_0 _27961_ (.A1(net2812),
    .A2(\inst$top.soc.cpu.gprf.mem[18][19] ),
    .B1(net2746),
    .Y(_08586_));
 sky130_fd_sc_hd__nor2_1 _27962_ (.A(net2812),
    .B(\inst$top.soc.cpu.gprf.mem[16][19] ),
    .Y(_08587_));
 sky130_fd_sc_hd__o21ai_0 _27963_ (.A1(\inst$top.soc.cpu.gprf.mem[17][19] ),
    .A2(net2405),
    .B1(net2343),
    .Y(_08588_));
 sky130_fd_sc_hd__o221ai_1 _27964_ (.A1(_08585_),
    .A2(_08586_),
    .B1(_08587_),
    .B2(_08588_),
    .C1(net2427),
    .Y(_08589_));
 sky130_fd_sc_hd__nand3_1 _27965_ (.A(_08584_),
    .B(_08589_),
    .C(net2439),
    .Y(_08590_));
 sky130_fd_sc_hd__nor2_1 _27966_ (.A(\inst$top.soc.cpu.gprf.mem[31][19] ),
    .B(net2404),
    .Y(_08591_));
 sky130_fd_sc_hd__o21ai_0 _27967_ (.A1(net2811),
    .A2(\inst$top.soc.cpu.gprf.mem[30][19] ),
    .B1(net2746),
    .Y(_08592_));
 sky130_fd_sc_hd__nor2_1 _27968_ (.A(net2811),
    .B(\inst$top.soc.cpu.gprf.mem[28][19] ),
    .Y(_08593_));
 sky130_fd_sc_hd__o21ai_0 _27969_ (.A1(\inst$top.soc.cpu.gprf.mem[29][19] ),
    .A2(net2404),
    .B1(net2343),
    .Y(_08594_));
 sky130_fd_sc_hd__o22ai_1 _27970_ (.A1(_08591_),
    .A2(_08592_),
    .B1(_08593_),
    .B2(_08594_),
    .Y(_08595_));
 sky130_fd_sc_hd__nor2_1 _27971_ (.A(\inst$top.soc.cpu.gprf.mem[27][19] ),
    .B(net2404),
    .Y(_08596_));
 sky130_fd_sc_hd__o21ai_0 _27972_ (.A1(net2801),
    .A2(\inst$top.soc.cpu.gprf.mem[26][19] ),
    .B1(net2747),
    .Y(_08597_));
 sky130_fd_sc_hd__nor2_1 _27973_ (.A(net2801),
    .B(\inst$top.soc.cpu.gprf.mem[24][19] ),
    .Y(_08598_));
 sky130_fd_sc_hd__o21ai_0 _27974_ (.A1(\inst$top.soc.cpu.gprf.mem[25][19] ),
    .A2(net2395),
    .B1(net2337),
    .Y(_08599_));
 sky130_fd_sc_hd__o22ai_1 _27975_ (.A1(_08596_),
    .A2(_08597_),
    .B1(_08598_),
    .B2(_08599_),
    .Y(_08600_));
 sky130_fd_sc_hd__nor2_1 _27976_ (.A(net2714),
    .B(_08600_),
    .Y(_08601_));
 sky130_fd_sc_hd__nor2_1 _27977_ (.A(net2440),
    .B(_08601_),
    .Y(_08602_));
 sky130_fd_sc_hd__o21ai_0 _27978_ (.A1(net2427),
    .A2(_08595_),
    .B1(_08602_),
    .Y(_08603_));
 sky130_fd_sc_hd__nor2_1 _27979_ (.A(\inst$top.soc.cpu.gprf.mem[11][19] ),
    .B(net2405),
    .Y(_08604_));
 sky130_fd_sc_hd__o21ai_0 _27980_ (.A1(net2812),
    .A2(\inst$top.soc.cpu.gprf.mem[10][19] ),
    .B1(net2747),
    .Y(_08605_));
 sky130_fd_sc_hd__nor2_1 _27981_ (.A(net2812),
    .B(\inst$top.soc.cpu.gprf.mem[8][19] ),
    .Y(_08606_));
 sky130_fd_sc_hd__o21ai_0 _27982_ (.A1(\inst$top.soc.cpu.gprf.mem[9][19] ),
    .A2(net2405),
    .B1(net2345),
    .Y(_08607_));
 sky130_fd_sc_hd__o22ai_1 _27983_ (.A1(_08604_),
    .A2(_08605_),
    .B1(_08606_),
    .B2(_08607_),
    .Y(_08608_));
 sky130_fd_sc_hd__nor2_1 _27984_ (.A(net2714),
    .B(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__nor2_1 _27985_ (.A(\inst$top.soc.cpu.gprf.mem[15][19] ),
    .B(net2405),
    .Y(_08610_));
 sky130_fd_sc_hd__o21ai_0 _27986_ (.A1(net2812),
    .A2(\inst$top.soc.cpu.gprf.mem[14][19] ),
    .B1(net2747),
    .Y(_08611_));
 sky130_fd_sc_hd__nor2_1 _27987_ (.A(net2812),
    .B(\inst$top.soc.cpu.gprf.mem[12][19] ),
    .Y(_08612_));
 sky130_fd_sc_hd__o21ai_0 _27988_ (.A1(\inst$top.soc.cpu.gprf.mem[13][19] ),
    .A2(net2405),
    .B1(net2345),
    .Y(_08613_));
 sky130_fd_sc_hd__o22ai_1 _27989_ (.A1(_08610_),
    .A2(_08611_),
    .B1(_08612_),
    .B2(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__o21ai_0 _27990_ (.A1(net2427),
    .A2(_08614_),
    .B1(net2698),
    .Y(_08615_));
 sky130_fd_sc_hd__nor2_1 _27991_ (.A(\inst$top.soc.cpu.gprf.mem[7][19] ),
    .B(net2404),
    .Y(_08616_));
 sky130_fd_sc_hd__o21ai_0 _27992_ (.A1(net2811),
    .A2(\inst$top.soc.cpu.gprf.mem[6][19] ),
    .B1(net2746),
    .Y(_08617_));
 sky130_fd_sc_hd__nor2_1 _27993_ (.A(net2811),
    .B(\inst$top.soc.cpu.gprf.mem[4][19] ),
    .Y(_08618_));
 sky130_fd_sc_hd__o21ai_0 _27994_ (.A1(\inst$top.soc.cpu.gprf.mem[5][19] ),
    .A2(net2404),
    .B1(net2343),
    .Y(_08619_));
 sky130_fd_sc_hd__o221ai_1 _27995_ (.A1(_08616_),
    .A2(_08617_),
    .B1(_08618_),
    .B2(_08619_),
    .C1(net2714),
    .Y(_08620_));
 sky130_fd_sc_hd__nor2_1 _27996_ (.A(\inst$top.soc.cpu.gprf.mem[3][19] ),
    .B(net2399),
    .Y(_08621_));
 sky130_fd_sc_hd__o21ai_0 _27997_ (.A1(net2806),
    .A2(\inst$top.soc.cpu.gprf.mem[2][19] ),
    .B1(net2746),
    .Y(_08622_));
 sky130_fd_sc_hd__nor2_1 _27998_ (.A(net2806),
    .B(\inst$top.soc.cpu.gprf.mem[0][19] ),
    .Y(_08623_));
 sky130_fd_sc_hd__o21ai_0 _27999_ (.A1(\inst$top.soc.cpu.gprf.mem[1][19] ),
    .A2(net2399),
    .B1(net2340),
    .Y(_08624_));
 sky130_fd_sc_hd__o221ai_1 _28000_ (.A1(_08621_),
    .A2(_08622_),
    .B1(_08623_),
    .B2(_08624_),
    .C1(net2426),
    .Y(_08625_));
 sky130_fd_sc_hd__nand3_1 _28001_ (.A(_08620_),
    .B(_08625_),
    .C(net2440),
    .Y(_08626_));
 sky130_fd_sc_hd__o21ai_0 _28002_ (.A1(_08609_),
    .A2(_08615_),
    .B1(_08626_),
    .Y(_08627_));
 sky130_fd_sc_hd__nor2_1 _28003_ (.A(net2693),
    .B(_08627_),
    .Y(_08628_));
 sky130_fd_sc_hd__a31oi_1 _28004_ (.A1(net2693),
    .A2(_08590_),
    .A3(_08603_),
    .B1(_08628_),
    .Y(_00042_));
 sky130_fd_sc_hd__nor2_1 _28005_ (.A(\inst$top.soc.cpu.gprf.mem[31][20] ),
    .B(net2379),
    .Y(_08629_));
 sky130_fd_sc_hd__o21ai_0 _28006_ (.A1(net2789),
    .A2(\inst$top.soc.cpu.gprf.mem[30][20] ),
    .B1(net2734),
    .Y(_08630_));
 sky130_fd_sc_hd__nor2_1 _28007_ (.A(net2782),
    .B(\inst$top.soc.cpu.gprf.mem[28][20] ),
    .Y(_08631_));
 sky130_fd_sc_hd__o21ai_0 _28008_ (.A1(\inst$top.soc.cpu.gprf.mem[29][20] ),
    .A2(net2379),
    .B1(net2330),
    .Y(_08632_));
 sky130_fd_sc_hd__o22ai_1 _28009_ (.A1(_08629_),
    .A2(_08630_),
    .B1(_08631_),
    .B2(_08632_),
    .Y(_08633_));
 sky130_fd_sc_hd__nor2_1 _28010_ (.A(\inst$top.soc.cpu.gprf.mem[27][20] ),
    .B(net2382),
    .Y(_08634_));
 sky130_fd_sc_hd__o21ai_0 _28011_ (.A1(net2785),
    .A2(\inst$top.soc.cpu.gprf.mem[26][20] ),
    .B1(net2734),
    .Y(_08635_));
 sky130_fd_sc_hd__nor2_1 _28012_ (.A(net2789),
    .B(\inst$top.soc.cpu.gprf.mem[24][20] ),
    .Y(_08636_));
 sky130_fd_sc_hd__o21ai_0 _28013_ (.A1(\inst$top.soc.cpu.gprf.mem[25][20] ),
    .A2(net2383),
    .B1(net2331),
    .Y(_08637_));
 sky130_fd_sc_hd__o22ai_1 _28014_ (.A1(_08634_),
    .A2(_08635_),
    .B1(_08636_),
    .B2(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__nor2_1 _28015_ (.A(net2708),
    .B(_08638_),
    .Y(_08639_));
 sky130_fd_sc_hd__nor2_1 _28016_ (.A(net2436),
    .B(_08639_),
    .Y(_08640_));
 sky130_fd_sc_hd__o21ai_0 _28017_ (.A1(net2422),
    .A2(_08633_),
    .B1(_08640_),
    .Y(_08641_));
 sky130_fd_sc_hd__nor2_1 _28018_ (.A(\inst$top.soc.cpu.gprf.mem[23][20] ),
    .B(net2385),
    .Y(_08642_));
 sky130_fd_sc_hd__o21ai_0 _28019_ (.A1(net2789),
    .A2(\inst$top.soc.cpu.gprf.mem[22][20] ),
    .B1(net2734),
    .Y(_08643_));
 sky130_fd_sc_hd__nor2_1 _28020_ (.A(net2789),
    .B(\inst$top.soc.cpu.gprf.mem[20][20] ),
    .Y(_08644_));
 sky130_fd_sc_hd__o21ai_0 _28021_ (.A1(\inst$top.soc.cpu.gprf.mem[21][20] ),
    .A2(net2383),
    .B1(net2331),
    .Y(_08645_));
 sky130_fd_sc_hd__o221ai_1 _28022_ (.A1(_08642_),
    .A2(_08643_),
    .B1(_08644_),
    .B2(_08645_),
    .C1(net2709),
    .Y(_08646_));
 sky130_fd_sc_hd__nor2_1 _28023_ (.A(\inst$top.soc.cpu.gprf.mem[19][20] ),
    .B(net2379),
    .Y(_08647_));
 sky130_fd_sc_hd__o21ai_0 _28024_ (.A1(net2782),
    .A2(\inst$top.soc.cpu.gprf.mem[18][20] ),
    .B1(net2732),
    .Y(_08648_));
 sky130_fd_sc_hd__nor2_1 _28025_ (.A(net2782),
    .B(\inst$top.soc.cpu.gprf.mem[16][20] ),
    .Y(_08649_));
 sky130_fd_sc_hd__o21ai_0 _28026_ (.A1(\inst$top.soc.cpu.gprf.mem[17][20] ),
    .A2(net2379),
    .B1(net2330),
    .Y(_08650_));
 sky130_fd_sc_hd__o221ai_1 _28027_ (.A1(_08647_),
    .A2(_08648_),
    .B1(_08649_),
    .B2(_08650_),
    .C1(net2421),
    .Y(_08651_));
 sky130_fd_sc_hd__nand3_1 _28028_ (.A(_08646_),
    .B(_08651_),
    .C(net2436),
    .Y(_08652_));
 sky130_fd_sc_hd__nor2_1 _28029_ (.A(\inst$top.soc.cpu.gprf.mem[7][20] ),
    .B(net2385),
    .Y(_08653_));
 sky130_fd_sc_hd__o21ai_0 _28030_ (.A1(net2789),
    .A2(\inst$top.soc.cpu.gprf.mem[6][20] ),
    .B1(net2734),
    .Y(_08654_));
 sky130_fd_sc_hd__nor2_1 _28031_ (.A(net2789),
    .B(\inst$top.soc.cpu.gprf.mem[4][20] ),
    .Y(_08655_));
 sky130_fd_sc_hd__o21ai_0 _28032_ (.A1(\inst$top.soc.cpu.gprf.mem[5][20] ),
    .A2(net2385),
    .B1(net2331),
    .Y(_08656_));
 sky130_fd_sc_hd__o221ai_1 _28033_ (.A1(_08653_),
    .A2(_08654_),
    .B1(_08655_),
    .B2(_08656_),
    .C1(net2708),
    .Y(_08657_));
 sky130_fd_sc_hd__nor2_1 _28034_ (.A(\inst$top.soc.cpu.gprf.mem[3][20] ),
    .B(net2379),
    .Y(_08658_));
 sky130_fd_sc_hd__o21ai_0 _28035_ (.A1(net2789),
    .A2(\inst$top.soc.cpu.gprf.mem[2][20] ),
    .B1(net2734),
    .Y(_08659_));
 sky130_fd_sc_hd__nor2_1 _28037_ (.A(net2789),
    .B(\inst$top.soc.cpu.gprf.mem[0][20] ),
    .Y(_08661_));
 sky130_fd_sc_hd__o21ai_0 _28038_ (.A1(\inst$top.soc.cpu.gprf.mem[1][20] ),
    .A2(net2385),
    .B1(net2331),
    .Y(_08662_));
 sky130_fd_sc_hd__o221ai_1 _28039_ (.A1(_08658_),
    .A2(_08659_),
    .B1(_08661_),
    .B2(_08662_),
    .C1(net2422),
    .Y(_08663_));
 sky130_fd_sc_hd__a31oi_1 _28040_ (.A1(_08657_),
    .A2(_08663_),
    .A3(net2435),
    .B1(net2694),
    .Y(_08664_));
 sky130_fd_sc_hd__nor2_1 _28041_ (.A(\inst$top.soc.cpu.gprf.mem[15][20] ),
    .B(net2383),
    .Y(_08665_));
 sky130_fd_sc_hd__o21ai_0 _28042_ (.A1(net2789),
    .A2(\inst$top.soc.cpu.gprf.mem[14][20] ),
    .B1(net2734),
    .Y(_08666_));
 sky130_fd_sc_hd__nor2_1 _28043_ (.A(net2789),
    .B(\inst$top.soc.cpu.gprf.mem[12][20] ),
    .Y(_08667_));
 sky130_fd_sc_hd__o21ai_0 _28044_ (.A1(\inst$top.soc.cpu.gprf.mem[13][20] ),
    .A2(net2383),
    .B1(net2331),
    .Y(_08668_));
 sky130_fd_sc_hd__o221ai_1 _28045_ (.A1(_08665_),
    .A2(_08666_),
    .B1(_08667_),
    .B2(_08668_),
    .C1(net2708),
    .Y(_08669_));
 sky130_fd_sc_hd__nor2_1 _28046_ (.A(\inst$top.soc.cpu.gprf.mem[11][20] ),
    .B(net2379),
    .Y(_08670_));
 sky130_fd_sc_hd__o21ai_0 _28047_ (.A1(net2782),
    .A2(\inst$top.soc.cpu.gprf.mem[10][20] ),
    .B1(net2732),
    .Y(_08671_));
 sky130_fd_sc_hd__nor2_1 _28048_ (.A(net2782),
    .B(\inst$top.soc.cpu.gprf.mem[8][20] ),
    .Y(_08672_));
 sky130_fd_sc_hd__o21ai_0 _28049_ (.A1(\inst$top.soc.cpu.gprf.mem[9][20] ),
    .A2(net2379),
    .B1(net2330),
    .Y(_08673_));
 sky130_fd_sc_hd__o221ai_1 _28050_ (.A1(_08670_),
    .A2(_08671_),
    .B1(_08672_),
    .B2(_08673_),
    .C1(net2421),
    .Y(_08674_));
 sky130_fd_sc_hd__nand3_1 _28051_ (.A(_08669_),
    .B(_08674_),
    .C(net2699),
    .Y(_08675_));
 sky130_fd_sc_hd__a32oi_1 _28052_ (.A1(net2694),
    .A2(_08641_),
    .A3(_08652_),
    .B1(_08664_),
    .B2(_08675_),
    .Y(_00044_));
 sky130_fd_sc_hd__nor2_1 _28053_ (.A(\inst$top.soc.cpu.gprf.mem[31][21] ),
    .B(net2399),
    .Y(_08676_));
 sky130_fd_sc_hd__o21ai_0 _28054_ (.A1(net2806),
    .A2(\inst$top.soc.cpu.gprf.mem[30][21] ),
    .B1(net2743),
    .Y(_08677_));
 sky130_fd_sc_hd__nor2_1 _28055_ (.A(net2806),
    .B(\inst$top.soc.cpu.gprf.mem[28][21] ),
    .Y(_08678_));
 sky130_fd_sc_hd__o21ai_0 _28056_ (.A1(\inst$top.soc.cpu.gprf.mem[29][21] ),
    .A2(net2399),
    .B1(net2340),
    .Y(_08679_));
 sky130_fd_sc_hd__o22ai_1 _28057_ (.A1(_08676_),
    .A2(_08677_),
    .B1(_08678_),
    .B2(_08679_),
    .Y(_08680_));
 sky130_fd_sc_hd__nor2_1 _28058_ (.A(\inst$top.soc.cpu.gprf.mem[27][21] ),
    .B(net2404),
    .Y(_08681_));
 sky130_fd_sc_hd__o21ai_0 _28059_ (.A1(net2811),
    .A2(\inst$top.soc.cpu.gprf.mem[26][21] ),
    .B1(net2746),
    .Y(_08682_));
 sky130_fd_sc_hd__nor2_1 _28060_ (.A(net2811),
    .B(\inst$top.soc.cpu.gprf.mem[24][21] ),
    .Y(_08683_));
 sky130_fd_sc_hd__o21ai_0 _28061_ (.A1(\inst$top.soc.cpu.gprf.mem[25][21] ),
    .A2(net2399),
    .B1(net2343),
    .Y(_08684_));
 sky130_fd_sc_hd__o22ai_1 _28062_ (.A1(_08681_),
    .A2(_08682_),
    .B1(_08683_),
    .B2(_08684_),
    .Y(_08685_));
 sky130_fd_sc_hd__nor2_1 _28063_ (.A(net2714),
    .B(_08685_),
    .Y(_08686_));
 sky130_fd_sc_hd__nor2_1 _28064_ (.A(net2439),
    .B(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__o21ai_0 _28065_ (.A1(net2426),
    .A2(_08680_),
    .B1(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__nor2_1 _28066_ (.A(\inst$top.soc.cpu.gprf.mem[23][21] ),
    .B(net2398),
    .Y(_08689_));
 sky130_fd_sc_hd__o21ai_0 _28067_ (.A1(net2805),
    .A2(\inst$top.soc.cpu.gprf.mem[22][21] ),
    .B1(net2743),
    .Y(_08690_));
 sky130_fd_sc_hd__nor2_1 _28068_ (.A(net2806),
    .B(\inst$top.soc.cpu.gprf.mem[20][21] ),
    .Y(_08691_));
 sky130_fd_sc_hd__o21ai_0 _28069_ (.A1(\inst$top.soc.cpu.gprf.mem[21][21] ),
    .A2(net2398),
    .B1(net2340),
    .Y(_08692_));
 sky130_fd_sc_hd__o221ai_1 _28070_ (.A1(_08689_),
    .A2(_08690_),
    .B1(_08691_),
    .B2(_08692_),
    .C1(net2713),
    .Y(_08693_));
 sky130_fd_sc_hd__nor2_1 _28071_ (.A(\inst$top.soc.cpu.gprf.mem[19][21] ),
    .B(net2398),
    .Y(_08694_));
 sky130_fd_sc_hd__o21ai_0 _28072_ (.A1(net2805),
    .A2(\inst$top.soc.cpu.gprf.mem[18][21] ),
    .B1(net2743),
    .Y(_08695_));
 sky130_fd_sc_hd__nor2_1 _28073_ (.A(net2805),
    .B(\inst$top.soc.cpu.gprf.mem[16][21] ),
    .Y(_08696_));
 sky130_fd_sc_hd__o21ai_0 _28074_ (.A1(\inst$top.soc.cpu.gprf.mem[17][21] ),
    .A2(net2399),
    .B1(net2340),
    .Y(_08697_));
 sky130_fd_sc_hd__o221ai_1 _28075_ (.A1(_08694_),
    .A2(_08695_),
    .B1(_08696_),
    .B2(_08697_),
    .C1(net2426),
    .Y(_08698_));
 sky130_fd_sc_hd__nand3_1 _28076_ (.A(_08693_),
    .B(_08698_),
    .C(net2439),
    .Y(_08699_));
 sky130_fd_sc_hd__nor2_1 _28077_ (.A(\inst$top.soc.cpu.gprf.mem[11][21] ),
    .B(net2403),
    .Y(_08700_));
 sky130_fd_sc_hd__o21ai_0 _28078_ (.A1(net2806),
    .A2(\inst$top.soc.cpu.gprf.mem[10][21] ),
    .B1(net2743),
    .Y(_08701_));
 sky130_fd_sc_hd__nor2_1 _28079_ (.A(net2807),
    .B(\inst$top.soc.cpu.gprf.mem[8][21] ),
    .Y(_08702_));
 sky130_fd_sc_hd__o21ai_0 _28080_ (.A1(\inst$top.soc.cpu.gprf.mem[9][21] ),
    .A2(net2403),
    .B1(net2342),
    .Y(_08703_));
 sky130_fd_sc_hd__o221ai_1 _28081_ (.A1(_08700_),
    .A2(_08701_),
    .B1(_08702_),
    .B2(_08703_),
    .C1(net2426),
    .Y(_08704_));
 sky130_fd_sc_hd__nor2_1 _28082_ (.A(\inst$top.soc.cpu.gprf.mem[15][21] ),
    .B(net2403),
    .Y(_08705_));
 sky130_fd_sc_hd__o21ai_0 _28083_ (.A1(net2806),
    .A2(\inst$top.soc.cpu.gprf.mem[14][21] ),
    .B1(net2743),
    .Y(_08706_));
 sky130_fd_sc_hd__nor2_1 _28084_ (.A(net2807),
    .B(\inst$top.soc.cpu.gprf.mem[12][21] ),
    .Y(_08707_));
 sky130_fd_sc_hd__o21ai_0 _28085_ (.A1(\inst$top.soc.cpu.gprf.mem[13][21] ),
    .A2(net2399),
    .B1(net2340),
    .Y(_08708_));
 sky130_fd_sc_hd__o221ai_1 _28086_ (.A1(_08705_),
    .A2(_08706_),
    .B1(_08707_),
    .B2(_08708_),
    .C1(net2713),
    .Y(_08709_));
 sky130_fd_sc_hd__a31oi_1 _28087_ (.A1(_08704_),
    .A2(_08709_),
    .A3(net2699),
    .B1(net2693),
    .Y(_08710_));
 sky130_fd_sc_hd__nor2_1 _28088_ (.A(\inst$top.soc.cpu.gprf.mem[7][21] ),
    .B(net2398),
    .Y(_08711_));
 sky130_fd_sc_hd__o21ai_0 _28089_ (.A1(net2806),
    .A2(\inst$top.soc.cpu.gprf.mem[6][21] ),
    .B1(net2745),
    .Y(_08712_));
 sky130_fd_sc_hd__nor2_1 _28090_ (.A(net2807),
    .B(\inst$top.soc.cpu.gprf.mem[4][21] ),
    .Y(_08713_));
 sky130_fd_sc_hd__o21ai_0 _28091_ (.A1(\inst$top.soc.cpu.gprf.mem[5][21] ),
    .A2(net2399),
    .B1(net2340),
    .Y(_08714_));
 sky130_fd_sc_hd__o221ai_1 _28092_ (.A1(_08711_),
    .A2(_08712_),
    .B1(_08713_),
    .B2(_08714_),
    .C1(net2713),
    .Y(_08715_));
 sky130_fd_sc_hd__nor2_1 _28093_ (.A(\inst$top.soc.cpu.gprf.mem[3][21] ),
    .B(net2398),
    .Y(_08716_));
 sky130_fd_sc_hd__o21ai_0 _28094_ (.A1(net2806),
    .A2(\inst$top.soc.cpu.gprf.mem[2][21] ),
    .B1(net2743),
    .Y(_08717_));
 sky130_fd_sc_hd__nor2_1 _28095_ (.A(net2806),
    .B(\inst$top.soc.cpu.gprf.mem[0][21] ),
    .Y(_08718_));
 sky130_fd_sc_hd__o21ai_0 _28096_ (.A1(\inst$top.soc.cpu.gprf.mem[1][21] ),
    .A2(net2399),
    .B1(net2340),
    .Y(_08719_));
 sky130_fd_sc_hd__o221ai_1 _28097_ (.A1(_08716_),
    .A2(_08717_),
    .B1(_08718_),
    .B2(_08719_),
    .C1(net2426),
    .Y(_08720_));
 sky130_fd_sc_hd__nand3_1 _28098_ (.A(_08715_),
    .B(_08720_),
    .C(net2439),
    .Y(_08721_));
 sky130_fd_sc_hd__a32oi_1 _28099_ (.A1(net2693),
    .A2(_08688_),
    .A3(_08699_),
    .B1(_08710_),
    .B2(_08721_),
    .Y(_00045_));
 sky130_fd_sc_hd__nor2_1 _28100_ (.A(\inst$top.soc.cpu.gprf.mem[7][22] ),
    .B(net2362),
    .Y(_08722_));
 sky130_fd_sc_hd__o21ai_0 _28101_ (.A1(net2763),
    .A2(\inst$top.soc.cpu.gprf.mem[6][22] ),
    .B1(net2722),
    .Y(_08723_));
 sky130_fd_sc_hd__nor2_1 _28102_ (.A(net2763),
    .B(\inst$top.soc.cpu.gprf.mem[4][22] ),
    .Y(_08724_));
 sky130_fd_sc_hd__o21ai_0 _28103_ (.A1(\inst$top.soc.cpu.gprf.mem[5][22] ),
    .A2(net2362),
    .B1(net2319),
    .Y(_08725_));
 sky130_fd_sc_hd__o221ai_1 _28104_ (.A1(_08722_),
    .A2(_08723_),
    .B1(_08724_),
    .B2(_08725_),
    .C1(net2702),
    .Y(_08726_));
 sky130_fd_sc_hd__nor2_1 _28105_ (.A(\inst$top.soc.cpu.gprf.mem[3][22] ),
    .B(net2362),
    .Y(_08727_));
 sky130_fd_sc_hd__o21ai_0 _28106_ (.A1(net2765),
    .A2(\inst$top.soc.cpu.gprf.mem[2][22] ),
    .B1(net2722),
    .Y(_08728_));
 sky130_fd_sc_hd__nor2_1 _28107_ (.A(net2763),
    .B(\inst$top.soc.cpu.gprf.mem[0][22] ),
    .Y(_08729_));
 sky130_fd_sc_hd__o21ai_0 _28108_ (.A1(\inst$top.soc.cpu.gprf.mem[1][22] ),
    .A2(net2362),
    .B1(net2319),
    .Y(_08730_));
 sky130_fd_sc_hd__o221ai_1 _28109_ (.A1(_08727_),
    .A2(_08728_),
    .B1(_08729_),
    .B2(_08730_),
    .C1(net2415),
    .Y(_08731_));
 sky130_fd_sc_hd__nand3_1 _28110_ (.A(_08726_),
    .B(_08731_),
    .C(net2431),
    .Y(_08732_));
 sky130_fd_sc_hd__nor2_1 _28111_ (.A(\inst$top.soc.cpu.gprf.mem[11][22] ),
    .B(net2364),
    .Y(_08733_));
 sky130_fd_sc_hd__o21ai_0 _28112_ (.A1(net2763),
    .A2(\inst$top.soc.cpu.gprf.mem[10][22] ),
    .B1(net2722),
    .Y(_08734_));
 sky130_fd_sc_hd__nor2_1 _28113_ (.A(net2763),
    .B(\inst$top.soc.cpu.gprf.mem[8][22] ),
    .Y(_08735_));
 sky130_fd_sc_hd__o21ai_0 _28114_ (.A1(\inst$top.soc.cpu.gprf.mem[9][22] ),
    .A2(net2364),
    .B1(net2321),
    .Y(_08736_));
 sky130_fd_sc_hd__o221ai_1 _28115_ (.A1(_08733_),
    .A2(_08734_),
    .B1(_08735_),
    .B2(_08736_),
    .C1(net2415),
    .Y(_08737_));
 sky130_fd_sc_hd__nor2_1 _28116_ (.A(\inst$top.soc.cpu.gprf.mem[15][22] ),
    .B(net2364),
    .Y(_08738_));
 sky130_fd_sc_hd__o21ai_0 _28117_ (.A1(net2765),
    .A2(\inst$top.soc.cpu.gprf.mem[14][22] ),
    .B1(net2722),
    .Y(_08739_));
 sky130_fd_sc_hd__nor2_1 _28118_ (.A(net2763),
    .B(\inst$top.soc.cpu.gprf.mem[12][22] ),
    .Y(_08740_));
 sky130_fd_sc_hd__o21ai_0 _28119_ (.A1(\inst$top.soc.cpu.gprf.mem[13][22] ),
    .A2(net2364),
    .B1(net2321),
    .Y(_08741_));
 sky130_fd_sc_hd__o221ai_1 _28120_ (.A1(_08738_),
    .A2(_08739_),
    .B1(_08740_),
    .B2(_08741_),
    .C1(net2702),
    .Y(_08742_));
 sky130_fd_sc_hd__nand3_1 _28121_ (.A(_08737_),
    .B(_08742_),
    .C(net2696),
    .Y(_08743_));
 sky130_fd_sc_hd__nor2_1 _28122_ (.A(\inst$top.soc.cpu.gprf.mem[31][22] ),
    .B(net2362),
    .Y(_08744_));
 sky130_fd_sc_hd__o21ai_0 _28123_ (.A1(net2764),
    .A2(\inst$top.soc.cpu.gprf.mem[30][22] ),
    .B1(net2722),
    .Y(_08745_));
 sky130_fd_sc_hd__nor2_1 _28124_ (.A(net2764),
    .B(\inst$top.soc.cpu.gprf.mem[28][22] ),
    .Y(_08746_));
 sky130_fd_sc_hd__o21ai_0 _28125_ (.A1(\inst$top.soc.cpu.gprf.mem[29][22] ),
    .A2(net2362),
    .B1(net2319),
    .Y(_08747_));
 sky130_fd_sc_hd__o221ai_1 _28126_ (.A1(_08744_),
    .A2(_08745_),
    .B1(_08746_),
    .B2(_08747_),
    .C1(net2702),
    .Y(_08748_));
 sky130_fd_sc_hd__nor2_1 _28127_ (.A(\inst$top.soc.cpu.gprf.mem[27][22] ),
    .B(net2362),
    .Y(_08749_));
 sky130_fd_sc_hd__o21ai_0 _28128_ (.A1(net2763),
    .A2(\inst$top.soc.cpu.gprf.mem[26][22] ),
    .B1(net2722),
    .Y(_08750_));
 sky130_fd_sc_hd__nor2_1 _28129_ (.A(net2763),
    .B(\inst$top.soc.cpu.gprf.mem[24][22] ),
    .Y(_08751_));
 sky130_fd_sc_hd__o21ai_0 _28130_ (.A1(\inst$top.soc.cpu.gprf.mem[25][22] ),
    .A2(net2362),
    .B1(net2319),
    .Y(_08752_));
 sky130_fd_sc_hd__o221ai_1 _28131_ (.A1(_08749_),
    .A2(_08750_),
    .B1(_08751_),
    .B2(_08752_),
    .C1(net2415),
    .Y(_08753_));
 sky130_fd_sc_hd__a31oi_1 _28132_ (.A1(_08748_),
    .A2(_08753_),
    .A3(net2696),
    .B1(net2445),
    .Y(_08754_));
 sky130_fd_sc_hd__nor2_1 _28133_ (.A(\inst$top.soc.cpu.gprf.mem[23][22] ),
    .B(net2361),
    .Y(_08755_));
 sky130_fd_sc_hd__o21ai_0 _28134_ (.A1(net2764),
    .A2(\inst$top.soc.cpu.gprf.mem[22][22] ),
    .B1(net2723),
    .Y(_08756_));
 sky130_fd_sc_hd__nor2_1 _28135_ (.A(net2764),
    .B(\inst$top.soc.cpu.gprf.mem[20][22] ),
    .Y(_08757_));
 sky130_fd_sc_hd__o21ai_0 _28136_ (.A1(\inst$top.soc.cpu.gprf.mem[21][22] ),
    .A2(net2361),
    .B1(net2319),
    .Y(_08758_));
 sky130_fd_sc_hd__o221ai_1 _28137_ (.A1(_08755_),
    .A2(_08756_),
    .B1(_08757_),
    .B2(_08758_),
    .C1(net2702),
    .Y(_08759_));
 sky130_fd_sc_hd__nor2_1 _28138_ (.A(\inst$top.soc.cpu.gprf.mem[19][22] ),
    .B(net2363),
    .Y(_08760_));
 sky130_fd_sc_hd__o21ai_0 _28139_ (.A1(net2765),
    .A2(\inst$top.soc.cpu.gprf.mem[18][22] ),
    .B1(net2722),
    .Y(_08761_));
 sky130_fd_sc_hd__nor2_1 _28140_ (.A(net2764),
    .B(\inst$top.soc.cpu.gprf.mem[16][22] ),
    .Y(_08762_));
 sky130_fd_sc_hd__o21ai_0 _28141_ (.A1(\inst$top.soc.cpu.gprf.mem[17][22] ),
    .A2(net2361),
    .B1(net2320),
    .Y(_08763_));
 sky130_fd_sc_hd__o221ai_1 _28142_ (.A1(_08760_),
    .A2(_08761_),
    .B1(_08762_),
    .B2(_08763_),
    .C1(net2416),
    .Y(_08764_));
 sky130_fd_sc_hd__nand3_1 _28143_ (.A(_08759_),
    .B(_08764_),
    .C(net2431),
    .Y(_08765_));
 sky130_fd_sc_hd__a32oi_1 _28144_ (.A1(_08732_),
    .A2(_08743_),
    .A3(net2445),
    .B1(_08754_),
    .B2(_08765_),
    .Y(_00046_));
 sky130_fd_sc_hd__nor2_1 _28145_ (.A(\inst$top.soc.cpu.gprf.mem[15][23] ),
    .B(net2378),
    .Y(_08766_));
 sky130_fd_sc_hd__o21ai_0 _28146_ (.A1(net2783),
    .A2(\inst$top.soc.cpu.gprf.mem[14][23] ),
    .B1(net2732),
    .Y(_08767_));
 sky130_fd_sc_hd__nor2_1 _28147_ (.A(net2783),
    .B(\inst$top.soc.cpu.gprf.mem[12][23] ),
    .Y(_08768_));
 sky130_fd_sc_hd__o21ai_0 _28148_ (.A1(\inst$top.soc.cpu.gprf.mem[13][23] ),
    .A2(net2378),
    .B1(net2330),
    .Y(_08769_));
 sky130_fd_sc_hd__o221ai_1 _28149_ (.A1(_08766_),
    .A2(_08767_),
    .B1(_08768_),
    .B2(_08769_),
    .C1(net2707),
    .Y(_08770_));
 sky130_fd_sc_hd__nor2_1 _28150_ (.A(\inst$top.soc.cpu.gprf.mem[11][23] ),
    .B(net2378),
    .Y(_08771_));
 sky130_fd_sc_hd__o21ai_0 _28151_ (.A1(net2782),
    .A2(\inst$top.soc.cpu.gprf.mem[10][23] ),
    .B1(net2732),
    .Y(_08772_));
 sky130_fd_sc_hd__nor2_1 _28152_ (.A(net2782),
    .B(\inst$top.soc.cpu.gprf.mem[8][23] ),
    .Y(_08773_));
 sky130_fd_sc_hd__o21ai_0 _28153_ (.A1(\inst$top.soc.cpu.gprf.mem[9][23] ),
    .A2(net2378),
    .B1(net2330),
    .Y(_08774_));
 sky130_fd_sc_hd__o221ai_1 _28154_ (.A1(_08771_),
    .A2(_08772_),
    .B1(_08773_),
    .B2(_08774_),
    .C1(net2421),
    .Y(_08775_));
 sky130_fd_sc_hd__nand3_1 _28155_ (.A(_08770_),
    .B(_08775_),
    .C(net2699),
    .Y(_08776_));
 sky130_fd_sc_hd__nor2_1 _28156_ (.A(\inst$top.soc.cpu.gprf.mem[7][23] ),
    .B(net2379),
    .Y(_08777_));
 sky130_fd_sc_hd__o21ai_0 _28157_ (.A1(net2782),
    .A2(\inst$top.soc.cpu.gprf.mem[6][23] ),
    .B1(net2732),
    .Y(_08778_));
 sky130_fd_sc_hd__nor2_1 _28158_ (.A(net2782),
    .B(\inst$top.soc.cpu.gprf.mem[4][23] ),
    .Y(_08779_));
 sky130_fd_sc_hd__o21ai_0 _28159_ (.A1(\inst$top.soc.cpu.gprf.mem[5][23] ),
    .A2(net2379),
    .B1(net2330),
    .Y(_08780_));
 sky130_fd_sc_hd__o221ai_1 _28160_ (.A1(_08777_),
    .A2(_08778_),
    .B1(_08779_),
    .B2(_08780_),
    .C1(net2707),
    .Y(_08781_));
 sky130_fd_sc_hd__nor2_1 _28161_ (.A(\inst$top.soc.cpu.gprf.mem[3][23] ),
    .B(net2378),
    .Y(_08782_));
 sky130_fd_sc_hd__o21ai_0 _28162_ (.A1(net2783),
    .A2(\inst$top.soc.cpu.gprf.mem[2][23] ),
    .B1(net2732),
    .Y(_08783_));
 sky130_fd_sc_hd__nor2_1 _28163_ (.A(net2783),
    .B(\inst$top.soc.cpu.gprf.mem[0][23] ),
    .Y(_08784_));
 sky130_fd_sc_hd__o21ai_0 _28164_ (.A1(\inst$top.soc.cpu.gprf.mem[1][23] ),
    .A2(net2378),
    .B1(net2330),
    .Y(_08785_));
 sky130_fd_sc_hd__o221ai_1 _28165_ (.A1(_08782_),
    .A2(_08783_),
    .B1(_08784_),
    .B2(_08785_),
    .C1(net2421),
    .Y(_08786_));
 sky130_fd_sc_hd__nand3_1 _28166_ (.A(_08781_),
    .B(_08786_),
    .C(net2435),
    .Y(_08787_));
 sky130_fd_sc_hd__nor2_1 _28167_ (.A(\inst$top.soc.cpu.gprf.mem[31][23] ),
    .B(net2379),
    .Y(_08788_));
 sky130_fd_sc_hd__o21ai_0 _28168_ (.A1(net2784),
    .A2(\inst$top.soc.cpu.gprf.mem[30][23] ),
    .B1(net2733),
    .Y(_08789_));
 sky130_fd_sc_hd__nor2_1 _28169_ (.A(net2784),
    .B(\inst$top.soc.cpu.gprf.mem[28][23] ),
    .Y(_08790_));
 sky130_fd_sc_hd__o21ai_0 _28170_ (.A1(\inst$top.soc.cpu.gprf.mem[29][23] ),
    .A2(net2380),
    .B1(net2329),
    .Y(_08791_));
 sky130_fd_sc_hd__o221ai_1 _28171_ (.A1(_08788_),
    .A2(_08789_),
    .B1(_08790_),
    .B2(_08791_),
    .C1(net2707),
    .Y(_08792_));
 sky130_fd_sc_hd__nor2_1 _28172_ (.A(\inst$top.soc.cpu.gprf.mem[27][23] ),
    .B(net2377),
    .Y(_08793_));
 sky130_fd_sc_hd__o21ai_0 _28173_ (.A1(net2781),
    .A2(\inst$top.soc.cpu.gprf.mem[26][23] ),
    .B1(net2732),
    .Y(_08794_));
 sky130_fd_sc_hd__nor2_1 _28174_ (.A(net2781),
    .B(\inst$top.soc.cpu.gprf.mem[24][23] ),
    .Y(_08795_));
 sky130_fd_sc_hd__o21ai_0 _28175_ (.A1(\inst$top.soc.cpu.gprf.mem[25][23] ),
    .A2(net2377),
    .B1(net2329),
    .Y(_08796_));
 sky130_fd_sc_hd__o221ai_1 _28176_ (.A1(_08793_),
    .A2(_08794_),
    .B1(_08795_),
    .B2(_08796_),
    .C1(net2421),
    .Y(_08797_));
 sky130_fd_sc_hd__a31oi_1 _28177_ (.A1(_08792_),
    .A2(_08797_),
    .A3(net2699),
    .B1(net2442),
    .Y(_08798_));
 sky130_fd_sc_hd__nor2_1 _28178_ (.A(\inst$top.soc.cpu.gprf.mem[23][23] ),
    .B(net2378),
    .Y(_08799_));
 sky130_fd_sc_hd__o21ai_0 _28179_ (.A1(net2782),
    .A2(\inst$top.soc.cpu.gprf.mem[22][23] ),
    .B1(net2733),
    .Y(_08800_));
 sky130_fd_sc_hd__nor2_1 _28180_ (.A(net2784),
    .B(\inst$top.soc.cpu.gprf.mem[20][23] ),
    .Y(_08801_));
 sky130_fd_sc_hd__o21ai_0 _28181_ (.A1(\inst$top.soc.cpu.gprf.mem[21][23] ),
    .A2(net2378),
    .B1(net2330),
    .Y(_08802_));
 sky130_fd_sc_hd__o221ai_1 _28182_ (.A1(_08799_),
    .A2(_08800_),
    .B1(_08801_),
    .B2(_08802_),
    .C1(net2707),
    .Y(_08803_));
 sky130_fd_sc_hd__nor2_1 _28183_ (.A(\inst$top.soc.cpu.gprf.mem[19][23] ),
    .B(net2378),
    .Y(_08804_));
 sky130_fd_sc_hd__o21ai_0 _28184_ (.A1(net2783),
    .A2(\inst$top.soc.cpu.gprf.mem[18][23] ),
    .B1(net2732),
    .Y(_08805_));
 sky130_fd_sc_hd__nor2_1 _28185_ (.A(net2783),
    .B(\inst$top.soc.cpu.gprf.mem[16][23] ),
    .Y(_08806_));
 sky130_fd_sc_hd__o21ai_0 _28186_ (.A1(\inst$top.soc.cpu.gprf.mem[17][23] ),
    .A2(net2378),
    .B1(net2330),
    .Y(_08807_));
 sky130_fd_sc_hd__o221ai_1 _28187_ (.A1(_08804_),
    .A2(_08805_),
    .B1(_08806_),
    .B2(_08807_),
    .C1(net2421),
    .Y(_08808_));
 sky130_fd_sc_hd__nand3_1 _28188_ (.A(_08803_),
    .B(_08808_),
    .C(net2435),
    .Y(_08809_));
 sky130_fd_sc_hd__a32oi_1 _28189_ (.A1(_08776_),
    .A2(_08787_),
    .A3(net2442),
    .B1(_08798_),
    .B2(_08809_),
    .Y(_00047_));
 sky130_fd_sc_hd__nor2_1 _28190_ (.A(\inst$top.soc.cpu.gprf.mem[11][24] ),
    .B(net2410),
    .Y(_08810_));
 sky130_fd_sc_hd__o21ai_0 _28191_ (.A1(net2816),
    .A2(\inst$top.soc.cpu.gprf.mem[10][24] ),
    .B1(net2749),
    .Y(_08811_));
 sky130_fd_sc_hd__nor2_1 _28192_ (.A(net2817),
    .B(\inst$top.soc.cpu.gprf.mem[8][24] ),
    .Y(_08812_));
 sky130_fd_sc_hd__o21ai_0 _28193_ (.A1(\inst$top.soc.cpu.gprf.mem[9][24] ),
    .A2(net2409),
    .B1(net2345),
    .Y(_08813_));
 sky130_fd_sc_hd__o22ai_1 _28194_ (.A1(_08810_),
    .A2(_08811_),
    .B1(_08812_),
    .B2(_08813_),
    .Y(_08814_));
 sky130_fd_sc_hd__nor2_1 _28195_ (.A(\inst$top.soc.cpu.gprf.mem[15][24] ),
    .B(net2409),
    .Y(_08815_));
 sky130_fd_sc_hd__o21ai_0 _28196_ (.A1(net2816),
    .A2(\inst$top.soc.cpu.gprf.mem[14][24] ),
    .B1(net2748),
    .Y(_08816_));
 sky130_fd_sc_hd__nor2_1 _28197_ (.A(net2816),
    .B(\inst$top.soc.cpu.gprf.mem[12][24] ),
    .Y(_08817_));
 sky130_fd_sc_hd__o21ai_0 _28198_ (.A1(\inst$top.soc.cpu.gprf.mem[13][24] ),
    .A2(net2409),
    .B1(net2344),
    .Y(_08818_));
 sky130_fd_sc_hd__o22ai_1 _28199_ (.A1(_08815_),
    .A2(_08816_),
    .B1(_08817_),
    .B2(_08818_),
    .Y(_08819_));
 sky130_fd_sc_hd__nor2_1 _28200_ (.A(net2428),
    .B(_08819_),
    .Y(_08820_));
 sky130_fd_sc_hd__nor2_1 _28201_ (.A(net2440),
    .B(_08820_),
    .Y(_08821_));
 sky130_fd_sc_hd__o21ai_0 _28202_ (.A1(net2714),
    .A2(_08814_),
    .B1(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__nor2_1 _28203_ (.A(\inst$top.soc.cpu.gprf.mem[7][24] ),
    .B(net2402),
    .Y(_08823_));
 sky130_fd_sc_hd__o21ai_0 _28204_ (.A1(net2809),
    .A2(\inst$top.soc.cpu.gprf.mem[6][24] ),
    .B1(net2744),
    .Y(_08824_));
 sky130_fd_sc_hd__nor2_1 _28205_ (.A(net2810),
    .B(\inst$top.soc.cpu.gprf.mem[4][24] ),
    .Y(_08825_));
 sky130_fd_sc_hd__o21ai_0 _28206_ (.A1(\inst$top.soc.cpu.gprf.mem[5][24] ),
    .A2(net2402),
    .B1(net2342),
    .Y(_08826_));
 sky130_fd_sc_hd__o221ai_1 _28207_ (.A1(_08823_),
    .A2(_08824_),
    .B1(_08825_),
    .B2(_08826_),
    .C1(net2713),
    .Y(_08827_));
 sky130_fd_sc_hd__nor2_1 _28208_ (.A(\inst$top.soc.cpu.gprf.mem[3][24] ),
    .B(net2402),
    .Y(_08828_));
 sky130_fd_sc_hd__o21ai_0 _28209_ (.A1(net2810),
    .A2(\inst$top.soc.cpu.gprf.mem[2][24] ),
    .B1(net2744),
    .Y(_08829_));
 sky130_fd_sc_hd__nor2_1 _28210_ (.A(net2809),
    .B(\inst$top.soc.cpu.gprf.mem[0][24] ),
    .Y(_08830_));
 sky130_fd_sc_hd__o21ai_0 _28211_ (.A1(\inst$top.soc.cpu.gprf.mem[1][24] ),
    .A2(net2402),
    .B1(net2342),
    .Y(_08831_));
 sky130_fd_sc_hd__o221ai_1 _28212_ (.A1(_08828_),
    .A2(_08829_),
    .B1(_08830_),
    .B2(_08831_),
    .C1(net2428),
    .Y(_08832_));
 sky130_fd_sc_hd__nand3_1 _28213_ (.A(_08827_),
    .B(_08832_),
    .C(net2439),
    .Y(_08833_));
 sky130_fd_sc_hd__nor2_1 _28214_ (.A(\inst$top.soc.cpu.gprf.mem[31][24] ),
    .B(net2402),
    .Y(_08834_));
 sky130_fd_sc_hd__o21ai_0 _28215_ (.A1(net2809),
    .A2(\inst$top.soc.cpu.gprf.mem[30][24] ),
    .B1(net2745),
    .Y(_08835_));
 sky130_fd_sc_hd__nor2_1 _28216_ (.A(net2809),
    .B(\inst$top.soc.cpu.gprf.mem[28][24] ),
    .Y(_08836_));
 sky130_fd_sc_hd__o21ai_0 _28217_ (.A1(\inst$top.soc.cpu.gprf.mem[29][24] ),
    .A2(net2402),
    .B1(net2341),
    .Y(_08837_));
 sky130_fd_sc_hd__o221ai_1 _28218_ (.A1(_08834_),
    .A2(_08835_),
    .B1(_08836_),
    .B2(_08837_),
    .C1(net2713),
    .Y(_08838_));
 sky130_fd_sc_hd__nor2_1 _28219_ (.A(\inst$top.soc.cpu.gprf.mem[27][24] ),
    .B(net2402),
    .Y(_08839_));
 sky130_fd_sc_hd__o21ai_0 _28220_ (.A1(net2809),
    .A2(\inst$top.soc.cpu.gprf.mem[26][24] ),
    .B1(net2745),
    .Y(_08840_));
 sky130_fd_sc_hd__nor2_1 _28221_ (.A(net2809),
    .B(\inst$top.soc.cpu.gprf.mem[24][24] ),
    .Y(_08841_));
 sky130_fd_sc_hd__o21ai_0 _28222_ (.A1(\inst$top.soc.cpu.gprf.mem[25][24] ),
    .A2(net2402),
    .B1(net2341),
    .Y(_08842_));
 sky130_fd_sc_hd__o221ai_1 _28223_ (.A1(_08839_),
    .A2(_08840_),
    .B1(_08841_),
    .B2(_08842_),
    .C1(net2428),
    .Y(_08843_));
 sky130_fd_sc_hd__a31oi_1 _28224_ (.A1(_08838_),
    .A2(_08843_),
    .A3(net2698),
    .B1(net2443),
    .Y(_08844_));
 sky130_fd_sc_hd__nor2_1 _28225_ (.A(\inst$top.soc.cpu.gprf.mem[23][24] ),
    .B(net2409),
    .Y(_08845_));
 sky130_fd_sc_hd__o21ai_0 _28226_ (.A1(net2816),
    .A2(\inst$top.soc.cpu.gprf.mem[22][24] ),
    .B1(net2749),
    .Y(_08846_));
 sky130_fd_sc_hd__nor2_1 _28227_ (.A(net2817),
    .B(\inst$top.soc.cpu.gprf.mem[20][24] ),
    .Y(_08847_));
 sky130_fd_sc_hd__o21ai_0 _28228_ (.A1(\inst$top.soc.cpu.gprf.mem[21][24] ),
    .A2(net2409),
    .B1(net2344),
    .Y(_08848_));
 sky130_fd_sc_hd__o221ai_1 _28229_ (.A1(_08845_),
    .A2(_08846_),
    .B1(_08847_),
    .B2(_08848_),
    .C1(net2714),
    .Y(_08849_));
 sky130_fd_sc_hd__nor2_1 _28230_ (.A(\inst$top.soc.cpu.gprf.mem[19][24] ),
    .B(net2409),
    .Y(_08850_));
 sky130_fd_sc_hd__o21ai_0 _28231_ (.A1(net2817),
    .A2(\inst$top.soc.cpu.gprf.mem[18][24] ),
    .B1(net2748),
    .Y(_08851_));
 sky130_fd_sc_hd__nor2_1 _28232_ (.A(net2816),
    .B(\inst$top.soc.cpu.gprf.mem[16][24] ),
    .Y(_08852_));
 sky130_fd_sc_hd__o21ai_0 _28233_ (.A1(\inst$top.soc.cpu.gprf.mem[17][24] ),
    .A2(net2409),
    .B1(net2345),
    .Y(_08853_));
 sky130_fd_sc_hd__o221ai_1 _28234_ (.A1(_08850_),
    .A2(_08851_),
    .B1(_08852_),
    .B2(_08853_),
    .C1(net2427),
    .Y(_08854_));
 sky130_fd_sc_hd__nand3_1 _28235_ (.A(_08849_),
    .B(_08854_),
    .C(net2439),
    .Y(_08855_));
 sky130_fd_sc_hd__a32oi_1 _28236_ (.A1(net2443),
    .A2(_08822_),
    .A3(_08833_),
    .B1(_08844_),
    .B2(_08855_),
    .Y(_00048_));
 sky130_fd_sc_hd__nor2_1 _28237_ (.A(\inst$top.soc.cpu.gprf.mem[7][25] ),
    .B(net2369),
    .Y(_08856_));
 sky130_fd_sc_hd__o21ai_0 _28238_ (.A1(net2777),
    .A2(\inst$top.soc.cpu.gprf.mem[6][25] ),
    .B1(net2729),
    .Y(_08857_));
 sky130_fd_sc_hd__nor2_1 _28239_ (.A(net2777),
    .B(\inst$top.soc.cpu.gprf.mem[4][25] ),
    .Y(_08858_));
 sky130_fd_sc_hd__o21ai_0 _28240_ (.A1(\inst$top.soc.cpu.gprf.mem[5][25] ),
    .A2(net2369),
    .B1(net2325),
    .Y(_08859_));
 sky130_fd_sc_hd__o221ai_1 _28241_ (.A1(_08856_),
    .A2(_08857_),
    .B1(_08858_),
    .B2(_08859_),
    .C1(net2705),
    .Y(_08860_));
 sky130_fd_sc_hd__nor2_1 _28242_ (.A(\inst$top.soc.cpu.gprf.mem[3][25] ),
    .B(net2369),
    .Y(_08861_));
 sky130_fd_sc_hd__o21ai_0 _28243_ (.A1(net2772),
    .A2(\inst$top.soc.cpu.gprf.mem[2][25] ),
    .B1(net2726),
    .Y(_08862_));
 sky130_fd_sc_hd__nor2_1 _28244_ (.A(net2772),
    .B(\inst$top.soc.cpu.gprf.mem[0][25] ),
    .Y(_08863_));
 sky130_fd_sc_hd__o21ai_0 _28245_ (.A1(\inst$top.soc.cpu.gprf.mem[1][25] ),
    .A2(net2369),
    .B1(net2325),
    .Y(_08864_));
 sky130_fd_sc_hd__o221ai_1 _28246_ (.A1(_08861_),
    .A2(_08862_),
    .B1(_08863_),
    .B2(_08864_),
    .C1(net2418),
    .Y(_08865_));
 sky130_fd_sc_hd__nand3_1 _28247_ (.A(_08860_),
    .B(_08865_),
    .C(net2433),
    .Y(_08866_));
 sky130_fd_sc_hd__nor2_1 _28248_ (.A(\inst$top.soc.cpu.gprf.mem[11][25] ),
    .B(net2373),
    .Y(_08867_));
 sky130_fd_sc_hd__o21ai_0 _28249_ (.A1(net2777),
    .A2(\inst$top.soc.cpu.gprf.mem[10][25] ),
    .B1(net2729),
    .Y(_08868_));
 sky130_fd_sc_hd__nor2_1 _28250_ (.A(net2777),
    .B(\inst$top.soc.cpu.gprf.mem[8][25] ),
    .Y(_08869_));
 sky130_fd_sc_hd__o21ai_0 _28251_ (.A1(\inst$top.soc.cpu.gprf.mem[9][25] ),
    .A2(net2373),
    .B1(net2327),
    .Y(_08870_));
 sky130_fd_sc_hd__o221ai_1 _28252_ (.A1(_08867_),
    .A2(_08868_),
    .B1(_08869_),
    .B2(_08870_),
    .C1(net2419),
    .Y(_08871_));
 sky130_fd_sc_hd__nor2_1 _28253_ (.A(\inst$top.soc.cpu.gprf.mem[15][25] ),
    .B(net2373),
    .Y(_08872_));
 sky130_fd_sc_hd__o21ai_0 _28254_ (.A1(net2777),
    .A2(\inst$top.soc.cpu.gprf.mem[14][25] ),
    .B1(net2729),
    .Y(_08873_));
 sky130_fd_sc_hd__nor2_1 _28255_ (.A(net2777),
    .B(\inst$top.soc.cpu.gprf.mem[12][25] ),
    .Y(_08874_));
 sky130_fd_sc_hd__o21ai_0 _28256_ (.A1(\inst$top.soc.cpu.gprf.mem[13][25] ),
    .A2(net2373),
    .B1(net2327),
    .Y(_08875_));
 sky130_fd_sc_hd__o221ai_1 _28257_ (.A1(_08872_),
    .A2(_08873_),
    .B1(_08874_),
    .B2(_08875_),
    .C1(net2705),
    .Y(_08876_));
 sky130_fd_sc_hd__nand3_1 _28258_ (.A(_08871_),
    .B(_08876_),
    .C(net2697),
    .Y(_08877_));
 sky130_fd_sc_hd__nor2_1 _28259_ (.A(\inst$top.soc.cpu.gprf.mem[31][25] ),
    .B(net2369),
    .Y(_08878_));
 sky130_fd_sc_hd__o21ai_0 _28260_ (.A1(net2772),
    .A2(\inst$top.soc.cpu.gprf.mem[30][25] ),
    .B1(net2727),
    .Y(_08879_));
 sky130_fd_sc_hd__nor2_1 _28261_ (.A(net2772),
    .B(\inst$top.soc.cpu.gprf.mem[28][25] ),
    .Y(_08880_));
 sky130_fd_sc_hd__o21ai_0 _28262_ (.A1(\inst$top.soc.cpu.gprf.mem[29][25] ),
    .A2(net2369),
    .B1(net2324),
    .Y(_08881_));
 sky130_fd_sc_hd__o221ai_1 _28263_ (.A1(_08878_),
    .A2(_08879_),
    .B1(_08880_),
    .B2(_08881_),
    .C1(net2704),
    .Y(_08882_));
 sky130_fd_sc_hd__nor2_1 _28264_ (.A(\inst$top.soc.cpu.gprf.mem[27][25] ),
    .B(net2369),
    .Y(_08883_));
 sky130_fd_sc_hd__o21ai_0 _28265_ (.A1(net2772),
    .A2(\inst$top.soc.cpu.gprf.mem[26][25] ),
    .B1(net2727),
    .Y(_08884_));
 sky130_fd_sc_hd__nor2_1 _28266_ (.A(net2772),
    .B(\inst$top.soc.cpu.gprf.mem[24][25] ),
    .Y(_08885_));
 sky130_fd_sc_hd__o21ai_0 _28267_ (.A1(\inst$top.soc.cpu.gprf.mem[25][25] ),
    .A2(net2369),
    .B1(net2324),
    .Y(_08886_));
 sky130_fd_sc_hd__o221ai_1 _28268_ (.A1(_08883_),
    .A2(_08884_),
    .B1(_08885_),
    .B2(_08886_),
    .C1(net2418),
    .Y(_08887_));
 sky130_fd_sc_hd__a31oi_1 _28269_ (.A1(_08882_),
    .A2(_08887_),
    .A3(net2697),
    .B1(net2442),
    .Y(_08888_));
 sky130_fd_sc_hd__nor2_1 _28270_ (.A(\inst$top.soc.cpu.gprf.mem[23][25] ),
    .B(net2369),
    .Y(_08889_));
 sky130_fd_sc_hd__o21ai_0 _28271_ (.A1(net2777),
    .A2(\inst$top.soc.cpu.gprf.mem[22][25] ),
    .B1(net2729),
    .Y(_08890_));
 sky130_fd_sc_hd__nor2_1 _28272_ (.A(net2777),
    .B(\inst$top.soc.cpu.gprf.mem[20][25] ),
    .Y(_08891_));
 sky130_fd_sc_hd__o21ai_0 _28273_ (.A1(\inst$top.soc.cpu.gprf.mem[21][25] ),
    .A2(net2369),
    .B1(net2325),
    .Y(_08892_));
 sky130_fd_sc_hd__o221ai_1 _28274_ (.A1(_08889_),
    .A2(_08890_),
    .B1(_08891_),
    .B2(_08892_),
    .C1(net2705),
    .Y(_08893_));
 sky130_fd_sc_hd__nor2_1 _28275_ (.A(\inst$top.soc.cpu.gprf.mem[19][25] ),
    .B(net2370),
    .Y(_08894_));
 sky130_fd_sc_hd__o21ai_0 _28276_ (.A1(net2773),
    .A2(\inst$top.soc.cpu.gprf.mem[18][25] ),
    .B1(net2726),
    .Y(_08895_));
 sky130_fd_sc_hd__nor2_1 _28277_ (.A(net2772),
    .B(\inst$top.soc.cpu.gprf.mem[16][25] ),
    .Y(_08896_));
 sky130_fd_sc_hd__o21ai_0 _28278_ (.A1(\inst$top.soc.cpu.gprf.mem[17][25] ),
    .A2(net2370),
    .B1(net2325),
    .Y(_08897_));
 sky130_fd_sc_hd__o221ai_1 _28279_ (.A1(_08894_),
    .A2(_08895_),
    .B1(_08896_),
    .B2(_08897_),
    .C1(net2420),
    .Y(_08898_));
 sky130_fd_sc_hd__nand3_1 _28280_ (.A(_08893_),
    .B(_08898_),
    .C(net2433),
    .Y(_08899_));
 sky130_fd_sc_hd__a32oi_1 _28281_ (.A1(_08866_),
    .A2(_08877_),
    .A3(net2442),
    .B1(_08888_),
    .B2(_08899_),
    .Y(_00049_));
 sky130_fd_sc_hd__nor2_1 _28282_ (.A(\inst$top.soc.cpu.gprf.mem[23][26] ),
    .B(net2359),
    .Y(_08900_));
 sky130_fd_sc_hd__o21ai_0 _28283_ (.A1(net2759),
    .A2(\inst$top.soc.cpu.gprf.mem[22][26] ),
    .B1(net2720),
    .Y(_08901_));
 sky130_fd_sc_hd__nor2_1 _28284_ (.A(net2758),
    .B(\inst$top.soc.cpu.gprf.mem[20][26] ),
    .Y(_08902_));
 sky130_fd_sc_hd__o21ai_0 _28285_ (.A1(\inst$top.soc.cpu.gprf.mem[21][26] ),
    .A2(net2356),
    .B1(net2317),
    .Y(_08903_));
 sky130_fd_sc_hd__o221ai_1 _28286_ (.A1(_08900_),
    .A2(_08901_),
    .B1(_08902_),
    .B2(_08903_),
    .C1(net2702),
    .Y(_08904_));
 sky130_fd_sc_hd__nor2_1 _28287_ (.A(\inst$top.soc.cpu.gprf.mem[19][26] ),
    .B(net2358),
    .Y(_08905_));
 sky130_fd_sc_hd__o21ai_0 _28288_ (.A1(net2762),
    .A2(\inst$top.soc.cpu.gprf.mem[18][26] ),
    .B1(net2720),
    .Y(_08906_));
 sky130_fd_sc_hd__nor2_1 _28289_ (.A(net2761),
    .B(\inst$top.soc.cpu.gprf.mem[16][26] ),
    .Y(_08907_));
 sky130_fd_sc_hd__o21ai_0 _28290_ (.A1(\inst$top.soc.cpu.gprf.mem[17][26] ),
    .A2(net2358),
    .B1(net2317),
    .Y(_08908_));
 sky130_fd_sc_hd__o221ai_1 _28291_ (.A1(_08905_),
    .A2(_08906_),
    .B1(_08907_),
    .B2(_08908_),
    .C1(net2416),
    .Y(_08909_));
 sky130_fd_sc_hd__nand3_1 _28292_ (.A(_08904_),
    .B(_08909_),
    .C(net2430),
    .Y(_08910_));
 sky130_fd_sc_hd__nor2_1 _28293_ (.A(\inst$top.soc.cpu.gprf.mem[31][26] ),
    .B(net2358),
    .Y(_08911_));
 sky130_fd_sc_hd__o21ai_0 _28294_ (.A1(net2761),
    .A2(\inst$top.soc.cpu.gprf.mem[30][26] ),
    .B1(net2720),
    .Y(_08912_));
 sky130_fd_sc_hd__nor2_1 _28295_ (.A(net2761),
    .B(\inst$top.soc.cpu.gprf.mem[28][26] ),
    .Y(_08913_));
 sky130_fd_sc_hd__o21ai_0 _28296_ (.A1(\inst$top.soc.cpu.gprf.mem[29][26] ),
    .A2(net2359),
    .B1(net2317),
    .Y(_08914_));
 sky130_fd_sc_hd__o22ai_1 _28297_ (.A1(_08911_),
    .A2(_08912_),
    .B1(_08913_),
    .B2(_08914_),
    .Y(_08915_));
 sky130_fd_sc_hd__nand2_1 _28298_ (.A(net2761),
    .B(\inst$top.soc.cpu.gprf.mem[25][26] ),
    .Y(_08916_));
 sky130_fd_sc_hd__o21ai_0 _28299_ (.A1(net2761),
    .A2(_07239_),
    .B1(_08916_),
    .Y(_08917_));
 sky130_fd_sc_hd__nor2_1 _28300_ (.A(\inst$top.soc.cpu.gprf.mem[27][26] ),
    .B(net2358),
    .Y(_08918_));
 sky130_fd_sc_hd__o21ai_0 _28301_ (.A1(net2761),
    .A2(\inst$top.soc.cpu.gprf.mem[26][26] ),
    .B1(net2720),
    .Y(_08919_));
 sky130_fd_sc_hd__nor2_1 _28302_ (.A(_08918_),
    .B(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__a21oi_1 _28303_ (.A1(net2317),
    .A2(_08917_),
    .B1(_08920_),
    .Y(_08921_));
 sky130_fd_sc_hd__a21oi_1 _28304_ (.A1(_08921_),
    .A2(net2414),
    .B1(net2431),
    .Y(_08922_));
 sky130_fd_sc_hd__o21ai_0 _28305_ (.A1(net2414),
    .A2(_08915_),
    .B1(_08922_),
    .Y(_08923_));
 sky130_fd_sc_hd__nor2_1 _28306_ (.A(\inst$top.soc.cpu.gprf.mem[7][26] ),
    .B(net2358),
    .Y(_08924_));
 sky130_fd_sc_hd__o21ai_0 _28307_ (.A1(net2760),
    .A2(\inst$top.soc.cpu.gprf.mem[6][26] ),
    .B1(net2720),
    .Y(_08925_));
 sky130_fd_sc_hd__nor2_1 _28308_ (.A(net2760),
    .B(\inst$top.soc.cpu.gprf.mem[4][26] ),
    .Y(_08926_));
 sky130_fd_sc_hd__o21ai_0 _28309_ (.A1(\inst$top.soc.cpu.gprf.mem[5][26] ),
    .A2(net2358),
    .B1(net2317),
    .Y(_08927_));
 sky130_fd_sc_hd__o221ai_1 _28310_ (.A1(_08924_),
    .A2(_08925_),
    .B1(_08926_),
    .B2(_08927_),
    .C1(net2701),
    .Y(_08928_));
 sky130_fd_sc_hd__nor2_1 _28311_ (.A(\inst$top.soc.cpu.gprf.mem[3][26] ),
    .B(net2353),
    .Y(_08929_));
 sky130_fd_sc_hd__o21ai_0 _28312_ (.A1(net2760),
    .A2(\inst$top.soc.cpu.gprf.mem[2][26] ),
    .B1(net2720),
    .Y(_08930_));
 sky130_fd_sc_hd__nor2_1 _28313_ (.A(net2760),
    .B(\inst$top.soc.cpu.gprf.mem[0][26] ),
    .Y(_08931_));
 sky130_fd_sc_hd__o21ai_0 _28314_ (.A1(\inst$top.soc.cpu.gprf.mem[1][26] ),
    .A2(net2353),
    .B1(net2315),
    .Y(_08932_));
 sky130_fd_sc_hd__o221ai_1 _28315_ (.A1(_08929_),
    .A2(_08930_),
    .B1(_08931_),
    .B2(_08932_),
    .C1(net2413),
    .Y(_08933_));
 sky130_fd_sc_hd__a31oi_1 _28316_ (.A1(_08928_),
    .A2(_08933_),
    .A3(net2430),
    .B1(net2689),
    .Y(_08934_));
 sky130_fd_sc_hd__nor2_1 _28317_ (.A(\inst$top.soc.cpu.gprf.mem[15][26] ),
    .B(net2355),
    .Y(_08935_));
 sky130_fd_sc_hd__o21ai_0 _28318_ (.A1(net2757),
    .A2(\inst$top.soc.cpu.gprf.mem[14][26] ),
    .B1(net2719),
    .Y(_08936_));
 sky130_fd_sc_hd__nor2_1 _28319_ (.A(net2759),
    .B(\inst$top.soc.cpu.gprf.mem[12][26] ),
    .Y(_08937_));
 sky130_fd_sc_hd__o21ai_0 _28320_ (.A1(\inst$top.soc.cpu.gprf.mem[13][26] ),
    .A2(net2355),
    .B1(net2316),
    .Y(_08938_));
 sky130_fd_sc_hd__o221ai_1 _28321_ (.A1(_08935_),
    .A2(_08936_),
    .B1(_08937_),
    .B2(_08938_),
    .C1(net2701),
    .Y(_08939_));
 sky130_fd_sc_hd__nor2_1 _28322_ (.A(\inst$top.soc.cpu.gprf.mem[11][26] ),
    .B(net2357),
    .Y(_08940_));
 sky130_fd_sc_hd__o21ai_0 _28323_ (.A1(net2759),
    .A2(\inst$top.soc.cpu.gprf.mem[10][26] ),
    .B1(net2719),
    .Y(_08941_));
 sky130_fd_sc_hd__nor2_1 _28324_ (.A(net2757),
    .B(\inst$top.soc.cpu.gprf.mem[8][26] ),
    .Y(_08942_));
 sky130_fd_sc_hd__o21ai_0 _28325_ (.A1(\inst$top.soc.cpu.gprf.mem[9][26] ),
    .A2(net2357),
    .B1(net2316),
    .Y(_08943_));
 sky130_fd_sc_hd__o221ai_1 _28326_ (.A1(_08940_),
    .A2(_08941_),
    .B1(_08942_),
    .B2(_08943_),
    .C1(net2416),
    .Y(_08944_));
 sky130_fd_sc_hd__nand3_1 _28327_ (.A(_08939_),
    .B(_08944_),
    .C(net2695),
    .Y(_08945_));
 sky130_fd_sc_hd__a32oi_1 _28328_ (.A1(net2689),
    .A2(_08910_),
    .A3(_08923_),
    .B1(_08934_),
    .B2(_08945_),
    .Y(_00050_));
 sky130_fd_sc_hd__nor2_1 _28329_ (.A(\inst$top.soc.cpu.gprf.mem[31][27] ),
    .B(net2389),
    .Y(_08946_));
 sky130_fd_sc_hd__o21ai_0 _28330_ (.A1(net2794),
    .A2(\inst$top.soc.cpu.gprf.mem[30][27] ),
    .B1(net2737),
    .Y(_08947_));
 sky130_fd_sc_hd__nor2_1 _28331_ (.A(net2794),
    .B(\inst$top.soc.cpu.gprf.mem[28][27] ),
    .Y(_08948_));
 sky130_fd_sc_hd__o21ai_0 _28332_ (.A1(\inst$top.soc.cpu.gprf.mem[29][27] ),
    .A2(net2387),
    .B1(net2334),
    .Y(_08949_));
 sky130_fd_sc_hd__o22ai_1 _28333_ (.A1(_08946_),
    .A2(_08947_),
    .B1(_08948_),
    .B2(_08949_),
    .Y(_08950_));
 sky130_fd_sc_hd__nor2_1 _28334_ (.A(\inst$top.soc.cpu.gprf.mem[27][27] ),
    .B(net2387),
    .Y(_08951_));
 sky130_fd_sc_hd__o21ai_0 _28335_ (.A1(net2792),
    .A2(\inst$top.soc.cpu.gprf.mem[26][27] ),
    .B1(net2737),
    .Y(_08952_));
 sky130_fd_sc_hd__nor2_1 _28336_ (.A(net2792),
    .B(\inst$top.soc.cpu.gprf.mem[24][27] ),
    .Y(_08953_));
 sky130_fd_sc_hd__o21ai_0 _28337_ (.A1(\inst$top.soc.cpu.gprf.mem[25][27] ),
    .A2(net2387),
    .B1(net2334),
    .Y(_08954_));
 sky130_fd_sc_hd__o22ai_1 _28338_ (.A1(_08951_),
    .A2(_08952_),
    .B1(_08953_),
    .B2(_08954_),
    .Y(_08955_));
 sky130_fd_sc_hd__nor2_1 _28339_ (.A(net2710),
    .B(_08955_),
    .Y(_08956_));
 sky130_fd_sc_hd__nor2_1 _28340_ (.A(net2437),
    .B(_08956_),
    .Y(_08957_));
 sky130_fd_sc_hd__o21ai_0 _28341_ (.A1(net2423),
    .A2(_08950_),
    .B1(_08957_),
    .Y(_08958_));
 sky130_fd_sc_hd__nor2_1 _28342_ (.A(\inst$top.soc.cpu.gprf.mem[23][27] ),
    .B(net2389),
    .Y(_08959_));
 sky130_fd_sc_hd__o21ai_0 _28343_ (.A1(net2792),
    .A2(\inst$top.soc.cpu.gprf.mem[22][27] ),
    .B1(net2737),
    .Y(_08960_));
 sky130_fd_sc_hd__nor2_1 _28344_ (.A(net2794),
    .B(\inst$top.soc.cpu.gprf.mem[20][27] ),
    .Y(_08961_));
 sky130_fd_sc_hd__o21ai_0 _28345_ (.A1(\inst$top.soc.cpu.gprf.mem[21][27] ),
    .A2(net2387),
    .B1(net2334),
    .Y(_08962_));
 sky130_fd_sc_hd__o221ai_1 _28346_ (.A1(_08959_),
    .A2(_08960_),
    .B1(_08961_),
    .B2(_08962_),
    .C1(net2710),
    .Y(_08963_));
 sky130_fd_sc_hd__nor2_1 _28347_ (.A(\inst$top.soc.cpu.gprf.mem[19][27] ),
    .B(net2389),
    .Y(_08964_));
 sky130_fd_sc_hd__o21ai_0 _28348_ (.A1(net2794),
    .A2(\inst$top.soc.cpu.gprf.mem[18][27] ),
    .B1(net2737),
    .Y(_08965_));
 sky130_fd_sc_hd__nor2_1 _28349_ (.A(net2792),
    .B(\inst$top.soc.cpu.gprf.mem[16][27] ),
    .Y(_08966_));
 sky130_fd_sc_hd__o21ai_0 _28350_ (.A1(\inst$top.soc.cpu.gprf.mem[17][27] ),
    .A2(net2389),
    .B1(net2334),
    .Y(_08967_));
 sky130_fd_sc_hd__o221ai_1 _28351_ (.A1(_08964_),
    .A2(_08965_),
    .B1(_08966_),
    .B2(_08967_),
    .C1(net2423),
    .Y(_08968_));
 sky130_fd_sc_hd__nand3_1 _28352_ (.A(_08963_),
    .B(_08968_),
    .C(net2437),
    .Y(_08969_));
 sky130_fd_sc_hd__nor2_1 _28353_ (.A(\inst$top.soc.cpu.gprf.mem[11][27] ),
    .B(net2388),
    .Y(_08970_));
 sky130_fd_sc_hd__o21ai_0 _28354_ (.A1(net2793),
    .A2(\inst$top.soc.cpu.gprf.mem[10][27] ),
    .B1(net2739),
    .Y(_08971_));
 sky130_fd_sc_hd__nor2_1 _28355_ (.A(net2793),
    .B(\inst$top.soc.cpu.gprf.mem[8][27] ),
    .Y(_08972_));
 sky130_fd_sc_hd__o21ai_0 _28356_ (.A1(\inst$top.soc.cpu.gprf.mem[9][27] ),
    .A2(net2388),
    .B1(net2334),
    .Y(_08973_));
 sky130_fd_sc_hd__o221ai_1 _28357_ (.A1(_08970_),
    .A2(_08971_),
    .B1(_08972_),
    .B2(_08973_),
    .C1(net2423),
    .Y(_08974_));
 sky130_fd_sc_hd__nor2_1 _28358_ (.A(\inst$top.soc.cpu.gprf.mem[15][27] ),
    .B(net2387),
    .Y(_08975_));
 sky130_fd_sc_hd__o21ai_0 _28359_ (.A1(net2792),
    .A2(\inst$top.soc.cpu.gprf.mem[14][27] ),
    .B1(net2737),
    .Y(_08976_));
 sky130_fd_sc_hd__nor2_1 _28360_ (.A(net2792),
    .B(\inst$top.soc.cpu.gprf.mem[12][27] ),
    .Y(_08977_));
 sky130_fd_sc_hd__o21ai_0 _28361_ (.A1(\inst$top.soc.cpu.gprf.mem[13][27] ),
    .A2(net2387),
    .B1(net2334),
    .Y(_08978_));
 sky130_fd_sc_hd__o221ai_1 _28362_ (.A1(_08975_),
    .A2(_08976_),
    .B1(_08977_),
    .B2(_08978_),
    .C1(net2710),
    .Y(_08979_));
 sky130_fd_sc_hd__a31oi_1 _28363_ (.A1(_08974_),
    .A2(_08979_),
    .A3(net2698),
    .B1(net2691),
    .Y(_08980_));
 sky130_fd_sc_hd__nor2_1 _28364_ (.A(\inst$top.soc.cpu.gprf.mem[7][27] ),
    .B(net2387),
    .Y(_08981_));
 sky130_fd_sc_hd__o21ai_0 _28365_ (.A1(net2792),
    .A2(\inst$top.soc.cpu.gprf.mem[6][27] ),
    .B1(net2737),
    .Y(_08982_));
 sky130_fd_sc_hd__nor2_1 _28366_ (.A(net2792),
    .B(\inst$top.soc.cpu.gprf.mem[4][27] ),
    .Y(_08983_));
 sky130_fd_sc_hd__o21ai_0 _28367_ (.A1(\inst$top.soc.cpu.gprf.mem[5][27] ),
    .A2(net2387),
    .B1(net2334),
    .Y(_08984_));
 sky130_fd_sc_hd__o221ai_1 _28368_ (.A1(_08981_),
    .A2(_08982_),
    .B1(_08983_),
    .B2(_08984_),
    .C1(net2710),
    .Y(_08985_));
 sky130_fd_sc_hd__nor2_1 _28369_ (.A(\inst$top.soc.cpu.gprf.mem[3][27] ),
    .B(net2387),
    .Y(_08986_));
 sky130_fd_sc_hd__o21ai_0 _28370_ (.A1(net2792),
    .A2(\inst$top.soc.cpu.gprf.mem[2][27] ),
    .B1(net2737),
    .Y(_08987_));
 sky130_fd_sc_hd__nor2_1 _28371_ (.A(net2792),
    .B(\inst$top.soc.cpu.gprf.mem[0][27] ),
    .Y(_08988_));
 sky130_fd_sc_hd__o21ai_0 _28372_ (.A1(\inst$top.soc.cpu.gprf.mem[1][27] ),
    .A2(net2387),
    .B1(net2334),
    .Y(_08989_));
 sky130_fd_sc_hd__o221ai_1 _28373_ (.A1(_08986_),
    .A2(_08987_),
    .B1(_08988_),
    .B2(_08989_),
    .C1(net2423),
    .Y(_08990_));
 sky130_fd_sc_hd__nand3_1 _28374_ (.A(_08985_),
    .B(_08990_),
    .C(net2437),
    .Y(_08991_));
 sky130_fd_sc_hd__a32oi_1 _28375_ (.A1(net2691),
    .A2(_08958_),
    .A3(_08969_),
    .B1(_08980_),
    .B2(_08991_),
    .Y(_00051_));
 sky130_fd_sc_hd__nor2_1 _28376_ (.A(\inst$top.soc.cpu.gprf.mem[23][28] ),
    .B(net2390),
    .Y(_08992_));
 sky130_fd_sc_hd__o21ai_0 _28377_ (.A1(net2795),
    .A2(\inst$top.soc.cpu.gprf.mem[22][28] ),
    .B1(net2738),
    .Y(_08993_));
 sky130_fd_sc_hd__nor2_1 _28378_ (.A(net2795),
    .B(\inst$top.soc.cpu.gprf.mem[20][28] ),
    .Y(_08994_));
 sky130_fd_sc_hd__o21ai_0 _28379_ (.A1(\inst$top.soc.cpu.gprf.mem[21][28] ),
    .A2(net2390),
    .B1(net2335),
    .Y(_08995_));
 sky130_fd_sc_hd__o221ai_1 _28380_ (.A1(_08992_),
    .A2(_08993_),
    .B1(_08994_),
    .B2(_08995_),
    .C1(net2710),
    .Y(_08996_));
 sky130_fd_sc_hd__nor2_1 _28381_ (.A(\inst$top.soc.cpu.gprf.mem[19][28] ),
    .B(net2390),
    .Y(_08997_));
 sky130_fd_sc_hd__o21ai_0 _28382_ (.A1(net2795),
    .A2(\inst$top.soc.cpu.gprf.mem[18][28] ),
    .B1(net2738),
    .Y(_08998_));
 sky130_fd_sc_hd__nor2_1 _28383_ (.A(net2795),
    .B(\inst$top.soc.cpu.gprf.mem[16][28] ),
    .Y(_08999_));
 sky130_fd_sc_hd__o21ai_0 _28384_ (.A1(\inst$top.soc.cpu.gprf.mem[17][28] ),
    .A2(net2390),
    .B1(net2335),
    .Y(_09000_));
 sky130_fd_sc_hd__o221ai_1 _28385_ (.A1(_08997_),
    .A2(_08998_),
    .B1(_08999_),
    .B2(_09000_),
    .C1(net2423),
    .Y(_09001_));
 sky130_fd_sc_hd__nand3_1 _28386_ (.A(_08996_),
    .B(_09001_),
    .C(net2437),
    .Y(_09002_));
 sky130_fd_sc_hd__nor2_1 _28387_ (.A(\inst$top.soc.cpu.gprf.mem[31][28] ),
    .B(net2391),
    .Y(_09003_));
 sky130_fd_sc_hd__o21ai_0 _28388_ (.A1(net2796),
    .A2(\inst$top.soc.cpu.gprf.mem[30][28] ),
    .B1(net2738),
    .Y(_09004_));
 sky130_fd_sc_hd__nor2_1 _28389_ (.A(net2804),
    .B(\inst$top.soc.cpu.gprf.mem[28][28] ),
    .Y(_09005_));
 sky130_fd_sc_hd__o21ai_0 _28390_ (.A1(\inst$top.soc.cpu.gprf.mem[29][28] ),
    .A2(net2391),
    .B1(net2335),
    .Y(_09006_));
 sky130_fd_sc_hd__o22ai_1 _28391_ (.A1(_09003_),
    .A2(_09004_),
    .B1(_09005_),
    .B2(_09006_),
    .Y(_09007_));
 sky130_fd_sc_hd__nor2_1 _28392_ (.A(\inst$top.soc.cpu.gprf.mem[27][28] ),
    .B(net2390),
    .Y(_09008_));
 sky130_fd_sc_hd__o21ai_0 _28393_ (.A1(net2795),
    .A2(\inst$top.soc.cpu.gprf.mem[26][28] ),
    .B1(net2738),
    .Y(_09009_));
 sky130_fd_sc_hd__nor2_1 _28394_ (.A(net2804),
    .B(\inst$top.soc.cpu.gprf.mem[24][28] ),
    .Y(_09010_));
 sky130_fd_sc_hd__o21ai_0 _28395_ (.A1(\inst$top.soc.cpu.gprf.mem[25][28] ),
    .A2(net2390),
    .B1(net2339),
    .Y(_09011_));
 sky130_fd_sc_hd__o22ai_1 _28396_ (.A1(_09008_),
    .A2(_09009_),
    .B1(_09010_),
    .B2(_09011_),
    .Y(_09012_));
 sky130_fd_sc_hd__nor2_1 _28397_ (.A(net2710),
    .B(_09012_),
    .Y(_09013_));
 sky130_fd_sc_hd__nor2_1 _28398_ (.A(net2437),
    .B(_09013_),
    .Y(_09014_));
 sky130_fd_sc_hd__o21ai_0 _28399_ (.A1(net2425),
    .A2(_09007_),
    .B1(_09014_),
    .Y(_09015_));
 sky130_fd_sc_hd__nor2_1 _28400_ (.A(\inst$top.soc.cpu.gprf.mem[11][28] ),
    .B(net2391),
    .Y(_09016_));
 sky130_fd_sc_hd__o21ai_0 _28401_ (.A1(net2795),
    .A2(\inst$top.soc.cpu.gprf.mem[10][28] ),
    .B1(net2739),
    .Y(_09017_));
 sky130_fd_sc_hd__nor2_1 _28402_ (.A(net2795),
    .B(\inst$top.soc.cpu.gprf.mem[8][28] ),
    .Y(_09018_));
 sky130_fd_sc_hd__o21ai_0 _28403_ (.A1(\inst$top.soc.cpu.gprf.mem[9][28] ),
    .A2(net2390),
    .B1(net2339),
    .Y(_09019_));
 sky130_fd_sc_hd__o22ai_1 _28404_ (.A1(_09016_),
    .A2(_09017_),
    .B1(_09018_),
    .B2(_09019_),
    .Y(_09020_));
 sky130_fd_sc_hd__nor2_1 _28405_ (.A(net2710),
    .B(_09020_),
    .Y(_09021_));
 sky130_fd_sc_hd__nor2_1 _28406_ (.A(\inst$top.soc.cpu.gprf.mem[15][28] ),
    .B(net2391),
    .Y(_09022_));
 sky130_fd_sc_hd__o21ai_0 _28407_ (.A1(net2796),
    .A2(\inst$top.soc.cpu.gprf.mem[14][28] ),
    .B1(net2738),
    .Y(_09023_));
 sky130_fd_sc_hd__nor2_1 _28408_ (.A(net2796),
    .B(\inst$top.soc.cpu.gprf.mem[12][28] ),
    .Y(_09024_));
 sky130_fd_sc_hd__o21ai_0 _28409_ (.A1(\inst$top.soc.cpu.gprf.mem[13][28] ),
    .A2(net2391),
    .B1(net2339),
    .Y(_09025_));
 sky130_fd_sc_hd__o22ai_1 _28410_ (.A1(_09022_),
    .A2(_09023_),
    .B1(_09024_),
    .B2(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__o21ai_0 _28411_ (.A1(net2423),
    .A2(_09026_),
    .B1(net2698),
    .Y(_09027_));
 sky130_fd_sc_hd__nor2_1 _28412_ (.A(\inst$top.soc.cpu.gprf.mem[7][28] ),
    .B(net2391),
    .Y(_09028_));
 sky130_fd_sc_hd__o21ai_0 _28413_ (.A1(net2796),
    .A2(\inst$top.soc.cpu.gprf.mem[6][28] ),
    .B1(net2738),
    .Y(_09029_));
 sky130_fd_sc_hd__nor2_1 _28414_ (.A(net2796),
    .B(\inst$top.soc.cpu.gprf.mem[4][28] ),
    .Y(_09030_));
 sky130_fd_sc_hd__o21ai_0 _28415_ (.A1(\inst$top.soc.cpu.gprf.mem[5][28] ),
    .A2(net2391),
    .B1(net2335),
    .Y(_09031_));
 sky130_fd_sc_hd__o221ai_1 _28416_ (.A1(_09028_),
    .A2(_09029_),
    .B1(_09030_),
    .B2(_09031_),
    .C1(net2710),
    .Y(_09032_));
 sky130_fd_sc_hd__nor2_1 _28417_ (.A(\inst$top.soc.cpu.gprf.mem[3][28] ),
    .B(net2391),
    .Y(_09033_));
 sky130_fd_sc_hd__o21ai_0 _28418_ (.A1(net2796),
    .A2(\inst$top.soc.cpu.gprf.mem[2][28] ),
    .B1(net2738),
    .Y(_09034_));
 sky130_fd_sc_hd__nor2_1 _28419_ (.A(net2796),
    .B(\inst$top.soc.cpu.gprf.mem[0][28] ),
    .Y(_09035_));
 sky130_fd_sc_hd__o21ai_0 _28420_ (.A1(\inst$top.soc.cpu.gprf.mem[1][28] ),
    .A2(net2391),
    .B1(net2339),
    .Y(_09036_));
 sky130_fd_sc_hd__o221ai_1 _28421_ (.A1(_09033_),
    .A2(_09034_),
    .B1(_09035_),
    .B2(_09036_),
    .C1(net2425),
    .Y(_09037_));
 sky130_fd_sc_hd__nand3_1 _28422_ (.A(_09032_),
    .B(_09037_),
    .C(net2437),
    .Y(_09038_));
 sky130_fd_sc_hd__o21ai_0 _28423_ (.A1(_09021_),
    .A2(_09027_),
    .B1(_09038_),
    .Y(_09039_));
 sky130_fd_sc_hd__nor2_1 _28424_ (.A(net2691),
    .B(_09039_),
    .Y(_09040_));
 sky130_fd_sc_hd__a31oi_1 _28425_ (.A1(net2691),
    .A2(_09002_),
    .A3(_09015_),
    .B1(_09040_),
    .Y(_00052_));
 sky130_fd_sc_hd__nor2_1 _28426_ (.A(\inst$top.soc.cpu.gprf.mem[31][29] ),
    .B(net2383),
    .Y(_09041_));
 sky130_fd_sc_hd__o21ai_0 _28427_ (.A1(net2787),
    .A2(\inst$top.soc.cpu.gprf.mem[30][29] ),
    .B1(net2736),
    .Y(_09042_));
 sky130_fd_sc_hd__nor2_1 _28428_ (.A(net2787),
    .B(\inst$top.soc.cpu.gprf.mem[28][29] ),
    .Y(_09043_));
 sky130_fd_sc_hd__o21ai_0 _28429_ (.A1(\inst$top.soc.cpu.gprf.mem[29][29] ),
    .A2(net2383),
    .B1(net2331),
    .Y(_09044_));
 sky130_fd_sc_hd__o22ai_1 _28430_ (.A1(_09041_),
    .A2(_09042_),
    .B1(_09043_),
    .B2(_09044_),
    .Y(_09045_));
 sky130_fd_sc_hd__nor2_1 _28431_ (.A(\inst$top.soc.cpu.gprf.mem[27][29] ),
    .B(net2384),
    .Y(_09046_));
 sky130_fd_sc_hd__o21ai_0 _28432_ (.A1(net2787),
    .A2(\inst$top.soc.cpu.gprf.mem[26][29] ),
    .B1(net2734),
    .Y(_09047_));
 sky130_fd_sc_hd__nor2_1 _28433_ (.A(net2787),
    .B(\inst$top.soc.cpu.gprf.mem[24][29] ),
    .Y(_09048_));
 sky130_fd_sc_hd__o21ai_0 _28434_ (.A1(\inst$top.soc.cpu.gprf.mem[25][29] ),
    .A2(net2384),
    .B1(net2333),
    .Y(_09049_));
 sky130_fd_sc_hd__o22ai_1 _28435_ (.A1(_09046_),
    .A2(_09047_),
    .B1(_09048_),
    .B2(_09049_),
    .Y(_09050_));
 sky130_fd_sc_hd__nor2_1 _28436_ (.A(net2708),
    .B(_09050_),
    .Y(_09051_));
 sky130_fd_sc_hd__nor2_1 _28437_ (.A(net2436),
    .B(_09051_),
    .Y(_09052_));
 sky130_fd_sc_hd__o21ai_0 _28438_ (.A1(net2422),
    .A2(_09045_),
    .B1(_09052_),
    .Y(_09053_));
 sky130_fd_sc_hd__nor2_1 _28439_ (.A(\inst$top.soc.cpu.gprf.mem[23][29] ),
    .B(net2383),
    .Y(_09054_));
 sky130_fd_sc_hd__o21ai_0 _28440_ (.A1(net2788),
    .A2(\inst$top.soc.cpu.gprf.mem[22][29] ),
    .B1(net2734),
    .Y(_09055_));
 sky130_fd_sc_hd__nor2_1 _28441_ (.A(net2788),
    .B(\inst$top.soc.cpu.gprf.mem[20][29] ),
    .Y(_09056_));
 sky130_fd_sc_hd__o21ai_0 _28442_ (.A1(\inst$top.soc.cpu.gprf.mem[21][29] ),
    .A2(net2383),
    .B1(net2331),
    .Y(_09057_));
 sky130_fd_sc_hd__o221ai_1 _28443_ (.A1(_09054_),
    .A2(_09055_),
    .B1(_09056_),
    .B2(_09057_),
    .C1(net2708),
    .Y(_09058_));
 sky130_fd_sc_hd__nor2_1 _28444_ (.A(\inst$top.soc.cpu.gprf.mem[19][29] ),
    .B(net2384),
    .Y(_09059_));
 sky130_fd_sc_hd__o21ai_0 _28445_ (.A1(net2788),
    .A2(\inst$top.soc.cpu.gprf.mem[18][29] ),
    .B1(net2736),
    .Y(_09060_));
 sky130_fd_sc_hd__nor2_1 _28446_ (.A(net2788),
    .B(\inst$top.soc.cpu.gprf.mem[16][29] ),
    .Y(_09061_));
 sky130_fd_sc_hd__o21ai_0 _28447_ (.A1(\inst$top.soc.cpu.gprf.mem[17][29] ),
    .A2(net2384),
    .B1(net2333),
    .Y(_09062_));
 sky130_fd_sc_hd__o221ai_1 _28448_ (.A1(_09059_),
    .A2(_09060_),
    .B1(_09061_),
    .B2(_09062_),
    .C1(net2422),
    .Y(_09063_));
 sky130_fd_sc_hd__nand3_1 _28449_ (.A(_09058_),
    .B(_09063_),
    .C(net2435),
    .Y(_09064_));
 sky130_fd_sc_hd__nor2_1 _28450_ (.A(\inst$top.soc.cpu.gprf.mem[7][29] ),
    .B(net2385),
    .Y(_09065_));
 sky130_fd_sc_hd__o21ai_0 _28451_ (.A1(net2787),
    .A2(\inst$top.soc.cpu.gprf.mem[6][29] ),
    .B1(net2736),
    .Y(_09066_));
 sky130_fd_sc_hd__nor2_1 _28452_ (.A(net2788),
    .B(\inst$top.soc.cpu.gprf.mem[4][29] ),
    .Y(_09067_));
 sky130_fd_sc_hd__o21ai_0 _28453_ (.A1(\inst$top.soc.cpu.gprf.mem[5][29] ),
    .A2(net2384),
    .B1(net2331),
    .Y(_09068_));
 sky130_fd_sc_hd__o221ai_1 _28454_ (.A1(_09065_),
    .A2(_09066_),
    .B1(_09067_),
    .B2(_09068_),
    .C1(net2708),
    .Y(_09069_));
 sky130_fd_sc_hd__nor2_1 _28455_ (.A(\inst$top.soc.cpu.gprf.mem[3][29] ),
    .B(net2383),
    .Y(_09070_));
 sky130_fd_sc_hd__o21ai_0 _28456_ (.A1(net2787),
    .A2(\inst$top.soc.cpu.gprf.mem[2][29] ),
    .B1(net2734),
    .Y(_09071_));
 sky130_fd_sc_hd__nor2_1 _28457_ (.A(net2788),
    .B(\inst$top.soc.cpu.gprf.mem[0][29] ),
    .Y(_09072_));
 sky130_fd_sc_hd__o21ai_0 _28458_ (.A1(\inst$top.soc.cpu.gprf.mem[1][29] ),
    .A2(net2383),
    .B1(net2331),
    .Y(_09073_));
 sky130_fd_sc_hd__o221ai_1 _28459_ (.A1(_09070_),
    .A2(_09071_),
    .B1(_09072_),
    .B2(_09073_),
    .C1(net2422),
    .Y(_09074_));
 sky130_fd_sc_hd__a31oi_1 _28460_ (.A1(_09069_),
    .A2(_09074_),
    .A3(net2435),
    .B1(net2693),
    .Y(_09075_));
 sky130_fd_sc_hd__nor2_1 _28461_ (.A(\inst$top.soc.cpu.gprf.mem[15][29] ),
    .B(net2384),
    .Y(_09076_));
 sky130_fd_sc_hd__o21ai_0 _28462_ (.A1(net2787),
    .A2(\inst$top.soc.cpu.gprf.mem[14][29] ),
    .B1(net2734),
    .Y(_09077_));
 sky130_fd_sc_hd__nor2_1 _28463_ (.A(net2787),
    .B(\inst$top.soc.cpu.gprf.mem[12][29] ),
    .Y(_09078_));
 sky130_fd_sc_hd__o21ai_0 _28464_ (.A1(\inst$top.soc.cpu.gprf.mem[13][29] ),
    .A2(net2384),
    .B1(net2331),
    .Y(_09079_));
 sky130_fd_sc_hd__o22ai_1 _28465_ (.A1(_09076_),
    .A2(_09077_),
    .B1(_09078_),
    .B2(_09079_),
    .Y(_09080_));
 sky130_fd_sc_hd__nor2_1 _28466_ (.A(\inst$top.soc.cpu.gprf.mem[11][29] ),
    .B(net2384),
    .Y(_09081_));
 sky130_fd_sc_hd__o21ai_0 _28467_ (.A1(net2787),
    .A2(\inst$top.soc.cpu.gprf.mem[10][29] ),
    .B1(net2736),
    .Y(_09082_));
 sky130_fd_sc_hd__nor2_1 _28468_ (.A(net2787),
    .B(\inst$top.soc.cpu.gprf.mem[8][29] ),
    .Y(_09083_));
 sky130_fd_sc_hd__o21ai_0 _28469_ (.A1(\inst$top.soc.cpu.gprf.mem[9][29] ),
    .A2(net2384),
    .B1(net2333),
    .Y(_09084_));
 sky130_fd_sc_hd__o22ai_1 _28470_ (.A1(_09081_),
    .A2(_09082_),
    .B1(_09083_),
    .B2(_09084_),
    .Y(_09085_));
 sky130_fd_sc_hd__nor2_1 _28471_ (.A(net2708),
    .B(_09085_),
    .Y(_09086_));
 sky130_fd_sc_hd__nor2_1 _28472_ (.A(net2436),
    .B(_09086_),
    .Y(_09087_));
 sky130_fd_sc_hd__o21ai_0 _28473_ (.A1(net2422),
    .A2(_09080_),
    .B1(_09087_),
    .Y(_09088_));
 sky130_fd_sc_hd__a32oi_1 _28474_ (.A1(net2694),
    .A2(_09053_),
    .A3(_09064_),
    .B1(_09075_),
    .B2(_09088_),
    .Y(_00053_));
 sky130_fd_sc_hd__nor2_1 _28475_ (.A(\inst$top.soc.cpu.gprf.mem[31][30] ),
    .B(net2359),
    .Y(_09089_));
 sky130_fd_sc_hd__o21ai_0 _28476_ (.A1(net2761),
    .A2(\inst$top.soc.cpu.gprf.mem[30][30] ),
    .B1(net2720),
    .Y(_09090_));
 sky130_fd_sc_hd__nor2_1 _28477_ (.A(net2762),
    .B(\inst$top.soc.cpu.gprf.mem[28][30] ),
    .Y(_09091_));
 sky130_fd_sc_hd__o21ai_0 _28478_ (.A1(\inst$top.soc.cpu.gprf.mem[29][30] ),
    .A2(net2359),
    .B1(net2318),
    .Y(_09092_));
 sky130_fd_sc_hd__o22ai_1 _28479_ (.A1(_09089_),
    .A2(_09090_),
    .B1(_09091_),
    .B2(_09092_),
    .Y(_09093_));
 sky130_fd_sc_hd__nor2_1 _28480_ (.A(\inst$top.soc.cpu.gprf.mem[27][30] ),
    .B(net2370),
    .Y(_09094_));
 sky130_fd_sc_hd__o21ai_0 _28481_ (.A1(net2771),
    .A2(\inst$top.soc.cpu.gprf.mem[26][30] ),
    .B1(net2726),
    .Y(_09095_));
 sky130_fd_sc_hd__nor2_1 _28482_ (.A(net2773),
    .B(\inst$top.soc.cpu.gprf.mem[24][30] ),
    .Y(_09096_));
 sky130_fd_sc_hd__o21ai_0 _28483_ (.A1(\inst$top.soc.cpu.gprf.mem[25][30] ),
    .A2(net2368),
    .B1(net2324),
    .Y(_09097_));
 sky130_fd_sc_hd__o22ai_1 _28484_ (.A1(_09094_),
    .A2(_09095_),
    .B1(_09096_),
    .B2(_09097_),
    .Y(_09098_));
 sky130_fd_sc_hd__nor2_1 _28485_ (.A(net2704),
    .B(_09098_),
    .Y(_09099_));
 sky130_fd_sc_hd__nor2_1 _28486_ (.A(net2431),
    .B(_09099_),
    .Y(_09100_));
 sky130_fd_sc_hd__o21ai_0 _28487_ (.A1(net2415),
    .A2(_09093_),
    .B1(_09100_),
    .Y(_09101_));
 sky130_fd_sc_hd__nor2_1 _28488_ (.A(\inst$top.soc.cpu.gprf.mem[23][30] ),
    .B(net2377),
    .Y(_09102_));
 sky130_fd_sc_hd__o21ai_0 _28489_ (.A1(net2780),
    .A2(\inst$top.soc.cpu.gprf.mem[22][30] ),
    .B1(net2731),
    .Y(_09103_));
 sky130_fd_sc_hd__nor2_1 _28490_ (.A(net2780),
    .B(\inst$top.soc.cpu.gprf.mem[20][30] ),
    .Y(_09104_));
 sky130_fd_sc_hd__o21ai_0 _28491_ (.A1(\inst$top.soc.cpu.gprf.mem[21][30] ),
    .A2(net2377),
    .B1(net2329),
    .Y(_09105_));
 sky130_fd_sc_hd__o221ai_1 _28492_ (.A1(_09102_),
    .A2(_09103_),
    .B1(_09104_),
    .B2(_09105_),
    .C1(net2707),
    .Y(_09106_));
 sky130_fd_sc_hd__nor2_1 _28493_ (.A(\inst$top.soc.cpu.gprf.mem[19][30] ),
    .B(net2377),
    .Y(_09107_));
 sky130_fd_sc_hd__o21ai_0 _28494_ (.A1(net2773),
    .A2(\inst$top.soc.cpu.gprf.mem[18][30] ),
    .B1(net2731),
    .Y(_09108_));
 sky130_fd_sc_hd__nor2_1 _28495_ (.A(net2780),
    .B(\inst$top.soc.cpu.gprf.mem[16][30] ),
    .Y(_09109_));
 sky130_fd_sc_hd__o21ai_0 _28496_ (.A1(\inst$top.soc.cpu.gprf.mem[17][30] ),
    .A2(net2370),
    .B1(net2324),
    .Y(_09110_));
 sky130_fd_sc_hd__o221ai_1 _28497_ (.A1(_09107_),
    .A2(_09108_),
    .B1(_09109_),
    .B2(_09110_),
    .C1(net2421),
    .Y(_09111_));
 sky130_fd_sc_hd__nand3_1 _28498_ (.A(_09106_),
    .B(_09111_),
    .C(net2435),
    .Y(_09112_));
 sky130_fd_sc_hd__nor2_1 _28499_ (.A(\inst$top.soc.cpu.gprf.mem[11][30] ),
    .B(net2376),
    .Y(_09113_));
 sky130_fd_sc_hd__o21ai_0 _28500_ (.A1(net2772),
    .A2(\inst$top.soc.cpu.gprf.mem[10][30] ),
    .B1(net2731),
    .Y(_09114_));
 sky130_fd_sc_hd__nor2_1 _28501_ (.A(net2772),
    .B(\inst$top.soc.cpu.gprf.mem[8][30] ),
    .Y(_09115_));
 sky130_fd_sc_hd__o21ai_0 _28502_ (.A1(\inst$top.soc.cpu.gprf.mem[9][30] ),
    .A2(net2370),
    .B1(net2324),
    .Y(_09116_));
 sky130_fd_sc_hd__o221ai_1 _28503_ (.A1(_09113_),
    .A2(_09114_),
    .B1(_09115_),
    .B2(_09116_),
    .C1(net2421),
    .Y(_09117_));
 sky130_fd_sc_hd__nor2_1 _28504_ (.A(\inst$top.soc.cpu.gprf.mem[15][30] ),
    .B(net2368),
    .Y(_09118_));
 sky130_fd_sc_hd__o21ai_0 _28505_ (.A1(net2772),
    .A2(\inst$top.soc.cpu.gprf.mem[14][30] ),
    .B1(net2726),
    .Y(_09119_));
 sky130_fd_sc_hd__nor2_1 _28506_ (.A(net2773),
    .B(\inst$top.soc.cpu.gprf.mem[12][30] ),
    .Y(_09120_));
 sky130_fd_sc_hd__o21ai_0 _28507_ (.A1(\inst$top.soc.cpu.gprf.mem[13][30] ),
    .A2(net2368),
    .B1(net2324),
    .Y(_09121_));
 sky130_fd_sc_hd__o221ai_1 _28508_ (.A1(_09118_),
    .A2(_09119_),
    .B1(_09120_),
    .B2(_09121_),
    .C1(net2704),
    .Y(_09122_));
 sky130_fd_sc_hd__a31oi_1 _28509_ (.A1(_09117_),
    .A2(_09122_),
    .A3(net2697),
    .B1(net2694),
    .Y(_09123_));
 sky130_fd_sc_hd__nor2_1 _28510_ (.A(\inst$top.soc.cpu.gprf.mem[7][30] ),
    .B(net2361),
    .Y(_09124_));
 sky130_fd_sc_hd__o21ai_0 _28511_ (.A1(net2764),
    .A2(\inst$top.soc.cpu.gprf.mem[6][30] ),
    .B1(net2722),
    .Y(_09125_));
 sky130_fd_sc_hd__nor2_1 _28512_ (.A(net2764),
    .B(\inst$top.soc.cpu.gprf.mem[4][30] ),
    .Y(_09126_));
 sky130_fd_sc_hd__o21ai_0 _28513_ (.A1(\inst$top.soc.cpu.gprf.mem[5][30] ),
    .A2(net2361),
    .B1(net2319),
    .Y(_09127_));
 sky130_fd_sc_hd__o221ai_1 _28514_ (.A1(_09124_),
    .A2(_09125_),
    .B1(_09126_),
    .B2(_09127_),
    .C1(net2702),
    .Y(_09128_));
 sky130_fd_sc_hd__nor2_1 _28515_ (.A(\inst$top.soc.cpu.gprf.mem[3][30] ),
    .B(net2361),
    .Y(_09129_));
 sky130_fd_sc_hd__o21ai_0 _28516_ (.A1(net2780),
    .A2(\inst$top.soc.cpu.gprf.mem[2][30] ),
    .B1(net2731),
    .Y(_09130_));
 sky130_fd_sc_hd__nor2_1 _28517_ (.A(net2780),
    .B(\inst$top.soc.cpu.gprf.mem[0][30] ),
    .Y(_09131_));
 sky130_fd_sc_hd__o21ai_0 _28518_ (.A1(\inst$top.soc.cpu.gprf.mem[1][30] ),
    .A2(net2361),
    .B1(net2329),
    .Y(_09132_));
 sky130_fd_sc_hd__o221ai_1 _28519_ (.A1(_09129_),
    .A2(_09130_),
    .B1(_09131_),
    .B2(_09132_),
    .C1(net2415),
    .Y(_09133_));
 sky130_fd_sc_hd__nand3_1 _28520_ (.A(_09128_),
    .B(_09133_),
    .C(net2431),
    .Y(_09134_));
 sky130_fd_sc_hd__a32oi_1 _28521_ (.A1(net2694),
    .A2(_09101_),
    .A3(_09112_),
    .B1(_09123_),
    .B2(_09134_),
    .Y(_00055_));
 sky130_fd_sc_hd__nor2_1 _28522_ (.A(\inst$top.soc.cpu.gprf.mem[7][31] ),
    .B(net2381),
    .Y(_09135_));
 sky130_fd_sc_hd__o21ai_0 _28523_ (.A1(net2786),
    .A2(\inst$top.soc.cpu.gprf.mem[6][31] ),
    .B1(net2735),
    .Y(_09136_));
 sky130_fd_sc_hd__nor2_1 _28524_ (.A(net2786),
    .B(\inst$top.soc.cpu.gprf.mem[4][31] ),
    .Y(_09137_));
 sky130_fd_sc_hd__o21ai_0 _28525_ (.A1(\inst$top.soc.cpu.gprf.mem[5][31] ),
    .A2(net2381),
    .B1(net2332),
    .Y(_09138_));
 sky130_fd_sc_hd__o221ai_1 _28526_ (.A1(_09135_),
    .A2(_09136_),
    .B1(_09137_),
    .B2(_09138_),
    .C1(net2708),
    .Y(_09139_));
 sky130_fd_sc_hd__nor2_1 _28527_ (.A(\inst$top.soc.cpu.gprf.mem[3][31] ),
    .B(net2381),
    .Y(_09140_));
 sky130_fd_sc_hd__o21ai_0 _28528_ (.A1(net2786),
    .A2(\inst$top.soc.cpu.gprf.mem[2][31] ),
    .B1(net2735),
    .Y(_09141_));
 sky130_fd_sc_hd__nor2_1 _28529_ (.A(net2786),
    .B(\inst$top.soc.cpu.gprf.mem[0][31] ),
    .Y(_09142_));
 sky130_fd_sc_hd__o21ai_0 _28530_ (.A1(\inst$top.soc.cpu.gprf.mem[1][31] ),
    .A2(net2381),
    .B1(net2332),
    .Y(_09143_));
 sky130_fd_sc_hd__o221ai_1 _28531_ (.A1(_09140_),
    .A2(_09141_),
    .B1(_09142_),
    .B2(_09143_),
    .C1(net2422),
    .Y(_09144_));
 sky130_fd_sc_hd__nand3_1 _28532_ (.A(_09139_),
    .B(_09144_),
    .C(net2435),
    .Y(_09145_));
 sky130_fd_sc_hd__nor2_1 _28533_ (.A(\inst$top.soc.cpu.gprf.mem[11][31] ),
    .B(net2381),
    .Y(_09146_));
 sky130_fd_sc_hd__o21ai_0 _28534_ (.A1(net2790),
    .A2(\inst$top.soc.cpu.gprf.mem[10][31] ),
    .B1(net2735),
    .Y(_09147_));
 sky130_fd_sc_hd__nor2_1 _28535_ (.A(net2786),
    .B(\inst$top.soc.cpu.gprf.mem[8][31] ),
    .Y(_09148_));
 sky130_fd_sc_hd__o21ai_0 _28536_ (.A1(\inst$top.soc.cpu.gprf.mem[9][31] ),
    .A2(net2382),
    .B1(net2332),
    .Y(_09149_));
 sky130_fd_sc_hd__o22ai_1 _28537_ (.A1(_09146_),
    .A2(_09147_),
    .B1(_09148_),
    .B2(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__nor2_1 _28538_ (.A(\inst$top.soc.cpu.gprf.mem[15][31] ),
    .B(net2381),
    .Y(_09151_));
 sky130_fd_sc_hd__o21ai_0 _28539_ (.A1(net2786),
    .A2(\inst$top.soc.cpu.gprf.mem[14][31] ),
    .B1(net2735),
    .Y(_09152_));
 sky130_fd_sc_hd__nor2_1 _28540_ (.A(net2786),
    .B(\inst$top.soc.cpu.gprf.mem[12][31] ),
    .Y(_09153_));
 sky130_fd_sc_hd__o21ai_0 _28541_ (.A1(\inst$top.soc.cpu.gprf.mem[13][31] ),
    .A2(net2381),
    .B1(net2332),
    .Y(_09154_));
 sky130_fd_sc_hd__o22ai_1 _28542_ (.A1(_09151_),
    .A2(_09152_),
    .B1(_09153_),
    .B2(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__nor2_1 _28543_ (.A(net2422),
    .B(_09155_),
    .Y(_09156_));
 sky130_fd_sc_hd__nor2_1 _28544_ (.A(net2436),
    .B(_09156_),
    .Y(_09157_));
 sky130_fd_sc_hd__o21ai_0 _28545_ (.A1(net2708),
    .A2(_09150_),
    .B1(_09157_),
    .Y(_09158_));
 sky130_fd_sc_hd__nor2_1 _28546_ (.A(\inst$top.soc.cpu.gprf.mem[31][31] ),
    .B(net2398),
    .Y(_09159_));
 sky130_fd_sc_hd__o21ai_0 _28547_ (.A1(net2805),
    .A2(\inst$top.soc.cpu.gprf.mem[30][31] ),
    .B1(net2743),
    .Y(_09160_));
 sky130_fd_sc_hd__nor2_1 _28548_ (.A(net2805),
    .B(\inst$top.soc.cpu.gprf.mem[28][31] ),
    .Y(_09161_));
 sky130_fd_sc_hd__o21ai_0 _28549_ (.A1(\inst$top.soc.cpu.gprf.mem[29][31] ),
    .A2(net2398),
    .B1(net2340),
    .Y(_09162_));
 sky130_fd_sc_hd__o22ai_1 _28550_ (.A1(_09159_),
    .A2(_09160_),
    .B1(_09161_),
    .B2(_09162_),
    .Y(_09163_));
 sky130_fd_sc_hd__nor2_1 _28551_ (.A(net2426),
    .B(_09163_),
    .Y(_09164_));
 sky130_fd_sc_hd__nor2_1 _28552_ (.A(\inst$top.soc.cpu.gprf.mem[27][31] ),
    .B(net2398),
    .Y(_09165_));
 sky130_fd_sc_hd__o21ai_0 _28553_ (.A1(net2805),
    .A2(\inst$top.soc.cpu.gprf.mem[26][31] ),
    .B1(net2743),
    .Y(_09166_));
 sky130_fd_sc_hd__nor2_1 _28554_ (.A(net2805),
    .B(\inst$top.soc.cpu.gprf.mem[24][31] ),
    .Y(_09167_));
 sky130_fd_sc_hd__o21ai_0 _28555_ (.A1(\inst$top.soc.cpu.gprf.mem[25][31] ),
    .A2(net2398),
    .B1(net2340),
    .Y(_09168_));
 sky130_fd_sc_hd__o22ai_1 _28556_ (.A1(_09165_),
    .A2(_09166_),
    .B1(_09167_),
    .B2(_09168_),
    .Y(_09169_));
 sky130_fd_sc_hd__o21ai_0 _28557_ (.A1(net2713),
    .A2(_09169_),
    .B1(net2698),
    .Y(_09170_));
 sky130_fd_sc_hd__nor2_1 _28558_ (.A(\inst$top.soc.cpu.gprf.mem[23][31] ),
    .B(net2381),
    .Y(_09171_));
 sky130_fd_sc_hd__o21ai_0 _28559_ (.A1(net2805),
    .A2(\inst$top.soc.cpu.gprf.mem[22][31] ),
    .B1(net2743),
    .Y(_09172_));
 sky130_fd_sc_hd__nor2_1 _28560_ (.A(net2786),
    .B(\inst$top.soc.cpu.gprf.mem[20][31] ),
    .Y(_09173_));
 sky130_fd_sc_hd__o21ai_0 _28561_ (.A1(\inst$top.soc.cpu.gprf.mem[21][31] ),
    .A2(net2381),
    .B1(net2332),
    .Y(_09174_));
 sky130_fd_sc_hd__o221ai_1 _28562_ (.A1(_09171_),
    .A2(_09172_),
    .B1(_09173_),
    .B2(_09174_),
    .C1(net2713),
    .Y(_09175_));
 sky130_fd_sc_hd__nor2_1 _28563_ (.A(\inst$top.soc.cpu.gprf.mem[19][31] ),
    .B(net2381),
    .Y(_09176_));
 sky130_fd_sc_hd__o21ai_0 _28564_ (.A1(net2805),
    .A2(\inst$top.soc.cpu.gprf.mem[18][31] ),
    .B1(net2743),
    .Y(_09177_));
 sky130_fd_sc_hd__nor2_1 _28565_ (.A(net2805),
    .B(\inst$top.soc.cpu.gprf.mem[16][31] ),
    .Y(_09178_));
 sky130_fd_sc_hd__o21ai_0 _28566_ (.A1(\inst$top.soc.cpu.gprf.mem[17][31] ),
    .A2(net2398),
    .B1(net2340),
    .Y(_09179_));
 sky130_fd_sc_hd__o221ai_1 _28567_ (.A1(_09176_),
    .A2(_09177_),
    .B1(_09178_),
    .B2(_09179_),
    .C1(net2426),
    .Y(_09180_));
 sky130_fd_sc_hd__nand3_1 _28568_ (.A(_09175_),
    .B(_09180_),
    .C(net2439),
    .Y(_09181_));
 sky130_fd_sc_hd__o21ai_0 _28569_ (.A1(_09164_),
    .A2(_09170_),
    .B1(_09181_),
    .Y(_09182_));
 sky130_fd_sc_hd__nor2_1 _28570_ (.A(net2443),
    .B(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__a31oi_1 _28571_ (.A1(net2443),
    .A2(_09145_),
    .A3(_09158_),
    .B1(_09183_),
    .Y(_00056_));
 sky130_fd_sc_hd__inv_2 _28572_ (.A(_02851_),
    .Y(_02542_));
 sky130_fd_sc_hd__inv_1 _28573_ (.A(net3032),
    .Y(_09184_));
 sky130_fd_sc_hd__nand2_1 _28575_ (.A(net2190),
    .B(_00096_),
    .Y(_09186_));
 sky130_fd_sc_hd__nand2_1 _28576_ (.A(_00064_),
    .B(net3030),
    .Y(_09187_));
 sky130_fd_sc_hd__nand2_1 _28577_ (.A(_09186_),
    .B(_09187_),
    .Y(\inst$top.soc.sram.read_port__data[0] ));
 sky130_fd_sc_hd__nand2_1 _28578_ (.A(net2190),
    .B(_00107_),
    .Y(_09188_));
 sky130_fd_sc_hd__nand2_1 _28580_ (.A(net3030),
    .B(_00075_),
    .Y(_09190_));
 sky130_fd_sc_hd__nand2_1 _28581_ (.A(_09188_),
    .B(_09190_),
    .Y(\inst$top.soc.sram.read_port__data[1] ));
 sky130_fd_sc_hd__nand2_1 _28583_ (.A(net2190),
    .B(_00118_),
    .Y(_09192_));
 sky130_fd_sc_hd__nand2_1 _28585_ (.A(net3030),
    .B(_00086_),
    .Y(_09194_));
 sky130_fd_sc_hd__nand2_1 _28586_ (.A(_09192_),
    .B(_09194_),
    .Y(\inst$top.soc.sram.read_port__data[2] ));
 sky130_fd_sc_hd__nand2_1 _28587_ (.A(net2190),
    .B(_00121_),
    .Y(_09195_));
 sky130_fd_sc_hd__nand2_1 _28588_ (.A(net3030),
    .B(_00089_),
    .Y(_09196_));
 sky130_fd_sc_hd__nand2_1 _28589_ (.A(_09195_),
    .B(_09196_),
    .Y(\inst$top.soc.sram.read_port__data[3] ));
 sky130_fd_sc_hd__nand2_1 _28590_ (.A(net2190),
    .B(_00122_),
    .Y(_09197_));
 sky130_fd_sc_hd__nand2_1 _28591_ (.A(net3030),
    .B(_00090_),
    .Y(_09198_));
 sky130_fd_sc_hd__nand2_1 _28592_ (.A(_09197_),
    .B(_09198_),
    .Y(\inst$top.soc.sram.read_port__data[4] ));
 sky130_fd_sc_hd__nand2_1 _28593_ (.A(net2191),
    .B(_00123_),
    .Y(_09199_));
 sky130_fd_sc_hd__nand2_1 _28594_ (.A(net3031),
    .B(_00091_),
    .Y(_09200_));
 sky130_fd_sc_hd__nand2_1 _28595_ (.A(_09199_),
    .B(_09200_),
    .Y(\inst$top.soc.sram.read_port__data[5] ));
 sky130_fd_sc_hd__nand2_1 _28596_ (.A(net2191),
    .B(_00124_),
    .Y(_09201_));
 sky130_fd_sc_hd__nand2_1 _28597_ (.A(net3031),
    .B(_00092_),
    .Y(_09202_));
 sky130_fd_sc_hd__nand2_1 _28598_ (.A(_09201_),
    .B(_09202_),
    .Y(\inst$top.soc.sram.read_port__data[6] ));
 sky130_fd_sc_hd__nand2_1 _28599_ (.A(net2192),
    .B(_00125_),
    .Y(_09203_));
 sky130_fd_sc_hd__nand2_1 _28600_ (.A(net3033),
    .B(_00093_),
    .Y(_09204_));
 sky130_fd_sc_hd__nand2_1 _28601_ (.A(_09203_),
    .B(_09204_),
    .Y(\inst$top.soc.sram.read_port__data[7] ));
 sky130_fd_sc_hd__nand2_1 _28602_ (.A(net2192),
    .B(_00126_),
    .Y(_09205_));
 sky130_fd_sc_hd__nand2_1 _28603_ (.A(net3033),
    .B(_00094_),
    .Y(_09206_));
 sky130_fd_sc_hd__nand2_1 _28604_ (.A(_09205_),
    .B(_09206_),
    .Y(\inst$top.soc.sram.read_port__data[8] ));
 sky130_fd_sc_hd__nand2_1 _28605_ (.A(net2192),
    .B(_00127_),
    .Y(_09207_));
 sky130_fd_sc_hd__nand2_1 _28606_ (.A(net3032),
    .B(_00095_),
    .Y(_09208_));
 sky130_fd_sc_hd__nand2_1 _28607_ (.A(_09207_),
    .B(_09208_),
    .Y(\inst$top.soc.sram.read_port__data[9] ));
 sky130_fd_sc_hd__nand2_1 _28608_ (.A(net2191),
    .B(_00097_),
    .Y(_09209_));
 sky130_fd_sc_hd__nand2_1 _28609_ (.A(net3031),
    .B(_00065_),
    .Y(_09210_));
 sky130_fd_sc_hd__nand2_1 _28610_ (.A(_09209_),
    .B(_09210_),
    .Y(\inst$top.soc.sram.read_port__data[10] ));
 sky130_fd_sc_hd__nand2_1 _28612_ (.A(net2192),
    .B(_00098_),
    .Y(_09212_));
 sky130_fd_sc_hd__nand2_1 _28613_ (.A(net3032),
    .B(_00066_),
    .Y(_09213_));
 sky130_fd_sc_hd__nand2_1 _28614_ (.A(_09212_),
    .B(_09213_),
    .Y(\inst$top.soc.sram.read_port__data[11] ));
 sky130_fd_sc_hd__nand2_1 _28615_ (.A(net2191),
    .B(_00099_),
    .Y(_09214_));
 sky130_fd_sc_hd__nand2_1 _28616_ (.A(net3033),
    .B(_00067_),
    .Y(_09215_));
 sky130_fd_sc_hd__nand2_1 _28617_ (.A(_09214_),
    .B(_09215_),
    .Y(\inst$top.soc.sram.read_port__data[12] ));
 sky130_fd_sc_hd__nand2_1 _28618_ (.A(net2190),
    .B(_00100_),
    .Y(_09216_));
 sky130_fd_sc_hd__nand2_1 _28619_ (.A(net3031),
    .B(_00068_),
    .Y(_09217_));
 sky130_fd_sc_hd__nand2_1 _28620_ (.A(_09216_),
    .B(_09217_),
    .Y(\inst$top.soc.sram.read_port__data[13] ));
 sky130_fd_sc_hd__nand2_1 _28621_ (.A(net2193),
    .B(_00101_),
    .Y(_09218_));
 sky130_fd_sc_hd__nand2_1 _28623_ (.A(net3033),
    .B(_00069_),
    .Y(_09220_));
 sky130_fd_sc_hd__nand2_1 _28624_ (.A(_09218_),
    .B(_09220_),
    .Y(\inst$top.soc.sram.read_port__data[14] ));
 sky130_fd_sc_hd__nand2_1 _28625_ (.A(net2192),
    .B(_00102_),
    .Y(_09221_));
 sky130_fd_sc_hd__nand2_1 _28626_ (.A(net3033),
    .B(_00070_),
    .Y(_09222_));
 sky130_fd_sc_hd__nand2_1 _28627_ (.A(_09221_),
    .B(_09222_),
    .Y(\inst$top.soc.sram.read_port__data[15] ));
 sky130_fd_sc_hd__nand2_1 _28628_ (.A(net2193),
    .B(_00103_),
    .Y(_09223_));
 sky130_fd_sc_hd__nand2_1 _28629_ (.A(net3032),
    .B(_00071_),
    .Y(_09224_));
 sky130_fd_sc_hd__nand2_1 _28630_ (.A(_09223_),
    .B(_09224_),
    .Y(\inst$top.soc.sram.read_port__data[16] ));
 sky130_fd_sc_hd__nand2_1 _28631_ (.A(net2193),
    .B(_00104_),
    .Y(_09225_));
 sky130_fd_sc_hd__nand2_1 _28632_ (.A(net3032),
    .B(_00072_),
    .Y(_09226_));
 sky130_fd_sc_hd__nand2_1 _28633_ (.A(_09225_),
    .B(_09226_),
    .Y(\inst$top.soc.sram.read_port__data[17] ));
 sky130_fd_sc_hd__nand2_1 _28634_ (.A(net2193),
    .B(_00105_),
    .Y(_09227_));
 sky130_fd_sc_hd__nand2_1 _28635_ (.A(net3033),
    .B(_00073_),
    .Y(_09228_));
 sky130_fd_sc_hd__nand2_1 _28636_ (.A(_09227_),
    .B(_09228_),
    .Y(\inst$top.soc.sram.read_port__data[18] ));
 sky130_fd_sc_hd__nand2_1 _28637_ (.A(net2193),
    .B(_00106_),
    .Y(_09229_));
 sky130_fd_sc_hd__nand2_1 _28638_ (.A(net3032),
    .B(_00074_),
    .Y(_09230_));
 sky130_fd_sc_hd__nand2_1 _28639_ (.A(_09229_),
    .B(_09230_),
    .Y(\inst$top.soc.sram.read_port__data[19] ));
 sky130_fd_sc_hd__nand2_1 _28640_ (.A(net2193),
    .B(_00108_),
    .Y(_09231_));
 sky130_fd_sc_hd__nand2_1 _28641_ (.A(net3033),
    .B(_00076_),
    .Y(_09232_));
 sky130_fd_sc_hd__nand2_1 _28642_ (.A(_09231_),
    .B(_09232_),
    .Y(\inst$top.soc.sram.read_port__data[20] ));
 sky130_fd_sc_hd__nand2_1 _28643_ (.A(net2192),
    .B(_00109_),
    .Y(_09233_));
 sky130_fd_sc_hd__nand2_1 _28644_ (.A(net3032),
    .B(_00077_),
    .Y(_09234_));
 sky130_fd_sc_hd__nand2_1 _28645_ (.A(_09233_),
    .B(_09234_),
    .Y(\inst$top.soc.sram.read_port__data[21] ));
 sky130_fd_sc_hd__nand2_1 _28646_ (.A(net2192),
    .B(_00110_),
    .Y(_09235_));
 sky130_fd_sc_hd__nand2_1 _28647_ (.A(net3032),
    .B(_00078_),
    .Y(_09236_));
 sky130_fd_sc_hd__nand2_1 _28648_ (.A(_09235_),
    .B(_09236_),
    .Y(\inst$top.soc.sram.read_port__data[22] ));
 sky130_fd_sc_hd__nand2_1 _28649_ (.A(net2192),
    .B(_00111_),
    .Y(_09237_));
 sky130_fd_sc_hd__nand2_1 _28650_ (.A(net3032),
    .B(_00079_),
    .Y(_09238_));
 sky130_fd_sc_hd__nand2_1 _28651_ (.A(_09237_),
    .B(_09238_),
    .Y(\inst$top.soc.sram.read_port__data[23] ));
 sky130_fd_sc_hd__nand2_1 _28652_ (.A(net2190),
    .B(_00112_),
    .Y(_09239_));
 sky130_fd_sc_hd__nand2_1 _28653_ (.A(net3030),
    .B(_00080_),
    .Y(_09240_));
 sky130_fd_sc_hd__nand2_1 _28654_ (.A(_09239_),
    .B(_09240_),
    .Y(\inst$top.soc.sram.read_port__data[24] ));
 sky130_fd_sc_hd__nand2_1 _28655_ (.A(net2190),
    .B(_00113_),
    .Y(_09241_));
 sky130_fd_sc_hd__nand2_1 _28656_ (.A(net3030),
    .B(_00081_),
    .Y(_09242_));
 sky130_fd_sc_hd__nand2_1 _28657_ (.A(_09241_),
    .B(_09242_),
    .Y(\inst$top.soc.sram.read_port__data[25] ));
 sky130_fd_sc_hd__nand2_1 _28658_ (.A(net2190),
    .B(_00114_),
    .Y(_09243_));
 sky130_fd_sc_hd__nand2_1 _28659_ (.A(net3030),
    .B(_00082_),
    .Y(_09244_));
 sky130_fd_sc_hd__nand2_1 _28660_ (.A(_09243_),
    .B(_09244_),
    .Y(\inst$top.soc.sram.read_port__data[26] ));
 sky130_fd_sc_hd__nand2_1 _28661_ (.A(net2190),
    .B(_00115_),
    .Y(_09245_));
 sky130_fd_sc_hd__nand2_1 _28662_ (.A(net3030),
    .B(_00083_),
    .Y(_09246_));
 sky130_fd_sc_hd__nand2_1 _28663_ (.A(_09245_),
    .B(_09246_),
    .Y(\inst$top.soc.sram.read_port__data[27] ));
 sky130_fd_sc_hd__nand2_1 _28664_ (.A(net2191),
    .B(_00116_),
    .Y(_09247_));
 sky130_fd_sc_hd__nand2_1 _28665_ (.A(net3030),
    .B(_00084_),
    .Y(_09248_));
 sky130_fd_sc_hd__nand2_1 _28666_ (.A(_09247_),
    .B(_09248_),
    .Y(\inst$top.soc.sram.read_port__data[28] ));
 sky130_fd_sc_hd__nand2_1 _28667_ (.A(net2192),
    .B(_00117_),
    .Y(_09249_));
 sky130_fd_sc_hd__nand2_1 _28668_ (.A(net3032),
    .B(_00085_),
    .Y(_09250_));
 sky130_fd_sc_hd__nand2_1 _28669_ (.A(_09249_),
    .B(_09250_),
    .Y(\inst$top.soc.sram.read_port__data[29] ));
 sky130_fd_sc_hd__nand2_1 _28670_ (.A(net2191),
    .B(_00119_),
    .Y(_09251_));
 sky130_fd_sc_hd__nand2_1 _28671_ (.A(net3031),
    .B(_00087_),
    .Y(_09252_));
 sky130_fd_sc_hd__nand2_1 _28672_ (.A(_09251_),
    .B(_09252_),
    .Y(\inst$top.soc.sram.read_port__data[30] ));
 sky130_fd_sc_hd__nand2_1 _28673_ (.A(net2192),
    .B(_00120_),
    .Y(_09253_));
 sky130_fd_sc_hd__nand2_1 _28674_ (.A(net3033),
    .B(_00088_),
    .Y(_09254_));
 sky130_fd_sc_hd__nand2_1 _28675_ (.A(_09253_),
    .B(_09254_),
    .Y(\inst$top.soc.sram.read_port__data[31] ));
 sky130_fd_sc_hd__inv_1 _28676_ (.A(\inst$top.soc.cpu.loadstore.dbus__sel[1] ),
    .Y(_09255_));
 sky130_fd_sc_hd__nand2_1 _28677_ (.A(net2566),
    .B(\inst$top.soc.cpu.loadstore.dbus__we ),
    .Y(_09256_));
 sky130_fd_sc_hd__nand2_1 _28678_ (.A(net2556),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[18] ),
    .Y(_09257_));
 sky130_fd_sc_hd__nand2_1 _28679_ (.A(net2559),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[18] ),
    .Y(_09258_));
 sky130_fd_sc_hd__nand2_1 _28680_ (.A(_09257_),
    .B(_09258_),
    .Y(_09259_));
 sky130_fd_sc_hd__or2_2 _28681_ (.A(\inst$top.soc.cpu.loadstore.dbus__adr[19] ),
    .B(net2556),
    .X(_09260_));
 sky130_fd_sc_hd__o21a_1 _28682_ (.A1(net2559),
    .A2(\inst$top.soc.cpu.fetch.ibus__adr[19] ),
    .B1(_09260_),
    .X(_09261_));
 sky130_fd_sc_hd__nor2_1 _28683_ (.A(_09259_),
    .B(_09261_),
    .Y(_09262_));
 sky130_fd_sc_hd__nand2_1 _28684_ (.A(net2557),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[21] ),
    .Y(_09263_));
 sky130_fd_sc_hd__nand2_1 _28685_ (.A(net2560),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[21] ),
    .Y(_09264_));
 sky130_fd_sc_hd__nand2_1 _28686_ (.A(_09263_),
    .B(_09264_),
    .Y(_09265_));
 sky130_fd_sc_hd__nand2_1 _28687_ (.A(net2556),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[20] ),
    .Y(_09266_));
 sky130_fd_sc_hd__nand2_1 _28688_ (.A(net2560),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[20] ),
    .Y(_09267_));
 sky130_fd_sc_hd__nand2_1 _28689_ (.A(_09266_),
    .B(_09267_),
    .Y(_09268_));
 sky130_fd_sc_hd__nor2_1 _28690_ (.A(_09265_),
    .B(_09268_),
    .Y(_09269_));
 sky130_fd_sc_hd__nand2_1 _28691_ (.A(_09262_),
    .B(_09269_),
    .Y(_09270_));
 sky130_fd_sc_hd__inv_1 _28692_ (.A(\inst$top.soc.cpu.loadstore.dbus__adr[25] ),
    .Y(_09271_));
 sky130_fd_sc_hd__nand2_1 _28693_ (.A(_09271_),
    .B(net2561),
    .Y(_09272_));
 sky130_fd_sc_hd__o21ai_0 _28694_ (.A1(net2561),
    .A2(\inst$top.soc.cpu.fetch.ibus__adr[25] ),
    .B1(_09272_),
    .Y(_09273_));
 sky130_fd_sc_hd__inv_1 _28695_ (.A(\inst$top.soc.cpu.loadstore.dbus__adr[24] ),
    .Y(_09274_));
 sky130_fd_sc_hd__nand2_1 _28696_ (.A(_09274_),
    .B(net2561),
    .Y(_09275_));
 sky130_fd_sc_hd__o21ai_0 _28697_ (.A1(net2561),
    .A2(\inst$top.soc.cpu.fetch.ibus__adr[24] ),
    .B1(_09275_),
    .Y(_09276_));
 sky130_fd_sc_hd__nand2_1 _28698_ (.A(_09273_),
    .B(_09276_),
    .Y(_09277_));
 sky130_fd_sc_hd__nand2_1 _28699_ (.A(net2557),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[27] ),
    .Y(_09278_));
 sky130_fd_sc_hd__nand2_1 _28700_ (.A(net2561),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[27] ),
    .Y(_09279_));
 sky130_fd_sc_hd__nand2_1 _28701_ (.A(_09278_),
    .B(_09279_),
    .Y(_09280_));
 sky130_fd_sc_hd__nand2_1 _28702_ (.A(net2556),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[8] ),
    .Y(_09281_));
 sky130_fd_sc_hd__nand2_1 _28703_ (.A(net2560),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[8] ),
    .Y(_09282_));
 sky130_fd_sc_hd__nand2_1 _28704_ (.A(_09281_),
    .B(_09282_),
    .Y(_09283_));
 sky130_fd_sc_hd__or2_2 _28705_ (.A(\inst$top.soc.cpu.loadstore.dbus__adr[9] ),
    .B(net2555),
    .X(_09284_));
 sky130_fd_sc_hd__o21ai_0 _28706_ (.A1(net2558),
    .A2(\inst$top.soc.cpu.fetch.ibus__adr[9] ),
    .B1(_09284_),
    .Y(_09285_));
 sky130_fd_sc_hd__inv_1 _28707_ (.A(_09285_),
    .Y(_09286_));
 sky130_fd_sc_hd__nor2_1 _28708_ (.A(_09283_),
    .B(_09286_),
    .Y(_09287_));
 sky130_fd_sc_hd__inv_1 _28709_ (.A(_09287_),
    .Y(_09288_));
 sky130_fd_sc_hd__mux2i_1 _28710_ (.A0(\inst$top.soc.cpu.fetch.ibus__adr[15] ),
    .A1(\inst$top.soc.cpu.loadstore.dbus__adr[15] ),
    .S(net2560),
    .Y(_09289_));
 sky130_fd_sc_hd__inv_1 _28711_ (.A(_09289_),
    .Y(_09290_));
 sky130_fd_sc_hd__mux2i_1 _28712_ (.A0(\inst$top.soc.cpu.fetch.ibus__adr[14] ),
    .A1(\inst$top.soc.cpu.loadstore.dbus__adr[14] ),
    .S(net2559),
    .Y(_09291_));
 sky130_fd_sc_hd__inv_1 _28713_ (.A(_09291_),
    .Y(_09292_));
 sky130_fd_sc_hd__nor2_1 _28714_ (.A(_09290_),
    .B(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__inv_1 _28715_ (.A(_09293_),
    .Y(_09294_));
 sky130_fd_sc_hd__nor2_1 _28716_ (.A(_09288_),
    .B(_09294_),
    .Y(_09295_));
 sky130_fd_sc_hd__nand2_1 _28717_ (.A(net2556),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[23] ),
    .Y(_09296_));
 sky130_fd_sc_hd__nand2_1 _28718_ (.A(net2560),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[23] ),
    .Y(_09297_));
 sky130_fd_sc_hd__nand2_1 _28719_ (.A(_09296_),
    .B(_09297_),
    .Y(_09298_));
 sky130_fd_sc_hd__or2_2 _28720_ (.A(\inst$top.soc.cpu.loadstore.dbus__adr[22] ),
    .B(net2557),
    .X(_09299_));
 sky130_fd_sc_hd__o21a_1 _28721_ (.A1(net2561),
    .A2(\inst$top.soc.cpu.fetch.ibus__adr[22] ),
    .B1(_09299_),
    .X(_09300_));
 sky130_fd_sc_hd__nor2_1 _28722_ (.A(_09298_),
    .B(_09300_),
    .Y(_09301_));
 sky130_fd_sc_hd__nand2_1 _28723_ (.A(net2557),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[26] ),
    .Y(_09302_));
 sky130_fd_sc_hd__nand2_1 _28724_ (.A(net2561),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[26] ),
    .Y(_09303_));
 sky130_fd_sc_hd__nand2_1 _28725_ (.A(_09302_),
    .B(_09303_),
    .Y(_09304_));
 sky130_fd_sc_hd__nand3_1 _28726_ (.A(_09295_),
    .B(_09301_),
    .C(_09304_),
    .Y(_09305_));
 sky130_fd_sc_hd__nor4_1 _28727_ (.A(_09270_),
    .B(_09277_),
    .C(_09280_),
    .D(_09305_),
    .Y(_09306_));
 sky130_fd_sc_hd__or2_1 _28728_ (.A(\inst$top.soc.cpu.loadstore.dbus__adr[29] ),
    .B(net2555),
    .X(_09307_));
 sky130_fd_sc_hd__o21a_1 _28729_ (.A1(net2558),
    .A2(\inst$top.soc.cpu.fetch.ibus__adr[29] ),
    .B1(_09307_),
    .X(_09308_));
 sky130_fd_sc_hd__nand2_1 _28730_ (.A(net2557),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[28] ),
    .Y(_09309_));
 sky130_fd_sc_hd__nand2_1 _28731_ (.A(net2561),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[28] ),
    .Y(_09310_));
 sky130_fd_sc_hd__nand2_1 _28732_ (.A(_09309_),
    .B(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__nand2_1 _28733_ (.A(net2556),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[13] ),
    .Y(_09312_));
 sky130_fd_sc_hd__nand2_1 _28734_ (.A(net2560),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[13] ),
    .Y(_09313_));
 sky130_fd_sc_hd__nand2_1 _28735_ (.A(_09312_),
    .B(_09313_),
    .Y(_09314_));
 sky130_fd_sc_hd__or2_2 _28736_ (.A(\inst$top.soc.cpu.loadstore.dbus__adr[10] ),
    .B(net2555),
    .X(_09315_));
 sky130_fd_sc_hd__o21ai_0 _28737_ (.A1(net2559),
    .A2(\inst$top.soc.cpu.fetch.ibus__adr[10] ),
    .B1(_09315_),
    .Y(_09316_));
 sky130_fd_sc_hd__inv_1 _28738_ (.A(_09316_),
    .Y(_09317_));
 sky130_fd_sc_hd__nor2_1 _28739_ (.A(_09314_),
    .B(_09317_),
    .Y(_09318_));
 sky130_fd_sc_hd__nand2_1 _28740_ (.A(net2556),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[11] ),
    .Y(_09319_));
 sky130_fd_sc_hd__nand2_1 _28741_ (.A(net2560),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[11] ),
    .Y(_09320_));
 sky130_fd_sc_hd__nand2_1 _28742_ (.A(_09319_),
    .B(_09320_),
    .Y(_09321_));
 sky130_fd_sc_hd__nand2_1 _28743_ (.A(net2556),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[12] ),
    .Y(_09322_));
 sky130_fd_sc_hd__nand2_1 _28744_ (.A(net2560),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[12] ),
    .Y(_09323_));
 sky130_fd_sc_hd__nand2_1 _28745_ (.A(_09322_),
    .B(_09323_),
    .Y(_09324_));
 sky130_fd_sc_hd__nor2_1 _28746_ (.A(_09321_),
    .B(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__nand2_1 _28747_ (.A(_09318_),
    .B(_09325_),
    .Y(_09326_));
 sky130_fd_sc_hd__nand2_1 _28748_ (.A(net2555),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[16] ),
    .Y(_09327_));
 sky130_fd_sc_hd__nand2_1 _28749_ (.A(net2558),
    .B(\inst$top.soc.cpu.loadstore.dbus__adr[16] ),
    .Y(_09328_));
 sky130_fd_sc_hd__nand2_1 _28750_ (.A(_09327_),
    .B(_09328_),
    .Y(_09329_));
 sky130_fd_sc_hd__mux2i_1 _28751_ (.A0(\inst$top.soc.cpu.fetch.ibus__adr[17] ),
    .A1(\inst$top.soc.cpu.loadstore.dbus__adr[17] ),
    .S(net2558),
    .Y(_09330_));
 sky130_fd_sc_hd__inv_1 _28752_ (.A(_09330_),
    .Y(_09331_));
 sky130_fd_sc_hd__nor2_1 _28753_ (.A(_09329_),
    .B(_09331_),
    .Y(_09332_));
 sky130_fd_sc_hd__inv_1 _28754_ (.A(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__nor4_1 _28755_ (.A(_09308_),
    .B(_09311_),
    .C(_09326_),
    .D(_09333_),
    .Y(_09334_));
 sky130_fd_sc_hd__nand2_1 _28756_ (.A(_09306_),
    .B(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__inv_1 _28757_ (.A(_09335_),
    .Y(_09336_));
 sky130_fd_sc_hd__inv_1 _28758_ (.A(\inst$top.soc.sram.wb_bus__ack ),
    .Y(_09337_));
 sky130_fd_sc_hd__nand2_1 _28759_ (.A(\inst$top.soc.cpu.loadstore.dbus__cyc ),
    .B(net2561),
    .Y(_09338_));
 sky130_fd_sc_hd__inv_1 _28760_ (.A(_09338_),
    .Y(_09339_));
 sky130_fd_sc_hd__inv_1 _28761_ (.A(\inst$top.soc.cpu.fetch.ibus__cyc ),
    .Y(_09340_));
 sky130_fd_sc_hd__nor2_1 _28762_ (.A(net2564),
    .B(_09340_),
    .Y(_09341_));
 sky130_fd_sc_hd__nand2_1 _28763_ (.A(net2557),
    .B(\inst$top.soc.cpu.fetch.ibus__stb ),
    .Y(_09342_));
 sky130_fd_sc_hd__nand2_1 _28764_ (.A(net2564),
    .B(\inst$top.soc.cpu.loadstore.dbus__stb ),
    .Y(_09343_));
 sky130_fd_sc_hd__nand2_1 _28765_ (.A(_09342_),
    .B(_09343_),
    .Y(_09344_));
 sky130_fd_sc_hd__o21ai_0 _28766_ (.A1(_09339_),
    .A2(_09341_),
    .B1(_09344_),
    .Y(_09345_));
 sky130_fd_sc_hd__inv_1 _28767_ (.A(_09345_),
    .Y(_09346_));
 sky130_fd_sc_hd__nand3_1 _28768_ (.A(_09336_),
    .B(_09337_),
    .C(_09346_),
    .Y(_09347_));
 sky130_fd_sc_hd__nor2_1 _28769_ (.A(_09256_),
    .B(_09347_),
    .Y(_09348_));
 sky130_fd_sc_hd__inv_2 _28770_ (.A(_09348_),
    .Y(\inst$top.soc.sram.read_port__en ));
 sky130_fd_sc_hd__nor2_4 _28771_ (.A(_09255_),
    .B(\inst$top.soc.sram.read_port__en ),
    .Y(\inst$top.soc.sram.write_port__en[1] ));
 sky130_fd_sc_hd__inv_1 _28772_ (.A(\inst$top.soc.cpu.loadstore.dbus__sel[0] ),
    .Y(_09349_));
 sky130_fd_sc_hd__nor2_4 _28773_ (.A(_09349_),
    .B(\inst$top.soc.sram.read_port__en ),
    .Y(\inst$top.soc.sram.write_port__en[0] ));
 sky130_fd_sc_hd__inv_1 _28774_ (.A(\inst$top.soc.cpu.loadstore.dbus__sel[3] ),
    .Y(_09350_));
 sky130_fd_sc_hd__nor2_4 _28775_ (.A(_09350_),
    .B(\inst$top.soc.sram.read_port__en ),
    .Y(\inst$top.soc.sram.write_port__en[3] ));
 sky130_fd_sc_hd__inv_1 _28776_ (.A(\inst$top.soc.cpu.loadstore.dbus__sel[2] ),
    .Y(_09351_));
 sky130_fd_sc_hd__nor2_4 _28777_ (.A(_09351_),
    .B(\inst$top.soc.sram.read_port__en ),
    .Y(\inst$top.soc.sram.write_port__en[2] ));
 sky130_fd_sc_hd__nor4_2 _28778_ (.A(net761),
    .B(net760),
    .C(net759),
    .D(net757),
    .Y(_00161_));
 sky130_fd_sc_hd__inv_2 _28779_ (.A(net1683),
    .Y(_09352_));
 sky130_fd_sc_hd__inv_2 _28781_ (.A(\inst$top.soc.cpu.multiplier.x_prod[0] ),
    .Y(_00162_));
 sky130_fd_sc_hd__nand2_1 _28782_ (.A(net1153),
    .B(net1077),
    .Y(_00172_));
 sky130_fd_sc_hd__nand2_1 _28783_ (.A(net1153),
    .B(net1394),
    .Y(_00181_));
 sky130_fd_sc_hd__nand2_1 _28784_ (.A(net1251),
    .B(net1351),
    .Y(_00184_));
 sky130_fd_sc_hd__nand2_1 _28785_ (.A(net1356),
    .B(net1251),
    .Y(_00190_));
 sky130_fd_sc_hd__nand2_1 _28786_ (.A(net1361),
    .B(net1251),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _28787_ (.A(net1155),
    .B(net1251),
    .Y(_00205_));
 sky130_fd_sc_hd__inv_2 _28788_ (.A(_03390_),
    .Y(_00263_));
 sky130_fd_sc_hd__inv_2 _28789_ (.A(_03397_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _28790_ (.A(net1355),
    .B(net1398),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _28791_ (.A(net1258),
    .B(net1397),
    .Y(_01069_));
 sky130_fd_sc_hd__nand2_1 _28792_ (.A(net1427),
    .B(net1309),
    .Y(_01183_));
 sky130_fd_sc_hd__nand2_1 _28793_ (.A(net1428),
    .B(net1305),
    .Y(_01301_));
 sky130_fd_sc_hd__inv_2 _28794_ (.A(_01450_),
    .Y(_01392_));
 sky130_fd_sc_hd__nand2_1 _28795_ (.A(_06033_),
    .B(net1396),
    .Y(_01620_));
 sky130_fd_sc_hd__inv_2 _28796_ (.A(_01769_),
    .Y(_01718_));
 sky130_fd_sc_hd__nand2_1 _28797_ (.A(net1459),
    .B(net1425),
    .Y(_01912_));
 sky130_fd_sc_hd__nand2_1 _28798_ (.A(net1273),
    .B(net1726),
    .Y(_02128_));
 sky130_fd_sc_hd__inv_2 _28799_ (.A(_02171_),
    .Y(_02138_));
 sky130_fd_sc_hd__nand2_1 _28800_ (.A(net1253),
    .B(net1216),
    .Y(_02194_));
 sky130_fd_sc_hd__nand2_1 _28801_ (.A(net1253),
    .B(net1457),
    .Y(_02322_));
 sky130_fd_sc_hd__inv_2 _28802_ (.A(_02366_),
    .Y(_02333_));
 sky130_fd_sc_hd__inv_2 _28803_ (.A(_02445_),
    .Y(_02419_));
 sky130_fd_sc_hd__nand2_1 _28804_ (.A(net1467),
    .B(net1480),
    .Y(_02477_));
 sky130_fd_sc_hd__inv_2 _28805_ (.A(_02497_),
    .Y(_02481_));
 sky130_fd_sc_hd__nand2_1 _28806_ (.A(_06033_),
    .B(net1473),
    .Y(_02511_));
 sky130_fd_sc_hd__nand2_1 _28807_ (.A(net1077),
    .B(net1262),
    .Y(_00182_));
 sky130_fd_sc_hd__nand2_1 _28808_ (.A(net1356),
    .B(net1385),
    .Y(_00185_));
 sky130_fd_sc_hd__inv_2 _28809_ (.A(_03365_),
    .Y(_00189_));
 sky130_fd_sc_hd__nand2_1 _28810_ (.A(net1361),
    .B(net1385),
    .Y(_00191_));
 sky130_fd_sc_hd__nand2_1 _28811_ (.A(net1155),
    .B(net1385),
    .Y(_00195_));
 sky130_fd_sc_hd__inv_2 _28812_ (.A(_03370_),
    .Y(_00198_));
 sky130_fd_sc_hd__inv_2 _28813_ (.A(_03374_),
    .Y(_00201_));
 sky130_fd_sc_hd__nand2_1 _28814_ (.A(_03082_),
    .B(net1389),
    .Y(_00206_));
 sky130_fd_sc_hd__inv_2 _28815_ (.A(_03391_),
    .Y(_00264_));
 sky130_fd_sc_hd__inv_2 _28816_ (.A(_03398_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _28817_ (.A(net1203),
    .B(net1262),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_1 _28818_ (.A(net1153),
    .B(net1203),
    .Y(_00320_));
 sky130_fd_sc_hd__nand2_1 _28819_ (.A(net1362),
    .B(net1203),
    .Y(_00347_));
 sky130_fd_sc_hd__nand2_1 _28820_ (.A(net1356),
    .B(net1203),
    .Y(_00384_));
 sky130_fd_sc_hd__inv_2 _28821_ (.A(_03423_),
    .Y(_00386_));
 sky130_fd_sc_hd__nand2_1 _28822_ (.A(net1341),
    .B(net1398),
    .Y(_00429_));
 sky130_fd_sc_hd__inv_2 _28823_ (.A(_03430_),
    .Y(_00451_));
 sky130_fd_sc_hd__nand2_1 _28824_ (.A(net1337),
    .B(net1398),
    .Y(_00463_));
 sky130_fd_sc_hd__nand2_1 _28825_ (.A(net1077),
    .B(net1322),
    .Y(_00467_));
 sky130_fd_sc_hd__inv_2 _28826_ (.A(_03438_),
    .Y(_00480_));
 sky130_fd_sc_hd__nand2_1 _28827_ (.A(net1077),
    .B(net1316),
    .Y(_00503_));
 sky130_fd_sc_hd__nand2_1 _28828_ (.A(net1076),
    .B(net1311),
    .Y(_00545_));
 sky130_fd_sc_hd__nand2_1 _28829_ (.A(net1427),
    .B(net1365),
    .Y(_00567_));
 sky130_fd_sc_hd__nand2_1 _28830_ (.A(net1076),
    .B(net1307),
    .Y(_00588_));
 sky130_fd_sc_hd__nand2_1 _28831_ (.A(net1335),
    .B(net1410),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _28832_ (.A(net1075),
    .B(net1302),
    .Y(_00638_));
 sky130_fd_sc_hd__nand2_1 _28833_ (.A(net1075),
    .B(net1296),
    .Y(_00686_));
 sky130_fd_sc_hd__nand2_1 _28834_ (.A(net1206),
    .B(net1321),
    .Y(_00721_));
 sky130_fd_sc_hd__nand2_1 _28835_ (.A(net1075),
    .B(net1294),
    .Y(_00736_));
 sky130_fd_sc_hd__inv_2 _28836_ (.A(_03501_),
    .Y(_00749_));
 sky130_fd_sc_hd__inv_2 _28837_ (.A(_03511_),
    .Y(_00765_));
 sky130_fd_sc_hd__nand2_1 _28838_ (.A(net1075),
    .B(net1288),
    .Y(_00790_));
 sky130_fd_sc_hd__nand2_1 _28839_ (.A(net1074),
    .B(net1283),
    .Y(_00844_));
 sky130_fd_sc_hd__nand2_1 _28840_ (.A(net1074),
    .B(net1278),
    .Y(_00901_));
 sky130_fd_sc_hd__nand2_1 _28841_ (.A(net1320),
    .B(net1422),
    .Y(_00939_));
 sky130_fd_sc_hd__nand2_1 _28842_ (.A(net1258),
    .B(net1073),
    .Y(_00956_));
 sky130_fd_sc_hd__nand2_1 _28843_ (.A(net1154),
    .B(net1723),
    .Y(_00980_));
 sky130_fd_sc_hd__nand2_1 _28844_ (.A(net1073),
    .B(net1273),
    .Y(_01016_));
 sky130_fd_sc_hd__nand2_1 _28845_ (.A(net1306),
    .B(net1418),
    .Y(_01061_));
 sky130_fd_sc_hd__nand2_1 _28846_ (.A(net1293),
    .B(net1205),
    .Y(_01064_));
 sky130_fd_sc_hd__nand2_1 _28847_ (.A(net1398),
    .B(net1278),
    .Y(_01070_));
 sky130_fd_sc_hd__inv_2 _28848_ (.A(_03589_),
    .Y(_01115_));
 sky130_fd_sc_hd__nand2_1 _28849_ (.A(net1287),
    .B(net1204),
    .Y(_01128_));
 sky130_fd_sc_hd__nand2_1 _28850_ (.A(net1204),
    .B(net1283),
    .Y(_01191_));
 sky130_fd_sc_hd__nand2_1 _28851_ (.A(net1204),
    .B(net1279),
    .Y(_01253_));
 sky130_fd_sc_hd__nand2_1 _28852_ (.A(net1408),
    .B(net1279),
    .Y(_01309_));
 sky130_fd_sc_hd__nand2_1 _28853_ (.A(net1274),
    .B(net1204),
    .Y(_01377_));
 sky130_fd_sc_hd__nand2_1 _28854_ (.A(net1427),
    .B(net1294),
    .Y(_01426_));
 sky130_fd_sc_hd__nand2_1 _28855_ (.A(net1205),
    .B(net1270),
    .Y(_01434_));
 sky130_fd_sc_hd__nand2_1 _28856_ (.A(net1255),
    .B(net1205),
    .Y(_01494_));
 sky130_fd_sc_hd__nand2_1 _28857_ (.A(net1252),
    .B(net1204),
    .Y(_01554_));
 sky130_fd_sc_hd__nand2_1 _28858_ (.A(net1452),
    .B(net1204),
    .Y(_01610_));
 sky130_fd_sc_hd__nand2_1 _28859_ (.A(net1132),
    .B(net1293),
    .Y(_01650_));
 sky130_fd_sc_hd__nand2_1 _28860_ (.A(net1459),
    .B(net1204),
    .Y(_01663_));
 sky130_fd_sc_hd__nand2_1 _28861_ (.A(net1466),
    .B(net1204),
    .Y(_01715_));
 sky130_fd_sc_hd__nand2_1 _28862_ (.A(net1432),
    .B(net1279),
    .Y(_01752_));
 sky130_fd_sc_hd__nand2_1 _28863_ (.A(net1477),
    .B(net1204),
    .Y(_01765_));
 sky130_fd_sc_hd__nand2_1 _28864_ (.A(net1270),
    .B(net1433),
    .Y(_01908_));
 sky130_fd_sc_hd__nand2_1 _28865_ (.A(net1427),
    .B(net1452),
    .Y(_01913_));
 sky130_fd_sc_hd__nand2_1 _28866_ (.A(net1446),
    .B(net1278),
    .Y(_01956_));
 sky130_fd_sc_hd__nand2_1 _28867_ (.A(net1255),
    .B(net1433),
    .Y(_01960_));
 sky130_fd_sc_hd__inv_2 _28868_ (.A(_01771_),
    .Y(_01772_));
 sky130_fd_sc_hd__nand2_1 _28869_ (.A(net1273),
    .B(net1442),
    .Y(_02004_));
 sky130_fd_sc_hd__nand2_1 _28870_ (.A(net1252),
    .B(net1434),
    .Y(_02007_));
 sky130_fd_sc_hd__nand2_1 _28871_ (.A(net1271),
    .B(net1442),
    .Y(_02051_));
 sky130_fd_sc_hd__nand2_1 _28872_ (.A(net1452),
    .B(net1434),
    .Y(_02055_));
 sky130_fd_sc_hd__nand2_1 _28873_ (.A(net1255),
    .B(net1442),
    .Y(_02097_));
 sky130_fd_sc_hd__nand2_1 _28874_ (.A(net1459),
    .B(net1434),
    .Y(_02100_));
 sky130_fd_sc_hd__nand2_1 _28875_ (.A(net1252),
    .B(net1442),
    .Y(_02133_));
 sky130_fd_sc_hd__nand2_1 _28876_ (.A(net1466),
    .B(net1434),
    .Y(_02136_));
 sky130_fd_sc_hd__nand2_1 _28877_ (.A(net1452),
    .B(net1442),
    .Y(_02165_));
 sky130_fd_sc_hd__nand2_1 _28878_ (.A(net1477),
    .B(net1434),
    .Y(_02168_));
 sky130_fd_sc_hd__nand2_1 _28879_ (.A(net1730),
    .B(net1272),
    .Y(_02195_));
 sky130_fd_sc_hd__nand2_1 _28880_ (.A(net1459),
    .B(net1443),
    .Y(_02199_));
 sky130_fd_sc_hd__nand2_1 _28881_ (.A(net1481),
    .B(net1434),
    .Y(_02202_));
 sky130_fd_sc_hd__inv_2 _28882_ (.A(_02309_),
    .Y(_02311_));
 sky130_fd_sc_hd__inv_2 _28883_ (.A(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hd__nand2_1 _28884_ (.A(net1045),
    .B(net1110),
    .Y(_02512_));
 sky130_fd_sc_hd__inv_2 _28885_ (.A(_02397_),
    .Y(_02424_));
 sky130_fd_sc_hd__inv_2 _28886_ (.A(_03072_),
    .Y(_00174_));
 sky130_fd_sc_hd__nand2_1 _28887_ (.A(net1361),
    .B(net1389),
    .Y(_00186_));
 sky130_fd_sc_hd__inv_2 _28888_ (.A(_03078_),
    .Y(_00192_));
 sky130_fd_sc_hd__nand2_1 _28889_ (.A(net1262),
    .B(net1389),
    .Y(_00196_));
 sky130_fd_sc_hd__inv_2 _28890_ (.A(_03081_),
    .Y(_00207_));
 sky130_fd_sc_hd__nand2_1 _28891_ (.A(_03082_),
    .B(net1411),
    .Y(_00296_));
 sky130_fd_sc_hd__nand2_1 _28892_ (.A(net1262),
    .B(net1411),
    .Y(_00321_));
 sky130_fd_sc_hd__inv_2 _28893_ (.A(_03056_),
    .Y(_00325_));
 sky130_fd_sc_hd__nand2_1 _28894_ (.A(net1153),
    .B(net1411),
    .Y(_00348_));
 sky130_fd_sc_hd__nand2_1 _28895_ (.A(net1362),
    .B(net1411),
    .Y(_00385_));
 sky130_fd_sc_hd__inv_2 _28896_ (.A(_00382_),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _28897_ (.A(_03045_),
    .B(net1346),
    .Y(_00430_));
 sky130_fd_sc_hd__inv_2 _28898_ (.A(_03439_),
    .Y(_00452_));
 sky130_fd_sc_hd__inv_2 _28899_ (.A(_00465_),
    .Y(_00464_));
 sky130_fd_sc_hd__nand2_1 _28900_ (.A(net1327),
    .B(net1396),
    .Y(_00468_));
 sky130_fd_sc_hd__inv_2 _28901_ (.A(_03450_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_1 _28902_ (.A(net1321),
    .B(net1396),
    .Y(_00504_));
 sky130_fd_sc_hd__inv_2 _28903_ (.A(_03447_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_1 _28904_ (.A(net1316),
    .B(net1395),
    .Y(_00546_));
 sky130_fd_sc_hd__inv_2 _28905_ (.A(_03457_),
    .Y(_00555_));
 sky130_fd_sc_hd__nand2_1 _28906_ (.A(net1428),
    .B(net1155),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _28907_ (.A(net1311),
    .B(net1395),
    .Y(_00589_));
 sky130_fd_sc_hd__inv_2 _28908_ (.A(_03465_),
    .Y(_00598_));
 sky130_fd_sc_hd__inv_2 _28909_ (.A(_03035_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand2_1 _28910_ (.A(net1307),
    .B(net1395),
    .Y(_00639_));
 sky130_fd_sc_hd__inv_2 _28911_ (.A(_03480_),
    .Y(_00648_));
 sky130_fd_sc_hd__nand2_1 _28912_ (.A(net1302),
    .B(net1395),
    .Y(_00687_));
 sky130_fd_sc_hd__inv_2 _28913_ (.A(_03488_),
    .Y(_00696_));
 sky130_fd_sc_hd__inv_2 _28914_ (.A(_03029_),
    .Y(_00722_));
 sky130_fd_sc_hd__nand2_1 _28915_ (.A(net1296),
    .B(net1395),
    .Y(_00737_));
 sky130_fd_sc_hd__inv_2 _28916_ (.A(_03500_),
    .Y(_00747_));
 sky130_fd_sc_hd__inv_2 _28917_ (.A(_03515_),
    .Y(_00750_));
 sky130_fd_sc_hd__inv_2 _28918_ (.A(_00761_),
    .Y(_00766_));
 sky130_fd_sc_hd__nand2_1 _28919_ (.A(net1292),
    .B(net1395),
    .Y(_00791_));
 sky130_fd_sc_hd__nand2_1 _28920_ (.A(net1288),
    .B(net1395),
    .Y(_00845_));
 sky130_fd_sc_hd__nand2_1 _28921_ (.A(net1396),
    .B(net1283),
    .Y(_00902_));
 sky130_fd_sc_hd__inv_2 _28922_ (.A(_03015_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand2_1 _28923_ (.A(net1395),
    .B(net1278),
    .Y(_00957_));
 sky130_fd_sc_hd__nand2_1 _28924_ (.A(net1727),
    .B(net1263),
    .Y(_00981_));
 sky130_fd_sc_hd__nand2_1 _28925_ (.A(net1258),
    .B(net1395),
    .Y(_01017_));
 sky130_fd_sc_hd__inv_2 _28926_ (.A(_03009_),
    .Y(_01062_));
 sky130_fd_sc_hd__nand2_1 _28927_ (.A(net1297),
    .B(net1409),
    .Y(_01065_));
 sky130_fd_sc_hd__inv_2 _28928_ (.A(_03598_),
    .Y(_01116_));
 sky130_fd_sc_hd__nand2_1 _28929_ (.A(net1293),
    .B(net1408),
    .Y(_01129_));
 sky130_fd_sc_hd__inv_2 _28930_ (.A(_03006_),
    .Y(_01185_));
 sky130_fd_sc_hd__nand2_1 _28931_ (.A(net1287),
    .B(net1408),
    .Y(_01192_));
 sky130_fd_sc_hd__nand2_1 _28932_ (.A(net1284),
    .B(net1408),
    .Y(_01254_));
 sky130_fd_sc_hd__inv_2 _28933_ (.A(_03000_),
    .Y(_01303_));
 sky130_fd_sc_hd__nand2_1 _28934_ (.A(net1284),
    .B(net1412),
    .Y(_01310_));
 sky130_fd_sc_hd__nand2_1 _28935_ (.A(net1258),
    .B(net1408),
    .Y(_01378_));
 sky130_fd_sc_hd__inv_2 _28936_ (.A(_01341_),
    .Y(_01394_));
 sky130_fd_sc_hd__inv_2 _28937_ (.A(_01428_),
    .Y(_01427_));
 sky130_fd_sc_hd__nand2_1 _28938_ (.A(net1273),
    .B(net1409),
    .Y(_01435_));
 sky130_fd_sc_hd__nand2_1 _28939_ (.A(net1270),
    .B(net1409),
    .Y(_01495_));
 sky130_fd_sc_hd__nand2_1 _28940_ (.A(net1255),
    .B(net1408),
    .Y(_01555_));
 sky130_fd_sc_hd__nand2_1 _28941_ (.A(net1252),
    .B(net1408),
    .Y(_01611_));
 sky130_fd_sc_hd__inv_2 _28942_ (.A(_01504_),
    .Y(_01622_));
 sky130_fd_sc_hd__inv_2 _28943_ (.A(_02981_),
    .Y(_01651_));
 sky130_fd_sc_hd__nand2_1 _28944_ (.A(net1452),
    .B(net1408),
    .Y(_01664_));
 sky130_fd_sc_hd__nand2_1 _28945_ (.A(net1459),
    .B(net1408),
    .Y(_01716_));
 sky130_fd_sc_hd__inv_2 _28946_ (.A(_01666_),
    .Y(_01720_));
 sky130_fd_sc_hd__inv_2 _28947_ (.A(_01451_),
    .Y(_01511_));
 sky130_fd_sc_hd__inv_2 _28948_ (.A(_02555_),
    .Y(_01753_));
 sky130_fd_sc_hd__nand2_1 _28949_ (.A(net1466),
    .B(net1408),
    .Y(_01766_));
 sky130_fd_sc_hd__nand2_1 _28950_ (.A(net1133),
    .B(net1273),
    .Y(_01909_));
 sky130_fd_sc_hd__inv_2 _28951_ (.A(_01958_),
    .Y(_01957_));
 sky130_fd_sc_hd__nand2_1 _28952_ (.A(net1133),
    .B(net1270),
    .Y(_01961_));
 sky130_fd_sc_hd__inv_2 _28953_ (.A(_01770_),
    .Y(_01820_));
 sky130_fd_sc_hd__nand2_1 _28954_ (.A(net1258),
    .B(net1446),
    .Y(_02005_));
 sky130_fd_sc_hd__nand2_1 _28955_ (.A(net1255),
    .B(net1134),
    .Y(_02008_));
 sky130_fd_sc_hd__inv_2 _28956_ (.A(_02053_),
    .Y(_02052_));
 sky130_fd_sc_hd__nand2_1 _28957_ (.A(net1252),
    .B(net1134),
    .Y(_02056_));
 sky130_fd_sc_hd__inv_2 _28958_ (.A(_01969_),
    .Y(_02018_));
 sky130_fd_sc_hd__nand2_1 _28959_ (.A(net1271),
    .B(net1446),
    .Y(_02098_));
 sky130_fd_sc_hd__nand2_1 _28960_ (.A(net1134),
    .B(net1452),
    .Y(_02101_));
 sky130_fd_sc_hd__inv_2 _28961_ (.A(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__inv_2 _28962_ (.A(_02603_),
    .Y(_02130_));
 sky130_fd_sc_hd__nand2_1 _28963_ (.A(net1255),
    .B(net1446),
    .Y(_02134_));
 sky130_fd_sc_hd__nand2_1 _28964_ (.A(net1459),
    .B(net1134),
    .Y(_02137_));
 sky130_fd_sc_hd__inv_2 _28965_ (.A(_02102_),
    .Y(_02140_));
 sky130_fd_sc_hd__nand2_1 _28966_ (.A(net1252),
    .B(net1446),
    .Y(_02166_));
 sky130_fd_sc_hd__nand2_1 _28967_ (.A(net1466),
    .B(net1134),
    .Y(_02169_));
 sky130_fd_sc_hd__inv_2 _28968_ (.A(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__nand2_1 _28969_ (.A(net1452),
    .B(net1447),
    .Y(_02200_));
 sky130_fd_sc_hd__nand2_1 _28970_ (.A(net1134),
    .B(net1476),
    .Y(_02203_));
 sky130_fd_sc_hd__inv_2 _28971_ (.A(_02641_),
    .Y(_02324_));
 sky130_fd_sc_hd__inv_2 _28972_ (.A(_02302_),
    .Y(_02335_));
 sky130_fd_sc_hd__inv_2 _28973_ (.A(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__inv_2 _28974_ (.A(_02269_),
    .Y(_02270_));
 sky130_fd_sc_hd__inv_2 _28975_ (.A(_02389_),
    .Y(_02421_));
 sky130_fd_sc_hd__inv_2 _28976_ (.A(_02678_),
    .Y(_02479_));
 sky130_fd_sc_hd__inv_2 _28977_ (.A(_02461_),
    .Y(_02483_));
 sky130_fd_sc_hd__inv_2 _28978_ (.A(_02691_),
    .Y(_02513_));
 sky130_fd_sc_hd__inv_2 _28979_ (.A(_00859_),
    .Y(_00860_));
 sky130_fd_sc_hd__inv_2 _28980_ (.A(_00916_),
    .Y(_00917_));
 sky130_fd_sc_hd__inv_2 _28981_ (.A(_00971_),
    .Y(_00972_));
 sky130_fd_sc_hd__inv_2 _28982_ (.A(_01031_),
    .Y(_01032_));
 sky130_fd_sc_hd__inv_2 _28983_ (.A(_01092_),
    .Y(_01093_));
 sky130_fd_sc_hd__inv_2 _28984_ (.A(_01158_),
    .Y(_01159_));
 sky130_fd_sc_hd__inv_2 _28985_ (.A(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__inv_2 _28986_ (.A(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__inv_2 _28987_ (.A(_01404_),
    .Y(_01405_));
 sky130_fd_sc_hd__inv_2 _28988_ (.A(_01462_),
    .Y(_01463_));
 sky130_fd_sc_hd__inv_2 _28989_ (.A(_01518_),
    .Y(_01519_));
 sky130_fd_sc_hd__inv_2 _28990_ (.A(_01576_),
    .Y(_01577_));
 sky130_fd_sc_hd__inv_2 _28991_ (.A(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__inv_2 _28992_ (.A(_01682_),
    .Y(_01683_));
 sky130_fd_sc_hd__inv_2 _28993_ (.A(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__inv_2 _28994_ (.A(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__inv_2 _28995_ (.A(_02066_),
    .Y(_02068_));
 sky130_fd_sc_hd__inv_2 _28996_ (.A(_02527_),
    .Y(_02528_));
 sky130_fd_sc_hd__inv_2 _28997_ (.A(_00179_),
    .Y(_00180_));
 sky130_fd_sc_hd__inv_2 _28998_ (.A(_00214_),
    .Y(_00221_));
 sky130_fd_sc_hd__inv_2 _28999_ (.A(_00219_),
    .Y(_00220_));
 sky130_fd_sc_hd__inv_2 _29000_ (.A(_00232_),
    .Y(_00240_));
 sky130_fd_sc_hd__inv_2 _29001_ (.A(_00237_),
    .Y(_00238_));
 sky130_fd_sc_hd__inv_2 _29002_ (.A(_00251_),
    .Y(_00259_));
 sky130_fd_sc_hd__inv_2 _29003_ (.A(_00256_),
    .Y(_00257_));
 sky130_fd_sc_hd__inv_2 _29004_ (.A(_00275_),
    .Y(_00283_));
 sky130_fd_sc_hd__inv_2 _29005_ (.A(_00280_),
    .Y(_00281_));
 sky130_fd_sc_hd__inv_2 _29006_ (.A(_00288_),
    .Y(_00291_));
 sky130_fd_sc_hd__inv_2 _29007_ (.A(_00306_),
    .Y(_00314_));
 sky130_fd_sc_hd__inv_2 _29008_ (.A(_00311_),
    .Y(_00312_));
 sky130_fd_sc_hd__inv_2 _29009_ (.A(_00333_),
    .Y(_00341_));
 sky130_fd_sc_hd__inv_2 _29010_ (.A(_00338_),
    .Y(_00339_));
 sky130_fd_sc_hd__inv_2 _29011_ (.A(_00354_),
    .Y(_00355_));
 sky130_fd_sc_hd__inv_2 _29012_ (.A(_00365_),
    .Y(_00373_));
 sky130_fd_sc_hd__inv_2 _29013_ (.A(_00370_),
    .Y(_00371_));
 sky130_fd_sc_hd__inv_2 _29014_ (.A(_00393_),
    .Y(_00395_));
 sky130_fd_sc_hd__inv_2 _29015_ (.A(_00400_),
    .Y(_00417_));
 sky130_fd_sc_hd__inv_2 _29016_ (.A(_00405_),
    .Y(_00413_));
 sky130_fd_sc_hd__inv_2 _29017_ (.A(_00410_),
    .Y(_00411_));
 sky130_fd_sc_hd__inv_2 _29018_ (.A(_00436_),
    .Y(_00444_));
 sky130_fd_sc_hd__inv_2 _29019_ (.A(_00441_),
    .Y(_00442_));
 sky130_fd_sc_hd__inv_2 _29020_ (.A(_00473_),
    .Y(_00474_));
 sky130_fd_sc_hd__inv_2 _29021_ (.A(_00500_),
    .Y(_00501_));
 sky130_fd_sc_hd__inv_2 _29022_ (.A(_00509_),
    .Y(_00510_));
 sky130_fd_sc_hd__inv_2 _29023_ (.A(_00517_),
    .Y(_00519_));
 sky130_fd_sc_hd__inv_2 _29024_ (.A(_00533_),
    .Y(_00534_));
 sky130_fd_sc_hd__inv_2 _29025_ (.A(_00541_),
    .Y(_00543_));
 sky130_fd_sc_hd__inv_2 _29026_ (.A(_00551_),
    .Y(_00552_));
 sky130_fd_sc_hd__inv_2 _29027_ (.A(_00583_),
    .Y(_00585_));
 sky130_fd_sc_hd__inv_2 _29028_ (.A(_00594_),
    .Y(_00595_));
 sky130_fd_sc_hd__inv_2 _29029_ (.A(_00603_),
    .Y(_00606_));
 sky130_fd_sc_hd__inv_2 _29030_ (.A(_00634_),
    .Y(_00636_));
 sky130_fd_sc_hd__inv_2 _29031_ (.A(_00644_),
    .Y(_00645_));
 sky130_fd_sc_hd__inv_2 _29032_ (.A(_00653_),
    .Y(_00656_));
 sky130_fd_sc_hd__inv_2 _29033_ (.A(_00682_),
    .Y(_00684_));
 sky130_fd_sc_hd__inv_2 _29034_ (.A(_00692_),
    .Y(_00693_));
 sky130_fd_sc_hd__inv_2 _29035_ (.A(_00701_),
    .Y(_00704_));
 sky130_fd_sc_hd__inv_2 _29036_ (.A(_00732_),
    .Y(_00734_));
 sky130_fd_sc_hd__inv_2 _29037_ (.A(_00742_),
    .Y(_00743_));
 sky130_fd_sc_hd__inv_2 _29038_ (.A(_00786_),
    .Y(_00788_));
 sky130_fd_sc_hd__inv_2 _29039_ (.A(_00796_),
    .Y(_00797_));
 sky130_fd_sc_hd__inv_2 _29040_ (.A(_00805_),
    .Y(_00807_));
 sky130_fd_sc_hd__inv_2 _29041_ (.A(_00828_),
    .Y(_00832_));
 sky130_fd_sc_hd__inv_2 _29042_ (.A(_00840_),
    .Y(_00842_));
 sky130_fd_sc_hd__inv_2 _29043_ (.A(_00850_),
    .Y(_00851_));
 sky130_fd_sc_hd__inv_2 _29044_ (.A(_00892_),
    .Y(_00919_));
 sky130_fd_sc_hd__inv_2 _29045_ (.A(_00897_),
    .Y(_00899_));
 sky130_fd_sc_hd__inv_2 _29046_ (.A(_00907_),
    .Y(_00908_));
 sky130_fd_sc_hd__inv_2 _29047_ (.A(_00952_),
    .Y(_00954_));
 sky130_fd_sc_hd__inv_2 _29048_ (.A(_00962_),
    .Y(_00963_));
 sky130_fd_sc_hd__inv_2 _29049_ (.A(_00996_),
    .Y(_00997_));
 sky130_fd_sc_hd__inv_2 _29050_ (.A(_01012_),
    .Y(_01014_));
 sky130_fd_sc_hd__inv_2 _29051_ (.A(_01022_),
    .Y(_01023_));
 sky130_fd_sc_hd__inv_2 _29052_ (.A(_01052_),
    .Y(_01068_));
 sky130_fd_sc_hd__inv_2 _29053_ (.A(_01057_),
    .Y(_01059_));
 sky130_fd_sc_hd__inv_2 _29054_ (.A(_01077_),
    .Y(_01084_));
 sky130_fd_sc_hd__inv_2 _29055_ (.A(_01082_),
    .Y(_01083_));
 sky130_fd_sc_hd__inv_2 _29056_ (.A(_01121_),
    .Y(_01123_));
 sky130_fd_sc_hd__inv_2 _29057_ (.A(_01136_),
    .Y(_01137_));
 sky130_fd_sc_hd__inv_2 _29058_ (.A(_01142_),
    .Y(_01150_));
 sky130_fd_sc_hd__inv_2 _29059_ (.A(_01147_),
    .Y(_01148_));
 sky130_fd_sc_hd__inv_2 _29060_ (.A(_01182_),
    .Y(_01193_));
 sky130_fd_sc_hd__inv_2 _29061_ (.A(_01198_),
    .Y(_01200_));
 sky130_fd_sc_hd__inv_2 _29062_ (.A(_01205_),
    .Y(_01213_));
 sky130_fd_sc_hd__inv_2 _29063_ (.A(_01210_),
    .Y(_01211_));
 sky130_fd_sc_hd__inv_2 _29064_ (.A(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hd__inv_2 _29065_ (.A(_01261_),
    .Y(_01263_));
 sky130_fd_sc_hd__inv_2 _29066_ (.A(_01268_),
    .Y(_01276_));
 sky130_fd_sc_hd__inv_2 _29067_ (.A(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hd__inv_2 _29068_ (.A(_01316_),
    .Y(_01318_));
 sky130_fd_sc_hd__inv_2 _29069_ (.A(_01323_),
    .Y(_01331_));
 sky130_fd_sc_hd__inv_2 _29070_ (.A(_01328_),
    .Y(_01329_));
 sky130_fd_sc_hd__inv_2 _29071_ (.A(_01345_),
    .Y(_01346_));
 sky130_fd_sc_hd__inv_2 _29072_ (.A(_01371_),
    .Y(_01372_));
 sky130_fd_sc_hd__inv_2 _29073_ (.A(_01384_),
    .Y(_01386_));
 sky130_fd_sc_hd__inv_2 _29074_ (.A(_01391_),
    .Y(_01396_));
 sky130_fd_sc_hd__inv_2 _29075_ (.A(_01441_),
    .Y(_01443_));
 sky130_fd_sc_hd__inv_2 _29076_ (.A(_01448_),
    .Y(_01455_));
 sky130_fd_sc_hd__inv_2 _29077_ (.A(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__inv_2 _29078_ (.A(_01488_),
    .Y(_01489_));
 sky130_fd_sc_hd__inv_2 _29079_ (.A(_01501_),
    .Y(_01503_));
 sky130_fd_sc_hd__inv_2 _29080_ (.A(_01508_),
    .Y(_01510_));
 sky130_fd_sc_hd__inv_2 _29081_ (.A(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__inv_2 _29082_ (.A(_01547_),
    .Y(_01549_));
 sky130_fd_sc_hd__inv_2 _29083_ (.A(_01561_),
    .Y(_01563_));
 sky130_fd_sc_hd__inv_2 _29084_ (.A(_01567_),
    .Y(_01569_));
 sky130_fd_sc_hd__inv_2 _29085_ (.A(_01602_),
    .Y(_01604_));
 sky130_fd_sc_hd__inv_2 _29086_ (.A(_01617_),
    .Y(_01619_));
 sky130_fd_sc_hd__inv_2 _29087_ (.A(_01656_),
    .Y(_01658_));
 sky130_fd_sc_hd__inv_2 _29088_ (.A(_01670_),
    .Y(_01672_));
 sky130_fd_sc_hd__inv_2 _29089_ (.A(_01708_),
    .Y(_01710_));
 sky130_fd_sc_hd__inv_2 _29090_ (.A(_01758_),
    .Y(_01760_));
 sky130_fd_sc_hd__inv_2 _29091_ (.A(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__inv_2 _29092_ (.A(_01807_),
    .Y(_01809_));
 sky130_fd_sc_hd__inv_2 _29093_ (.A(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__inv_2 _29094_ (.A(_01827_),
    .Y(_01829_));
 sky130_fd_sc_hd__inv_2 _29095_ (.A(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__inv_2 _29096_ (.A(_01852_),
    .Y(_01856_));
 sky130_fd_sc_hd__inv_2 _29097_ (.A(_01861_),
    .Y(_01863_));
 sky130_fd_sc_hd__inv_2 _29098_ (.A(_01870_),
    .Y(_01871_));
 sky130_fd_sc_hd__inv_2 _29099_ (.A(_01880_),
    .Y(_01882_));
 sky130_fd_sc_hd__inv_2 _29100_ (.A(_01899_),
    .Y(_01901_));
 sky130_fd_sc_hd__inv_2 _29101_ (.A(_01906_),
    .Y(_01911_));
 sky130_fd_sc_hd__inv_2 _29102_ (.A(_01920_),
    .Y(_01924_));
 sky130_fd_sc_hd__inv_2 _29103_ (.A(_01933_),
    .Y(_01935_));
 sky130_fd_sc_hd__inv_2 _29104_ (.A(_01952_),
    .Y(_01954_));
 sky130_fd_sc_hd__inv_2 _29105_ (.A(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__inv_2 _29106_ (.A(_01972_),
    .Y(_01974_));
 sky130_fd_sc_hd__inv_2 _29107_ (.A(_01977_),
    .Y(_02073_));
 sky130_fd_sc_hd__inv_2 _29108_ (.A(_01981_),
    .Y(_01983_));
 sky130_fd_sc_hd__inv_2 _29109_ (.A(_02000_),
    .Y(_02002_));
 sky130_fd_sc_hd__inv_2 _29110_ (.A(_02013_),
    .Y(_02015_));
 sky130_fd_sc_hd__inv_2 _29111_ (.A(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__inv_2 _29112_ (.A(_02028_),
    .Y(_02030_));
 sky130_fd_sc_hd__inv_2 _29113_ (.A(_02047_),
    .Y(_02049_));
 sky130_fd_sc_hd__inv_2 _29114_ (.A(_02061_),
    .Y(_02063_));
 sky130_fd_sc_hd__inv_2 _29115_ (.A(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__inv_2 _29116_ (.A(_02093_),
    .Y(_02095_));
 sky130_fd_sc_hd__inv_2 _29117_ (.A(_02106_),
    .Y(_02108_));
 sky130_fd_sc_hd__inv_2 _29118_ (.A(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__inv_2 _29119_ (.A(_02143_),
    .Y(_02145_));
 sky130_fd_sc_hd__inv_2 _29120_ (.A(_02162_),
    .Y(_02163_));
 sky130_fd_sc_hd__inv_2 _29121_ (.A(_02173_),
    .Y(_02174_));
 sky130_fd_sc_hd__inv_2 _29122_ (.A(_02192_),
    .Y(_02193_));
 sky130_fd_sc_hd__inv_2 _29123_ (.A(_02219_),
    .Y(_02220_));
 sky130_fd_sc_hd__inv_2 _29124_ (.A(_02225_),
    .Y(_02226_));
 sky130_fd_sc_hd__inv_2 _29125_ (.A(_02232_),
    .Y(_02238_));
 sky130_fd_sc_hd__inv_2 _29126_ (.A(_02253_),
    .Y(_02254_));
 sky130_fd_sc_hd__inv_2 _29127_ (.A(_02259_),
    .Y(_02261_));
 sky130_fd_sc_hd__inv_2 _29128_ (.A(_02267_),
    .Y(_02272_));
 sky130_fd_sc_hd__inv_2 _29129_ (.A(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__inv_2 _29130_ (.A(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__inv_2 _29131_ (.A(_02298_),
    .Y(_02300_));
 sky130_fd_sc_hd__inv_2 _29132_ (.A(_02306_),
    .Y(_02308_));
 sky130_fd_sc_hd__inv_2 _29133_ (.A(_02329_),
    .Y(_02331_));
 sky130_fd_sc_hd__inv_2 _29134_ (.A(_02350_),
    .Y(_02357_));
 sky130_fd_sc_hd__inv_2 _29135_ (.A(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__inv_2 _29136_ (.A(_02362_),
    .Y(_02364_));
 sky130_fd_sc_hd__inv_2 _29137_ (.A(_02380_),
    .Y(_02388_));
 sky130_fd_sc_hd__inv_2 _29138_ (.A(_02385_),
    .Y(_02386_));
 sky130_fd_sc_hd__inv_2 _29139_ (.A(_02393_),
    .Y(_02395_));
 sky130_fd_sc_hd__inv_2 _29140_ (.A(_02398_),
    .Y(_02399_));
 sky130_fd_sc_hd__inv_2 _29141_ (.A(_02410_),
    .Y(_02418_));
 sky130_fd_sc_hd__inv_2 _29142_ (.A(_02415_),
    .Y(_02416_));
 sky130_fd_sc_hd__inv_2 _29143_ (.A(_02435_),
    .Y(_02443_));
 sky130_fd_sc_hd__inv_2 _29144_ (.A(_02440_),
    .Y(_02441_));
 sky130_fd_sc_hd__inv_2 _29145_ (.A(_02447_),
    .Y(_02448_));
 sky130_fd_sc_hd__inv_2 _29146_ (.A(_02460_),
    .Y(_02468_));
 sky130_fd_sc_hd__inv_2 _29147_ (.A(_02465_),
    .Y(_02466_));
 sky130_fd_sc_hd__inv_2 _29148_ (.A(_02501_),
    .Y(_02504_));
 sky130_fd_sc_hd__inv_2 _29149_ (.A(_02524_),
    .Y(_02529_));
 sky130_fd_sc_hd__inv_2 _29150_ (.A(_00178_),
    .Y(_00222_));
 sky130_fd_sc_hd__inv_2 _29151_ (.A(_00208_),
    .Y(_03381_));
 sky130_fd_sc_hd__inv_2 _29152_ (.A(_00213_),
    .Y(_00239_));
 sky130_fd_sc_hd__inv_2 _29153_ (.A(_00218_),
    .Y(_00241_));
 sky130_fd_sc_hd__inv_2 _29154_ (.A(_00231_),
    .Y(_00258_));
 sky130_fd_sc_hd__inv_2 _29155_ (.A(_00236_),
    .Y(_00260_));
 sky130_fd_sc_hd__inv_2 _29156_ (.A(_00250_),
    .Y(_00282_));
 sky130_fd_sc_hd__inv_2 _29157_ (.A(_00255_),
    .Y(_00284_));
 sky130_fd_sc_hd__inv_2 _29158_ (.A(_00274_),
    .Y(_00313_));
 sky130_fd_sc_hd__inv_2 _29159_ (.A(_00279_),
    .Y(_00315_));
 sky130_fd_sc_hd__inv_2 _29160_ (.A(_00301_),
    .Y(_00326_));
 sky130_fd_sc_hd__inv_2 _29161_ (.A(_00305_),
    .Y(_00340_));
 sky130_fd_sc_hd__inv_2 _29162_ (.A(_00310_),
    .Y(_00342_));
 sky130_fd_sc_hd__inv_2 _29163_ (.A(_00332_),
    .Y(_00372_));
 sky130_fd_sc_hd__inv_2 _29164_ (.A(_00337_),
    .Y(_00374_));
 sky130_fd_sc_hd__inv_2 _29165_ (.A(_00353_),
    .Y(_00394_));
 sky130_fd_sc_hd__inv_2 _29166_ (.A(_00360_),
    .Y(_00416_));
 sky130_fd_sc_hd__inv_2 _29167_ (.A(_00364_),
    .Y(_00412_));
 sky130_fd_sc_hd__inv_2 _29168_ (.A(_00369_),
    .Y(_00414_));
 sky130_fd_sc_hd__inv_2 _29169_ (.A(_00381_),
    .Y(_00426_));
 sky130_fd_sc_hd__inv_2 _29170_ (.A(_00392_),
    .Y(_00431_));
 sky130_fd_sc_hd__inv_2 _29171_ (.A(_00399_),
    .Y(_00447_));
 sky130_fd_sc_hd__inv_2 _29172_ (.A(_00404_),
    .Y(_00443_));
 sky130_fd_sc_hd__inv_2 _29173_ (.A(_00409_),
    .Y(_00445_));
 sky130_fd_sc_hd__inv_2 _29174_ (.A(_00435_),
    .Y(_00475_));
 sky130_fd_sc_hd__inv_2 _29175_ (.A(_00440_),
    .Y(_00476_));
 sky130_fd_sc_hd__inv_2 _29176_ (.A(_00472_),
    .Y(_00511_));
 sky130_fd_sc_hd__inv_2 _29177_ (.A(_00499_),
    .Y(_00542_));
 sky130_fd_sc_hd__inv_2 _29178_ (.A(_00508_),
    .Y(_00553_));
 sky130_fd_sc_hd__inv_2 _29179_ (.A(_00514_),
    .Y(_03471_));
 sky130_fd_sc_hd__inv_2 _29180_ (.A(_00516_),
    .Y(_00562_));
 sky130_fd_sc_hd__inv_2 _29181_ (.A(_00532_),
    .Y(_00586_));
 sky130_fd_sc_hd__inv_2 _29182_ (.A(_00540_),
    .Y(_00584_));
 sky130_fd_sc_hd__inv_2 _29183_ (.A(_00550_),
    .Y(_00596_));
 sky130_fd_sc_hd__inv_2 _29184_ (.A(_00556_),
    .Y(_03482_));
 sky130_fd_sc_hd__inv_2 _29185_ (.A(_00582_),
    .Y(_00635_));
 sky130_fd_sc_hd__inv_2 _29186_ (.A(_00593_),
    .Y(_00646_));
 sky130_fd_sc_hd__inv_2 _29187_ (.A(_00599_),
    .Y(_03491_));
 sky130_fd_sc_hd__inv_2 _29188_ (.A(_00602_),
    .Y(_00655_));
 sky130_fd_sc_hd__inv_2 _29189_ (.A(_00621_),
    .Y(_00675_));
 sky130_fd_sc_hd__inv_2 _29190_ (.A(_00633_),
    .Y(_00683_));
 sky130_fd_sc_hd__inv_2 _29191_ (.A(_00643_),
    .Y(_00694_));
 sky130_fd_sc_hd__inv_2 _29192_ (.A(_00649_),
    .Y(_03503_));
 sky130_fd_sc_hd__inv_2 _29193_ (.A(_00652_),
    .Y(_00703_));
 sky130_fd_sc_hd__inv_2 _29194_ (.A(_00681_),
    .Y(_00733_));
 sky130_fd_sc_hd__inv_2 _29195_ (.A(_00691_),
    .Y(_00744_));
 sky130_fd_sc_hd__inv_2 _29196_ (.A(_00697_),
    .Y(_03517_));
 sky130_fd_sc_hd__inv_2 _29197_ (.A(_00700_),
    .Y(_00752_));
 sky130_fd_sc_hd__inv_2 _29198_ (.A(_00727_),
    .Y(_00778_));
 sky130_fd_sc_hd__inv_2 _29199_ (.A(_00731_),
    .Y(_00787_));
 sky130_fd_sc_hd__inv_2 _29200_ (.A(_00741_),
    .Y(_00798_));
 sky130_fd_sc_hd__inv_2 _29201_ (.A(_00748_),
    .Y(_03528_));
 sky130_fd_sc_hd__inv_2 _29202_ (.A(_00760_),
    .Y(_00818_));
 sky130_fd_sc_hd__inv_2 _29203_ (.A(_00785_),
    .Y(_00841_));
 sky130_fd_sc_hd__inv_2 _29204_ (.A(_00795_),
    .Y(_00852_));
 sky130_fd_sc_hd__inv_2 _29205_ (.A(_00804_),
    .Y(_00864_));
 sky130_fd_sc_hd__inv_2 _29206_ (.A(_00827_),
    .Y(_00886_));
 sky130_fd_sc_hd__inv_2 _29207_ (.A(_00839_),
    .Y(_00898_));
 sky130_fd_sc_hd__inv_2 _29208_ (.A(_00849_),
    .Y(_00909_));
 sky130_fd_sc_hd__inv_2 _29209_ (.A(_00891_),
    .Y(_00973_));
 sky130_fd_sc_hd__inv_2 _29210_ (.A(_00896_),
    .Y(_00953_));
 sky130_fd_sc_hd__inv_2 _29211_ (.A(_00906_),
    .Y(_00964_));
 sky130_fd_sc_hd__inv_2 _29212_ (.A(_00951_),
    .Y(_01013_));
 sky130_fd_sc_hd__inv_2 _29213_ (.A(_00961_),
    .Y(_01024_));
 sky130_fd_sc_hd__inv_2 _29214_ (.A(_00995_),
    .Y(_01058_));
 sky130_fd_sc_hd__inv_2 _29215_ (.A(_01011_),
    .Y(_01072_));
 sky130_fd_sc_hd__inv_2 _29216_ (.A(_01021_),
    .Y(_01085_));
 sky130_fd_sc_hd__inv_2 _29217_ (.A(_01051_),
    .Y(_01131_));
 sky130_fd_sc_hd__inv_2 _29218_ (.A(_01056_),
    .Y(_01122_));
 sky130_fd_sc_hd__inv_2 _29219_ (.A(_01076_),
    .Y(_01149_));
 sky130_fd_sc_hd__inv_2 _29220_ (.A(_01081_),
    .Y(_01151_));
 sky130_fd_sc_hd__inv_2 _29221_ (.A(_01120_),
    .Y(_01186_));
 sky130_fd_sc_hd__inv_2 _29222_ (.A(_01135_),
    .Y(_01199_));
 sky130_fd_sc_hd__inv_2 _29223_ (.A(_01141_),
    .Y(_01212_));
 sky130_fd_sc_hd__inv_2 _29224_ (.A(_01146_),
    .Y(_01214_));
 sky130_fd_sc_hd__inv_2 _29225_ (.A(_01181_),
    .Y(_01256_));
 sky130_fd_sc_hd__inv_2 _29226_ (.A(_01197_),
    .Y(_01262_));
 sky130_fd_sc_hd__inv_2 _29227_ (.A(_01204_),
    .Y(_01275_));
 sky130_fd_sc_hd__inv_2 _29228_ (.A(_01209_),
    .Y(_01277_));
 sky130_fd_sc_hd__inv_2 _29229_ (.A(_01246_),
    .Y(_01304_));
 sky130_fd_sc_hd__inv_2 _29230_ (.A(_01260_),
    .Y(_01317_));
 sky130_fd_sc_hd__inv_2 _29231_ (.A(_01267_),
    .Y(_01330_));
 sky130_fd_sc_hd__inv_2 _29232_ (.A(_01272_),
    .Y(_01332_));
 sky130_fd_sc_hd__inv_2 _29233_ (.A(_01315_),
    .Y(_01385_));
 sky130_fd_sc_hd__inv_2 _29234_ (.A(_01322_),
    .Y(_01395_));
 sky130_fd_sc_hd__inv_2 _29235_ (.A(_01327_),
    .Y(_01397_));
 sky130_fd_sc_hd__inv_2 _29236_ (.A(_01344_),
    .Y(_01407_));
 sky130_fd_sc_hd__inv_2 _29237_ (.A(_01370_),
    .Y(_01429_));
 sky130_fd_sc_hd__inv_2 _29238_ (.A(_01383_),
    .Y(_01442_));
 sky130_fd_sc_hd__inv_2 _29239_ (.A(_01390_),
    .Y(_01454_));
 sky130_fd_sc_hd__inv_2 _29240_ (.A(_01440_),
    .Y(_01502_));
 sky130_fd_sc_hd__inv_2 _29241_ (.A(_01447_),
    .Y(_01509_));
 sky130_fd_sc_hd__inv_2 _29242_ (.A(_01487_),
    .Y(_01548_));
 sky130_fd_sc_hd__inv_2 _29243_ (.A(_01500_),
    .Y(_01562_));
 sky130_fd_sc_hd__inv_2 _29244_ (.A(_01507_),
    .Y(_01568_));
 sky130_fd_sc_hd__inv_2 _29245_ (.A(_01540_),
    .Y(_01605_));
 sky130_fd_sc_hd__inv_2 _29246_ (.A(_01546_),
    .Y(_01603_));
 sky130_fd_sc_hd__inv_2 _29247_ (.A(_01560_),
    .Y(_01618_));
 sky130_fd_sc_hd__inv_2 _29248_ (.A(_01566_),
    .Y(_01623_));
 sky130_fd_sc_hd__inv_2 _29249_ (.A(_01601_),
    .Y(_01657_));
 sky130_fd_sc_hd__inv_2 _29250_ (.A(_01616_),
    .Y(_01671_));
 sky130_fd_sc_hd__inv_2 _29251_ (.A(_01655_),
    .Y(_01709_));
 sky130_fd_sc_hd__inv_2 _29252_ (.A(_01669_),
    .Y(_01721_));
 sky130_fd_sc_hd__inv_2 _29253_ (.A(_01707_),
    .Y(_01759_));
 sky130_fd_sc_hd__inv_2 _29254_ (.A(_01757_),
    .Y(_01808_));
 sky130_fd_sc_hd__inv_2 _29255_ (.A(_01779_),
    .Y(_01828_));
 sky130_fd_sc_hd__inv_2 _29256_ (.A(_01806_),
    .Y(_01862_));
 sky130_fd_sc_hd__inv_2 _29257_ (.A(_01816_),
    .Y(_01873_));
 sky130_fd_sc_hd__inv_2 _29258_ (.A(_01826_),
    .Y(_01881_));
 sky130_fd_sc_hd__inv_2 _29259_ (.A(_01845_),
    .Y(_01900_));
 sky130_fd_sc_hd__inv_2 _29260_ (.A(_01851_),
    .Y(_01910_));
 sky130_fd_sc_hd__inv_2 _29261_ (.A(_01860_),
    .Y(_01915_));
 sky130_fd_sc_hd__inv_2 _29262_ (.A(_01869_),
    .Y(_01926_));
 sky130_fd_sc_hd__inv_2 _29263_ (.A(_01879_),
    .Y(_01934_));
 sky130_fd_sc_hd__inv_2 _29264_ (.A(_01898_),
    .Y(_01953_));
 sky130_fd_sc_hd__inv_2 _29265_ (.A(_01905_),
    .Y(_01962_));
 sky130_fd_sc_hd__inv_2 _29266_ (.A(_01919_),
    .Y(_01973_));
 sky130_fd_sc_hd__inv_2 _29267_ (.A(_01932_),
    .Y(_01982_));
 sky130_fd_sc_hd__inv_2 _29268_ (.A(_01951_),
    .Y(_02001_));
 sky130_fd_sc_hd__inv_2 _29269_ (.A(_01966_),
    .Y(_02014_));
 sky130_fd_sc_hd__inv_2 _29270_ (.A(_01976_),
    .Y(_02072_));
 sky130_fd_sc_hd__inv_2 _29271_ (.A(_01980_),
    .Y(_02029_));
 sky130_fd_sc_hd__inv_2 _29272_ (.A(_01999_),
    .Y(_02048_));
 sky130_fd_sc_hd__inv_2 _29273_ (.A(_02012_),
    .Y(_02062_));
 sky130_fd_sc_hd__inv_2 _29274_ (.A(_02022_),
    .Y(_02071_));
 sky130_fd_sc_hd__inv_2 _29275_ (.A(_02026_),
    .Y(_02075_));
 sky130_fd_sc_hd__inv_2 _29276_ (.A(_02027_),
    .Y(_02076_));
 sky130_fd_sc_hd__inv_2 _29277_ (.A(_02046_),
    .Y(_02094_));
 sky130_fd_sc_hd__inv_2 _29278_ (.A(_02060_),
    .Y(_02107_));
 sky130_fd_sc_hd__inv_2 _29279_ (.A(_02092_),
    .Y(_02131_));
 sky130_fd_sc_hd__inv_2 _29280_ (.A(_02105_),
    .Y(_02141_));
 sky130_fd_sc_hd__inv_2 _29281_ (.A(_02113_),
    .Y(_02144_));
 sky130_fd_sc_hd__inv_2 _29282_ (.A(_02142_),
    .Y(_02177_));
 sky130_fd_sc_hd__inv_2 _29283_ (.A(_02161_),
    .Y(_02197_));
 sky130_fd_sc_hd__inv_2 _29284_ (.A(_02172_),
    .Y(_02204_));
 sky130_fd_sc_hd__inv_2 _29285_ (.A(_02191_),
    .Y(_02227_));
 sky130_fd_sc_hd__inv_2 _29286_ (.A(_02218_),
    .Y(_02262_));
 sky130_fd_sc_hd__inv_2 _29287_ (.A(_02224_),
    .Y(_02260_));
 sky130_fd_sc_hd__inv_2 _29288_ (.A(_02231_),
    .Y(_02271_));
 sky130_fd_sc_hd__inv_2 _29289_ (.A(_02252_),
    .Y(_02301_));
 sky130_fd_sc_hd__inv_2 _29290_ (.A(_02258_),
    .Y(_02299_));
 sky130_fd_sc_hd__inv_2 _29291_ (.A(_02266_),
    .Y(_02307_));
 sky130_fd_sc_hd__inv_2 _29292_ (.A(_02274_),
    .Y(_02310_));
 sky130_fd_sc_hd__inv_2 _29293_ (.A(_02276_),
    .Y(_02312_));
 sky130_fd_sc_hd__inv_2 _29294_ (.A(_02291_),
    .Y(_02332_));
 sky130_fd_sc_hd__inv_2 _29295_ (.A(_02297_),
    .Y(_02330_));
 sky130_fd_sc_hd__inv_2 _29296_ (.A(_02305_),
    .Y(_02336_));
 sky130_fd_sc_hd__inv_2 _29297_ (.A(_02328_),
    .Y(_02363_));
 sky130_fd_sc_hd__inv_2 _29298_ (.A(_02337_),
    .Y(_02369_));
 sky130_fd_sc_hd__inv_2 _29299_ (.A(_02349_),
    .Y(_02387_));
 sky130_fd_sc_hd__inv_2 _29300_ (.A(_02354_),
    .Y(_02396_));
 sky130_fd_sc_hd__inv_2 _29301_ (.A(_02361_),
    .Y(_02394_));
 sky130_fd_sc_hd__inv_2 _29302_ (.A(_02379_),
    .Y(_02417_));
 sky130_fd_sc_hd__inv_2 _29303_ (.A(_02384_),
    .Y(_02423_));
 sky130_fd_sc_hd__inv_2 _29304_ (.A(_02392_),
    .Y(_02422_));
 sky130_fd_sc_hd__inv_2 _29305_ (.A(_02409_),
    .Y(_02442_));
 sky130_fd_sc_hd__inv_2 _29306_ (.A(_02414_),
    .Y(_02449_));
 sky130_fd_sc_hd__inv_2 _29307_ (.A(_02434_),
    .Y(_02467_));
 sky130_fd_sc_hd__inv_2 _29308_ (.A(_02439_),
    .Y(_02470_));
 sky130_fd_sc_hd__inv_2 _29309_ (.A(_02446_),
    .Y(_02469_));
 sky130_fd_sc_hd__inv_2 _29310_ (.A(_02459_),
    .Y(_02484_));
 sky130_fd_sc_hd__inv_2 _29311_ (.A(_02464_),
    .Y(_02485_));
 sky130_fd_sc_hd__inv_2 _29312_ (.A(_02495_),
    .Y(_02515_));
 sky130_fd_sc_hd__inv_2 _29313_ (.A(_02498_),
    .Y(_02518_));
 sky130_fd_sc_hd__inv_2 _29314_ (.A(_01673_),
    .Y(_01724_));
 sky130_fd_sc_hd__inv_2 _29315_ (.A(_01728_),
    .Y(_01730_));
 sky130_fd_sc_hd__inv_2 _29316_ (.A(_01677_),
    .Y(_01729_));
 sky130_fd_sc_hd__inv_2 _29317_ (.A(_01675_),
    .Y(_02549_));
 sky130_fd_sc_hd__inv_2 _29318_ (.A(_01686_),
    .Y(_02551_));
 sky130_fd_sc_hd__inv_2 _29319_ (.A(_01774_),
    .Y(_01776_));
 sky130_fd_sc_hd__inv_2 _29320_ (.A(_01722_),
    .Y(_01775_));
 sky130_fd_sc_hd__inv_2 _29321_ (.A(_01723_),
    .Y(_01778_));
 sky130_fd_sc_hd__inv_2 _29322_ (.A(_01736_),
    .Y(_02557_));
 sky130_fd_sc_hd__inv_2 _29323_ (.A(_01822_),
    .Y(_01824_));
 sky130_fd_sc_hd__inv_2 _29324_ (.A(_01773_),
    .Y(_01823_));
 sky130_fd_sc_hd__inv_2 _29325_ (.A(_01782_),
    .Y(_02561_));
 sky130_fd_sc_hd__inv_2 _29326_ (.A(_01785_),
    .Y(_02563_));
 sky130_fd_sc_hd__nor2_1 _29327_ (.A(net1129),
    .B(net1211),
    .Y(_01848_));
 sky130_fd_sc_hd__inv_2 _29328_ (.A(_01875_),
    .Y(_01877_));
 sky130_fd_sc_hd__inv_2 _29329_ (.A(_01821_),
    .Y(_01876_));
 sky130_fd_sc_hd__inv_2 _29330_ (.A(_01830_),
    .Y(_02567_));
 sky130_fd_sc_hd__inv_2 _29331_ (.A(_01833_),
    .Y(_02569_));
 sky130_fd_sc_hd__nor2_1 _29332_ (.A(net1323),
    .B(net1108),
    .Y(_01921_));
 sky130_fd_sc_hd__inv_2 _29333_ (.A(_01928_),
    .Y(_01930_));
 sky130_fd_sc_hd__inv_2 _29334_ (.A(_01874_),
    .Y(_01929_));
 sky130_fd_sc_hd__inv_2 _29335_ (.A(_01883_),
    .Y(_02573_));
 sky130_fd_sc_hd__inv_2 _29336_ (.A(_01886_),
    .Y(_02575_));
 sky130_fd_sc_hd__inv_2 _29337_ (.A(_01927_),
    .Y(_01978_));
 sky130_fd_sc_hd__inv_2 _29338_ (.A(_01936_),
    .Y(_02579_));
 sky130_fd_sc_hd__inv_2 _29339_ (.A(_01939_),
    .Y(_02581_));
 sky130_fd_sc_hd__inv_2 _29340_ (.A(_01975_),
    .Y(_02025_));
 sky130_fd_sc_hd__inv_2 _29341_ (.A(_01984_),
    .Y(_02585_));
 sky130_fd_sc_hd__inv_2 _29342_ (.A(_01987_),
    .Y(_02587_));
 sky130_fd_sc_hd__inv_2 _29343_ (.A(_02019_),
    .Y(_02067_));
 sky130_fd_sc_hd__inv_2 _29344_ (.A(_02031_),
    .Y(_02591_));
 sky130_fd_sc_hd__inv_2 _29345_ (.A(_02034_),
    .Y(_02593_));
 sky130_fd_sc_hd__inv_2 _29346_ (.A(_02065_),
    .Y(_02109_));
 sky130_fd_sc_hd__inv_2 _29347_ (.A(_02074_),
    .Y(_02112_));
 sky130_fd_sc_hd__inv_2 _29348_ (.A(_02077_),
    .Y(_02597_));
 sky130_fd_sc_hd__inv_2 _29349_ (.A(_02080_),
    .Y(_02599_));
 sky130_fd_sc_hd__inv_2 _29350_ (.A(_02116_),
    .Y(_02604_));
 sky130_fd_sc_hd__inv_2 _29351_ (.A(_02119_),
    .Y(_02606_));
 sky130_fd_sc_hd__inv_2 _29352_ (.A(_02146_),
    .Y(_02610_));
 sky130_fd_sc_hd__inv_2 _29353_ (.A(_02149_),
    .Y(_02612_));
 sky130_fd_sc_hd__inv_2 _29354_ (.A(_02179_),
    .Y(_02617_));
 sky130_fd_sc_hd__inv_2 _29355_ (.A(_02182_),
    .Y(_02619_));
 sky130_fd_sc_hd__inv_2 _29356_ (.A(_02206_),
    .Y(_02623_));
 sky130_fd_sc_hd__inv_2 _29357_ (.A(_02209_),
    .Y(_02625_));
 sky130_fd_sc_hd__inv_2 _29358_ (.A(_02235_),
    .Y(_02273_));
 sky130_fd_sc_hd__inv_2 _29359_ (.A(_02239_),
    .Y(_02275_));
 sky130_fd_sc_hd__inv_2 _29360_ (.A(_02240_),
    .Y(_02629_));
 sky130_fd_sc_hd__inv_2 _29361_ (.A(_02243_),
    .Y(_02631_));
 sky130_fd_sc_hd__inv_2 _29362_ (.A(_02279_),
    .Y(_02635_));
 sky130_fd_sc_hd__inv_2 _29363_ (.A(_02282_),
    .Y(_02637_));
 sky130_fd_sc_hd__inv_2 _29364_ (.A(_02313_),
    .Y(_02642_));
 sky130_fd_sc_hd__inv_2 _29365_ (.A(_02316_),
    .Y(_02644_));
 sky130_fd_sc_hd__inv_2 _29366_ (.A(_02340_),
    .Y(_02648_));
 sky130_fd_sc_hd__inv_2 _29367_ (.A(_02343_),
    .Y(_02650_));
 sky130_fd_sc_hd__inv_2 _29368_ (.A(_02370_),
    .Y(_02654_));
 sky130_fd_sc_hd__inv_2 _29369_ (.A(_02373_),
    .Y(_02656_));
 sky130_fd_sc_hd__inv_2 _29370_ (.A(_02400_),
    .Y(_02660_));
 sky130_fd_sc_hd__inv_2 _29371_ (.A(_02403_),
    .Y(_02662_));
 sky130_fd_sc_hd__inv_2 _29372_ (.A(_02425_),
    .Y(_02666_));
 sky130_fd_sc_hd__inv_2 _29373_ (.A(_02428_),
    .Y(_02668_));
 sky130_fd_sc_hd__inv_2 _29374_ (.A(_02450_),
    .Y(_02672_));
 sky130_fd_sc_hd__inv_2 _29375_ (.A(_02453_),
    .Y(_02674_));
 sky130_fd_sc_hd__inv_2 _29376_ (.A(_02471_),
    .Y(_02679_));
 sky130_fd_sc_hd__inv_2 _29377_ (.A(_02474_),
    .Y(_02681_));
 sky130_fd_sc_hd__inv_2 _29378_ (.A(_02480_),
    .Y(_02500_));
 sky130_fd_sc_hd__inv_2 _29379_ (.A(_02486_),
    .Y(_02685_));
 sky130_fd_sc_hd__inv_2 _29380_ (.A(_02489_),
    .Y(_02687_));
 sky130_fd_sc_hd__inv_2 _29381_ (.A(_02503_),
    .Y(_02525_));
 sky130_fd_sc_hd__inv_2 _29382_ (.A(_02505_),
    .Y(_02692_));
 sky130_fd_sc_hd__inv_2 _29383_ (.A(_02508_),
    .Y(_02695_));
 sky130_fd_sc_hd__inv_2 _29384_ (.A(\inst$top.soc.uart_0._phy.tx.lower.bitno[0] ),
    .Y(_02702_));
 sky130_fd_sc_hd__inv_2 _29385_ (.A(\inst$top.soc.uart_0._phy.rx.lower.bitno[0] ),
    .Y(_02714_));
 sky130_fd_sc_hd__inv_1 _29386_ (.A(net1668),
    .Y(_09353_));
 sky130_fd_sc_hd__a21oi_1 _29387_ (.A1(_09353_),
    .A2(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[1] ),
    .B1(\inst$top.soc.uart_0._phy.rx.lower.timer[1] ),
    .Y(_02719_));
 sky130_fd_sc_hd__inv_2 _29388_ (.A(\inst$top.soc.spiflash.ctrl.i_data_count[0] ),
    .Y(_02732_));
 sky130_fd_sc_hd__inv_2 _29389_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[0] ),
    .Y(_02739_));
 sky130_fd_sc_hd__inv_2 _29390_ (.A(\inst$top.soc.cpu.divider.timer[0] ),
    .Y(_02857_));
 sky130_fd_sc_hd__inv_2 _29391_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__2._storage[0] ),
    .Y(_02868_));
 sky130_fd_sc_hd__inv_2 _29392_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__0._storage[0] ),
    .Y(_02871_));
 sky130_fd_sc_hd__inv_2 _29393_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__3._storage[0] ),
    .Y(_02874_));
 sky130_fd_sc_hd__inv_2 _29394_ (.A(\inst$top.soc.uart_0._phy.rx.lower.fsm_state[0] ),
    .Y(_02877_));
 sky130_fd_sc_hd__inv_2 _29395_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__1._storage[0] ),
    .Y(_02884_));
 sky130_fd_sc_hd__inv_2 _29396_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__0._storage[0] ),
    .Y(_02887_));
 sky130_fd_sc_hd__inv_2 _29397_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__2._storage[0] ),
    .Y(_02890_));
 sky130_fd_sc_hd__inv_2 _29398_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__1._storage[0] ),
    .Y(_02893_));
 sky130_fd_sc_hd__inv_2 _29399_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__3._storage[0] ),
    .Y(_02896_));
 sky130_fd_sc_hd__inv_2 _29400_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__7._storage[0] ),
    .Y(_02899_));
 sky130_fd_sc_hd__inv_2 _29401_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__6._storage[0] ),
    .Y(_02902_));
 sky130_fd_sc_hd__inv_2 _29402_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__5._storage[0] ),
    .Y(_02905_));
 sky130_fd_sc_hd__inv_2 _29403_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__4._storage[0] ),
    .Y(_02908_));
 sky130_fd_sc_hd__inv_2 _29404_ (.A(_00209_),
    .Y(_02914_));
 sky130_fd_sc_hd__inv_2 _29405_ (.A(_03095_),
    .Y(_03091_));
 sky130_fd_sc_hd__inv_2 _29406_ (.A(_03307_),
    .Y(_03303_));
 sky130_fd_sc_hd__inv_2 _29407_ (.A(_00188_),
    .Y(_03366_));
 sky130_fd_sc_hd__inv_2 _29408_ (.A(_00199_),
    .Y(_03371_));
 sky130_fd_sc_hd__inv_2 _29409_ (.A(_00200_),
    .Y(_03375_));
 sky130_fd_sc_hd__inv_2 _29410_ (.A(_00204_),
    .Y(_03380_));
 sky130_fd_sc_hd__inv_2 _29411_ (.A(_00224_),
    .Y(_03384_));
 sky130_fd_sc_hd__inv_2 _29412_ (.A(_00187_),
    .Y(_03385_));
 sky130_fd_sc_hd__inv_2 _29413_ (.A(_00243_),
    .Y(_03388_));
 sky130_fd_sc_hd__inv_2 _29414_ (.A(_00223_),
    .Y(_03389_));
 sky130_fd_sc_hd__inv_2 _29415_ (.A(_00262_),
    .Y(_03394_));
 sky130_fd_sc_hd__inv_2 _29416_ (.A(_00242_),
    .Y(_03396_));
 sky130_fd_sc_hd__inv_2 _29417_ (.A(_00286_),
    .Y(_00287_));
 sky130_fd_sc_hd__inv_2 _29418_ (.A(_00261_),
    .Y(_03405_));
 sky130_fd_sc_hd__inv_2 _29419_ (.A(_00266_),
    .Y(_03406_));
 sky130_fd_sc_hd__inv_2 _29420_ (.A(_00317_),
    .Y(_00318_));
 sky130_fd_sc_hd__inv_2 _29421_ (.A(_00285_),
    .Y(_03411_));
 sky130_fd_sc_hd__inv_2 _29422_ (.A(_00292_),
    .Y(_03412_));
 sky130_fd_sc_hd__inv_2 _29423_ (.A(_00322_),
    .Y(_03415_));
 sky130_fd_sc_hd__inv_2 _29424_ (.A(_00344_),
    .Y(_00345_));
 sky130_fd_sc_hd__inv_2 _29425_ (.A(_00316_),
    .Y(_03418_));
 sky130_fd_sc_hd__inv_2 _29426_ (.A(_00349_),
    .Y(_03424_));
 sky130_fd_sc_hd__inv_2 _29427_ (.A(_00357_),
    .Y(_00359_));
 sky130_fd_sc_hd__inv_2 _29428_ (.A(_00327_),
    .Y(_00358_));
 sky130_fd_sc_hd__inv_2 _29429_ (.A(_00376_),
    .Y(_00377_));
 sky130_fd_sc_hd__inv_2 _29430_ (.A(_00343_),
    .Y(_03425_));
 sky130_fd_sc_hd__nor2_1 _29431_ (.A(net1707),
    .B(_03017_),
    .Y(_00379_));
 sky130_fd_sc_hd__nor2_1 _29432_ (.A(net1318),
    .B(net1367),
    .Y(_00378_));
 sky130_fd_sc_hd__inv_2 _29433_ (.A(_00396_),
    .Y(_00398_));
 sky130_fd_sc_hd__inv_2 _29434_ (.A(_00356_),
    .Y(_00397_));
 sky130_fd_sc_hd__inv_2 _29435_ (.A(_00375_),
    .Y(_03431_));
 sky130_fd_sc_hd__inv_2 _29436_ (.A(_00427_),
    .Y(_03434_));
 sky130_fd_sc_hd__inv_2 _29437_ (.A(_00418_),
    .Y(_03436_));
 sky130_fd_sc_hd__inv_2 _29438_ (.A(_00415_),
    .Y(_03440_));
 sky130_fd_sc_hd__inv_2 _29439_ (.A(_00461_),
    .Y(_03446_));
 sky130_fd_sc_hd__inv_2 _29440_ (.A(_00448_),
    .Y(_03448_));
 sky130_fd_sc_hd__inv_2 _29441_ (.A(_00446_),
    .Y(_03451_));
 sky130_fd_sc_hd__inv_2 _29442_ (.A(_00495_),
    .Y(_03456_));
 sky130_fd_sc_hd__inv_2 _29443_ (.A(_00515_),
    .Y(_03458_));
 sky130_fd_sc_hd__inv_2 _29444_ (.A(_00477_),
    .Y(_03460_));
 sky130_fd_sc_hd__inv_2 _29445_ (.A(_00483_),
    .Y(_03461_));
 sky130_fd_sc_hd__nor2_1 _29446_ (.A(net1407),
    .B(net1157),
    .Y(_00529_));
 sky130_fd_sc_hd__inv_2 _29447_ (.A(_00535_),
    .Y(_00536_));
 sky130_fd_sc_hd__inv_2 _29448_ (.A(_00557_),
    .Y(_03467_));
 sky130_fd_sc_hd__inv_2 _29449_ (.A(_00512_),
    .Y(_03470_));
 sky130_fd_sc_hd__inv_2 _29450_ (.A(_00520_),
    .Y(_03473_));
 sky130_fd_sc_hd__inv_2 _29451_ (.A(_00577_),
    .Y(_00578_));
 sky130_fd_sc_hd__inv_2 _29452_ (.A(_00600_),
    .Y(_00601_));
 sky130_fd_sc_hd__inv_2 _29453_ (.A(_00554_),
    .Y(_03481_));
 sky130_fd_sc_hd__inv_2 _29454_ (.A(_00563_),
    .Y(_03484_));
 sky130_fd_sc_hd__inv_2 _29455_ (.A(_00618_),
    .Y(_00620_));
 sky130_fd_sc_hd__inv_2 _29456_ (.A(_00569_),
    .Y(_00619_));
 sky130_fd_sc_hd__inv_2 _29457_ (.A(_00628_),
    .Y(_00629_));
 sky130_fd_sc_hd__inv_2 _29458_ (.A(_00650_),
    .Y(_00651_));
 sky130_fd_sc_hd__inv_2 _29459_ (.A(_00597_),
    .Y(_03490_));
 sky130_fd_sc_hd__inv_2 _29460_ (.A(_00608_),
    .Y(_03493_));
 sky130_fd_sc_hd__inv_2 _29461_ (.A(_00664_),
    .Y(_03497_));
 sky130_fd_sc_hd__inv_2 _29462_ (.A(_00698_),
    .Y(_00699_));
 sky130_fd_sc_hd__inv_2 _29463_ (.A(_00647_),
    .Y(_03502_));
 sky130_fd_sc_hd__inv_2 _29464_ (.A(_00658_),
    .Y(_03505_));
 sky130_fd_sc_hd__inv_2 _29465_ (.A(_00712_),
    .Y(_03512_));
 sky130_fd_sc_hd__inv_2 _29466_ (.A(_00668_),
    .Y(_00725_));
 sky130_fd_sc_hd__inv_2 _29467_ (.A(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hd__inv_2 _29468_ (.A(_00676_),
    .Y(_03514_));
 sky130_fd_sc_hd__inv_2 _29469_ (.A(_00695_),
    .Y(_03516_));
 sky130_fd_sc_hd__inv_2 _29470_ (.A(_00706_),
    .Y(_03519_));
 sky130_fd_sc_hd__nor2_1 _29471_ (.A(net1708),
    .B(net1211),
    .Y(_00758_));
 sky130_fd_sc_hd__nor2_1 _29472_ (.A(net1438),
    .B(net1368),
    .Y(_00757_));
 sky130_fd_sc_hd__inv_2 _29473_ (.A(_00781_),
    .Y(_03525_));
 sky130_fd_sc_hd__inv_2 _29474_ (.A(_00801_),
    .Y(_00803_));
 sky130_fd_sc_hd__inv_2 _29475_ (.A(_00746_),
    .Y(_00802_));
 sky130_fd_sc_hd__inv_2 _29476_ (.A(_00745_),
    .Y(_03527_));
 sky130_fd_sc_hd__inv_2 _29477_ (.A(_00754_),
    .Y(_03530_));
 sky130_fd_sc_hd__inv_2 _29478_ (.A(_00767_),
    .Y(_03534_));
 sky130_fd_sc_hd__nor2_1 _29479_ (.A(_03017_),
    .B(_05912_),
    .Y(_00824_));
 sky130_fd_sc_hd__inv_2 _29480_ (.A(_00835_),
    .Y(_03538_));
 sky130_fd_sc_hd__inv_2 _29481_ (.A(_00855_),
    .Y(_00857_));
 sky130_fd_sc_hd__inv_2 _29482_ (.A(_00800_),
    .Y(_00856_));
 sky130_fd_sc_hd__inv_2 _29483_ (.A(_00799_),
    .Y(_03541_));
 sky130_fd_sc_hd__inv_2 _29484_ (.A(_00809_),
    .Y(_03543_));
 sky130_fd_sc_hd__inv_2 _29485_ (.A(_00819_),
    .Y(_03549_));
 sky130_fd_sc_hd__inv_2 _29486_ (.A(_00889_),
    .Y(_00890_));
 sky130_fd_sc_hd__inv_2 _29487_ (.A(_00912_),
    .Y(_00914_));
 sky130_fd_sc_hd__inv_2 _29488_ (.A(_00854_),
    .Y(_00913_));
 sky130_fd_sc_hd__inv_2 _29489_ (.A(_00853_),
    .Y(_03553_));
 sky130_fd_sc_hd__inv_2 _29490_ (.A(_00866_),
    .Y(_03555_));
 sky130_fd_sc_hd__inv_2 _29491_ (.A(_00875_),
    .Y(_03560_));
 sky130_fd_sc_hd__inv_2 _29492_ (.A(_00967_),
    .Y(_00969_));
 sky130_fd_sc_hd__inv_2 _29493_ (.A(_00911_),
    .Y(_00968_));
 sky130_fd_sc_hd__inv_2 _29494_ (.A(_00910_),
    .Y(_03565_));
 sky130_fd_sc_hd__inv_2 _29495_ (.A(_00922_),
    .Y(_03567_));
 sky130_fd_sc_hd__inv_2 _29496_ (.A(_00991_),
    .Y(_03574_));
 sky130_fd_sc_hd__inv_2 _29497_ (.A(_01027_),
    .Y(_01029_));
 sky130_fd_sc_hd__inv_2 _29498_ (.A(_00966_),
    .Y(_01028_));
 sky130_fd_sc_hd__inv_2 _29499_ (.A(_00965_),
    .Y(_03577_));
 sky130_fd_sc_hd__inv_2 _29500_ (.A(_00976_),
    .Y(_03579_));
 sky130_fd_sc_hd__nor2_1 _29501_ (.A(net1708),
    .B(_05826_),
    .Y(_03583_));
 sky130_fd_sc_hd__inv_2 _29502_ (.A(_00982_),
    .Y(_03586_));
 sky130_fd_sc_hd__inv_2 _29503_ (.A(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__inv_2 _29504_ (.A(_01088_),
    .Y(_01090_));
 sky130_fd_sc_hd__inv_2 _29505_ (.A(_01026_),
    .Y(_01089_));
 sky130_fd_sc_hd__inv_2 _29506_ (.A(_01025_),
    .Y(_03590_));
 sky130_fd_sc_hd__inv_2 _29507_ (.A(_01035_),
    .Y(_03592_));
 sky130_fd_sc_hd__inv_2 _29508_ (.A(_01107_),
    .Y(_03596_));
 sky130_fd_sc_hd__inv_2 _29509_ (.A(_01154_),
    .Y(_01156_));
 sky130_fd_sc_hd__inv_2 _29510_ (.A(_01087_),
    .Y(_01155_));
 sky130_fd_sc_hd__inv_2 _29511_ (.A(_01086_),
    .Y(_03599_));
 sky130_fd_sc_hd__inv_2 _29512_ (.A(_01096_),
    .Y(_03601_));
 sky130_fd_sc_hd__inv_2 _29513_ (.A(_01168_),
    .Y(_03605_));
 sky130_fd_sc_hd__inv_2 _29514_ (.A(_01172_),
    .Y(_03608_));
 sky130_fd_sc_hd__inv_2 _29515_ (.A(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__inv_2 _29516_ (.A(_01216_),
    .Y(_01218_));
 sky130_fd_sc_hd__inv_2 _29517_ (.A(_01153_),
    .Y(_01217_));
 sky130_fd_sc_hd__inv_2 _29518_ (.A(_01152_),
    .Y(_03610_));
 sky130_fd_sc_hd__inv_2 _29519_ (.A(_01162_),
    .Y(_03612_));
 sky130_fd_sc_hd__inv_2 _29520_ (.A(_01230_),
    .Y(_03619_));
 sky130_fd_sc_hd__inv_2 _29521_ (.A(_01215_),
    .Y(_03622_));
 sky130_fd_sc_hd__inv_2 _29522_ (.A(_01224_),
    .Y(_03624_));
 sky130_fd_sc_hd__nor2_1 _29523_ (.A(net1740),
    .B(net1708),
    .Y(_03628_));
 sky130_fd_sc_hd__inv_2 _29524_ (.A(_01335_),
    .Y(_01337_));
 sky130_fd_sc_hd__inv_2 _29525_ (.A(_01279_),
    .Y(_01336_));
 sky130_fd_sc_hd__inv_2 _29526_ (.A(_01278_),
    .Y(_01342_));
 sky130_fd_sc_hd__inv_2 _29527_ (.A(_01283_),
    .Y(_03632_));
 sky130_fd_sc_hd__inv_2 _29528_ (.A(_01400_),
    .Y(_01402_));
 sky130_fd_sc_hd__inv_2 _29529_ (.A(_01334_),
    .Y(_01401_));
 sky130_fd_sc_hd__inv_2 _29530_ (.A(_01333_),
    .Y(_03636_));
 sky130_fd_sc_hd__inv_2 _29531_ (.A(_01348_),
    .Y(_03638_));
 sky130_fd_sc_hd__inv_2 _29532_ (.A(_01458_),
    .Y(_01460_));
 sky130_fd_sc_hd__inv_2 _29533_ (.A(_01399_),
    .Y(_01459_));
 sky130_fd_sc_hd__inv_2 _29534_ (.A(_01398_),
    .Y(_03642_));
 sky130_fd_sc_hd__inv_2 _29535_ (.A(_01408_),
    .Y(_03644_));
 sky130_fd_sc_hd__inv_2 _29536_ (.A(_01514_),
    .Y(_01516_));
 sky130_fd_sc_hd__inv_2 _29537_ (.A(_01457_),
    .Y(_01515_));
 sky130_fd_sc_hd__inv_2 _29538_ (.A(_01456_),
    .Y(_03648_));
 sky130_fd_sc_hd__inv_2 _29539_ (.A(_01466_),
    .Y(_03650_));
 sky130_fd_sc_hd__nor2_1 _29540_ (.A(_02983_),
    .B(net1140),
    .Y(_01537_));
 sky130_fd_sc_hd__inv_2 _29541_ (.A(_01572_),
    .Y(_01574_));
 sky130_fd_sc_hd__inv_2 _29542_ (.A(_01513_),
    .Y(_01573_));
 sky130_fd_sc_hd__inv_2 _29543_ (.A(_01512_),
    .Y(_03654_));
 sky130_fd_sc_hd__inv_2 _29544_ (.A(_01522_),
    .Y(_03656_));
 sky130_fd_sc_hd__inv_2 _29545_ (.A(_01626_),
    .Y(_01628_));
 sky130_fd_sc_hd__inv_2 _29546_ (.A(_01571_),
    .Y(_01627_));
 sky130_fd_sc_hd__inv_2 _29547_ (.A(_01570_),
    .Y(_03660_));
 sky130_fd_sc_hd__inv_2 _29548_ (.A(_01580_),
    .Y(_03662_));
 sky130_fd_sc_hd__inv_2 _29549_ (.A(_01678_),
    .Y(_01680_));
 sky130_fd_sc_hd__inv_2 _29550_ (.A(_01625_),
    .Y(_01679_));
 sky130_fd_sc_hd__inv_2 _29551_ (.A(_01624_),
    .Y(_03666_));
 sky130_fd_sc_hd__inv_2 _29552_ (.A(_01634_),
    .Y(_03668_));
 sky130_fd_sc_hd__inv_2 _29553_ (.A(_01674_),
    .Y(_01676_));
 sky130_fd_sc_hd__inv_2 _29554_ (.A(_01665_),
    .Y(_01731_));
 sky130_fd_sc_hd__inv_2 _29555_ (.A(_01737_),
    .Y(_02552_));
 sky130_fd_sc_hd__nor2_1 _29556_ (.A(net1718),
    .B(net1123),
    .Y(_01756_));
 sky130_fd_sc_hd__inv_2 _29557_ (.A(_01717_),
    .Y(_01777_));
 sky130_fd_sc_hd__inv_2 _29558_ (.A(_01786_),
    .Y(_02558_));
 sky130_fd_sc_hd__nor2_1 _29559_ (.A(net1121),
    .B(net1717),
    .Y(_01805_));
 sky130_fd_sc_hd__inv_2 _29560_ (.A(_01767_),
    .Y(_01825_));
 sky130_fd_sc_hd__inv_2 _29561_ (.A(_01834_),
    .Y(_02564_));
 sky130_fd_sc_hd__nor2_1 _29562_ (.A(net1141),
    .B(net1266),
    .Y(_01844_));
 sky130_fd_sc_hd__nor2_1 _29563_ (.A(net1212),
    .B(net3042),
    .Y(_01849_));
 sky130_fd_sc_hd__nor2_1 _29564_ (.A(net1718),
    .B(net1672),
    .Y(_01859_));
 sky130_fd_sc_hd__nor2_1 _29565_ (.A(net1323),
    .B(net1223),
    .Y(_01868_));
 sky130_fd_sc_hd__inv_2 _29566_ (.A(_01819_),
    .Y(_01878_));
 sky130_fd_sc_hd__inv_2 _29567_ (.A(_01887_),
    .Y(_02570_));
 sky130_fd_sc_hd__nor2_1 _29568_ (.A(net1140),
    .B(net1266),
    .Y(_01897_));
 sky130_fd_sc_hd__nor2_1 _29569_ (.A(net1129),
    .B(net1212),
    .Y(_01904_));
 sky130_fd_sc_hd__nor2_1 _29570_ (.A(_03011_),
    .B(net1115),
    .Y(_01918_));
 sky130_fd_sc_hd__nor2_1 _29571_ (.A(net1407),
    .B(net1108),
    .Y(_01867_));
 sky130_fd_sc_hd__inv_2 _29572_ (.A(_01872_),
    .Y(_01931_));
 sky130_fd_sc_hd__inv_2 _29573_ (.A(_01940_),
    .Y(_02576_));
 sky130_fd_sc_hd__nor2_1 _29574_ (.A(net1265),
    .B(net1138),
    .Y(_01950_));
 sky130_fd_sc_hd__inv_2 _29575_ (.A(_01925_),
    .Y(_01979_));
 sky130_fd_sc_hd__inv_2 _29576_ (.A(_01988_),
    .Y(_02582_));
 sky130_fd_sc_hd__nor2_1 _29577_ (.A(net1266),
    .B(net3042),
    .Y(_01998_));
 sky130_fd_sc_hd__inv_2 _29578_ (.A(_02035_),
    .Y(_02588_));
 sky130_fd_sc_hd__nor2_1 _29579_ (.A(net1129),
    .B(net1266),
    .Y(_02045_));
 sky130_fd_sc_hd__inv_2 _29580_ (.A(_02081_),
    .Y(_02594_));
 sky130_fd_sc_hd__nor2_1 _29581_ (.A(net1126),
    .B(net1266),
    .Y(_02091_));
 sky130_fd_sc_hd__inv_2 _29582_ (.A(_02120_),
    .Y(_02600_));
 sky130_fd_sc_hd__inv_2 _29583_ (.A(_02150_),
    .Y(_02607_));
 sky130_fd_sc_hd__nor2_1 _29584_ (.A(net1266),
    .B(net1123),
    .Y(_02160_));
 sky130_fd_sc_hd__inv_2 _29585_ (.A(_02183_),
    .Y(_02613_));
 sky130_fd_sc_hd__nor2_1 _29586_ (.A(net1127),
    .B(net1218),
    .Y(_02190_));
 sky130_fd_sc_hd__inv_2 _29587_ (.A(_02210_),
    .Y(_02620_));
 sky130_fd_sc_hd__nor2_1 _29588_ (.A(net1218),
    .B(net3044),
    .Y(_02217_));
 sky130_fd_sc_hd__inv_2 _29589_ (.A(_02244_),
    .Y(_02626_));
 sky130_fd_sc_hd__nor2_1 _29590_ (.A(net1218),
    .B(net1124),
    .Y(_02251_));
 sky130_fd_sc_hd__inv_2 _29591_ (.A(_02283_),
    .Y(_02632_));
 sky130_fd_sc_hd__nor2_1 _29592_ (.A(net1122),
    .B(net1218),
    .Y(_02290_));
 sky130_fd_sc_hd__inv_2 _29593_ (.A(_02317_),
    .Y(_02638_));
 sky130_fd_sc_hd__inv_2 _29594_ (.A(_02344_),
    .Y(_02645_));
 sky130_fd_sc_hd__nor2_1 _29595_ (.A(net1275),
    .B(_06005_),
    .Y(_02348_));
 sky130_fd_sc_hd__inv_2 _29596_ (.A(_02374_),
    .Y(_02651_));
 sky130_fd_sc_hd__inv_2 _29597_ (.A(_02404_),
    .Y(_02657_));
 sky130_fd_sc_hd__inv_2 _29598_ (.A(_02429_),
    .Y(_02663_));
 sky130_fd_sc_hd__inv_2 _29599_ (.A(_02454_),
    .Y(_02669_));
 sky130_fd_sc_hd__inv_2 _29600_ (.A(_02475_),
    .Y(_02675_));
 sky130_fd_sc_hd__inv_2 _29601_ (.A(_02490_),
    .Y(_02682_));
 sky130_fd_sc_hd__inv_2 _29602_ (.A(_02509_),
    .Y(_02688_));
 sky130_fd_sc_hd__inv_2 _29603_ (.A(_02517_),
    .Y(_02522_));
 sky130_fd_sc_hd__inv_2 _29604_ (.A(_02539_),
    .Y(_02696_));
 sky130_fd_sc_hd__inv_2 _29605_ (.A(\inst$top.soc.uart_0._phy.tx.lower.bitno[1] ),
    .Y(_02703_));
 sky130_fd_sc_hd__inv_2 _29606_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[1] ),
    .Y(_02707_));
 sky130_fd_sc_hd__inv_2 _29607_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[1] ),
    .Y(_02711_));
 sky130_fd_sc_hd__inv_2 _29608_ (.A(\inst$top.soc.uart_0._phy.rx.lower.bitno[1] ),
    .Y(_02715_));
 sky130_fd_sc_hd__inv_2 _29609_ (.A(\inst$top.soc.spiflash.ctrl.o_addr_count[1] ),
    .Y(_02724_));
 sky130_fd_sc_hd__inv_2 _29610_ (.A(\inst$top.soc.spiflash.ctrl.i_data_count[1] ),
    .Y(_02733_));
 sky130_fd_sc_hd__inv_2 _29611_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[1] ),
    .Y(_02740_));
 sky130_fd_sc_hd__inv_2 _29612_ (.A(\inst$top.soc.cpu.divider.divisor[31] ),
    .Y(_02751_));
 sky130_fd_sc_hd__inv_2 _29613_ (.A(\inst$top.soc.cpu.divider.divisor[30] ),
    .Y(_02754_));
 sky130_fd_sc_hd__inv_2 _29614_ (.A(\inst$top.soc.cpu.divider.divisor[29] ),
    .Y(_02757_));
 sky130_fd_sc_hd__inv_2 _29615_ (.A(\inst$top.soc.cpu.divider.divisor[28] ),
    .Y(_02760_));
 sky130_fd_sc_hd__inv_2 _29616_ (.A(\inst$top.soc.cpu.divider.divisor[27] ),
    .Y(_02763_));
 sky130_fd_sc_hd__inv_2 _29617_ (.A(\inst$top.soc.cpu.divider.divisor[26] ),
    .Y(_02766_));
 sky130_fd_sc_hd__inv_2 _29618_ (.A(\inst$top.soc.cpu.divider.divisor[25] ),
    .Y(_02769_));
 sky130_fd_sc_hd__inv_2 _29619_ (.A(\inst$top.soc.cpu.divider.divisor[24] ),
    .Y(_02772_));
 sky130_fd_sc_hd__inv_2 _29620_ (.A(\inst$top.soc.cpu.divider.divisor[23] ),
    .Y(_02775_));
 sky130_fd_sc_hd__inv_2 _29621_ (.A(\inst$top.soc.cpu.divider.divisor[22] ),
    .Y(_02778_));
 sky130_fd_sc_hd__inv_2 _29622_ (.A(\inst$top.soc.cpu.divider.divisor[21] ),
    .Y(_02781_));
 sky130_fd_sc_hd__inv_2 _29623_ (.A(\inst$top.soc.cpu.divider.divisor[20] ),
    .Y(_02784_));
 sky130_fd_sc_hd__inv_2 _29624_ (.A(\inst$top.soc.cpu.divider.divisor[19] ),
    .Y(_02787_));
 sky130_fd_sc_hd__inv_2 _29625_ (.A(\inst$top.soc.cpu.divider.divisor[18] ),
    .Y(_02790_));
 sky130_fd_sc_hd__inv_2 _29626_ (.A(\inst$top.soc.cpu.divider.divisor[17] ),
    .Y(_02793_));
 sky130_fd_sc_hd__inv_2 _29627_ (.A(\inst$top.soc.cpu.divider.divisor[16] ),
    .Y(_02796_));
 sky130_fd_sc_hd__inv_2 _29628_ (.A(\inst$top.soc.cpu.divider.divisor[15] ),
    .Y(_02799_));
 sky130_fd_sc_hd__inv_2 _29629_ (.A(\inst$top.soc.cpu.divider.divisor[14] ),
    .Y(_02802_));
 sky130_fd_sc_hd__inv_2 _29630_ (.A(\inst$top.soc.cpu.divider.divisor[13] ),
    .Y(_02805_));
 sky130_fd_sc_hd__inv_2 _29631_ (.A(\inst$top.soc.cpu.divider.divisor[12] ),
    .Y(_02808_));
 sky130_fd_sc_hd__inv_2 _29632_ (.A(\inst$top.soc.cpu.divider.divisor[11] ),
    .Y(_02811_));
 sky130_fd_sc_hd__inv_2 _29633_ (.A(\inst$top.soc.cpu.divider.divisor[10] ),
    .Y(_02814_));
 sky130_fd_sc_hd__inv_2 _29634_ (.A(\inst$top.soc.cpu.divider.divisor[9] ),
    .Y(_02817_));
 sky130_fd_sc_hd__inv_2 _29635_ (.A(\inst$top.soc.cpu.divider.divisor[8] ),
    .Y(_02820_));
 sky130_fd_sc_hd__inv_2 _29636_ (.A(\inst$top.soc.cpu.divider.divisor[7] ),
    .Y(_02823_));
 sky130_fd_sc_hd__inv_2 _29637_ (.A(\inst$top.soc.cpu.divider.divisor[6] ),
    .Y(_02826_));
 sky130_fd_sc_hd__inv_2 _29638_ (.A(\inst$top.soc.cpu.divider.divisor[5] ),
    .Y(_02829_));
 sky130_fd_sc_hd__inv_2 _29639_ (.A(\inst$top.soc.cpu.divider.divisor[4] ),
    .Y(_02832_));
 sky130_fd_sc_hd__inv_2 _29640_ (.A(\inst$top.soc.cpu.divider.divisor[3] ),
    .Y(_02835_));
 sky130_fd_sc_hd__inv_2 _29641_ (.A(\inst$top.soc.cpu.divider.divisor[2] ),
    .Y(_02838_));
 sky130_fd_sc_hd__inv_2 _29642_ (.A(\inst$top.soc.cpu.divider.divisor[1] ),
    .Y(_02541_));
 sky130_fd_sc_hd__inv_2 _29643_ (.A(\inst$top.soc.cpu.divider.quotient[1] ),
    .Y(_02847_));
 sky130_fd_sc_hd__inv_2 _29644_ (.A(\inst$top.soc.cpu.divider.remainder[1] ),
    .Y(_02854_));
 sky130_fd_sc_hd__inv_2 _29645_ (.A(\inst$top.soc.cpu.divider.timer[1] ),
    .Y(_02858_));
 sky130_fd_sc_hd__inv_2 _29646_ (.A(\inst$top.soc.cpu.d.sink__payload$6.branch_predict_taken ),
    .Y(_02864_));
 sky130_fd_sc_hd__inv_2 _29647_ (.A(\inst$top.soc.uart_0._phy.rx.lower.fsm_state[1] ),
    .Y(_02878_));
 sky130_fd_sc_hd__inv_2 _29648_ (.A(_00193_),
    .Y(_03372_));
 sky130_fd_sc_hd__inv_2 _29649_ (.A(_00203_),
    .Y(_03376_));
 sky130_fd_sc_hd__inv_2 _29650_ (.A(_00197_),
    .Y(_03378_));
 sky130_fd_sc_hd__inv_2 _29651_ (.A(_00267_),
    .Y(_03400_));
 sky130_fd_sc_hd__inv_2 _29652_ (.A(_00293_),
    .Y(_03407_));
 sky130_fd_sc_hd__inv_2 _29653_ (.A(_00297_),
    .Y(_03410_));
 sky130_fd_sc_hd__inv_2 _29654_ (.A(_00328_),
    .Y(_03417_));
 sky130_fd_sc_hd__nor2_1 _29655_ (.A(net1693),
    .B(_03011_),
    .Y(_00380_));
 sky130_fd_sc_hd__inv_2 _29656_ (.A(_00419_),
    .Y(_03428_));
 sky130_fd_sc_hd__inv_2 _29657_ (.A(_00388_),
    .Y(_03429_));
 sky130_fd_sc_hd__inv_2 _29658_ (.A(_00449_),
    .Y(_03437_));
 sky130_fd_sc_hd__inv_2 _29659_ (.A(_00453_),
    .Y(_00454_));
 sky130_fd_sc_hd__inv_2 _29660_ (.A(_00478_),
    .Y(_03449_));
 sky130_fd_sc_hd__inv_2 _29661_ (.A(_00484_),
    .Y(_03453_));
 sky130_fd_sc_hd__nor2_1 _29662_ (.A(net1402),
    .B(_05907_),
    .Y(_00498_));
 sky130_fd_sc_hd__inv_2 _29663_ (.A(_00521_),
    .Y(_03462_));
 sky130_fd_sc_hd__nor2_1 _29664_ (.A(net1323),
    .B(net1158),
    .Y(_00530_));
 sky130_fd_sc_hd__nor2_1 _29665_ (.A(net1402),
    .B(net1156),
    .Y(_00539_));
 sky130_fd_sc_hd__inv_2 _29666_ (.A(_00564_),
    .Y(_03474_));
 sky130_fd_sc_hd__inv_2 _29667_ (.A(_00570_),
    .Y(_03479_));
 sky130_fd_sc_hd__nor2_1 _29668_ (.A(net1402),
    .B(_05912_),
    .Y(_00581_));
 sky130_fd_sc_hd__inv_2 _29669_ (.A(_00609_),
    .Y(_03485_));
 sky130_fd_sc_hd__inv_2 _29670_ (.A(_00614_),
    .Y(_03489_));
 sky130_fd_sc_hd__nor2_1 _29671_ (.A(net1399),
    .B(net1151),
    .Y(_00632_));
 sky130_fd_sc_hd__inv_2 _29672_ (.A(_00659_),
    .Y(_03494_));
 sky130_fd_sc_hd__inv_2 _29673_ (.A(_00677_),
    .Y(_03499_));
 sky130_fd_sc_hd__nor2_1 _29674_ (.A(net1401),
    .B(net1148),
    .Y(_00680_));
 sky130_fd_sc_hd__inv_2 _29675_ (.A(_00707_),
    .Y(_03506_));
 sky130_fd_sc_hd__inv_2 _29676_ (.A(_00716_),
    .Y(_00726_));
 sky130_fd_sc_hd__nor2_1 _29677_ (.A(net1401),
    .B(net1146),
    .Y(_00730_));
 sky130_fd_sc_hd__inv_2 _29678_ (.A(_00755_),
    .Y(_03520_));
 sky130_fd_sc_hd__nor2_1 _29679_ (.A(net1694),
    .B(net1212),
    .Y(_00759_));
 sky130_fd_sc_hd__inv_2 _29680_ (.A(_00768_),
    .Y(_03523_));
 sky130_fd_sc_hd__nor2_1 _29681_ (.A(net1401),
    .B(net1144),
    .Y(_00784_));
 sky130_fd_sc_hd__inv_2 _29682_ (.A(_00810_),
    .Y(_03531_));
 sky130_fd_sc_hd__inv_2 _29683_ (.A(_00820_),
    .Y(_03535_));
 sky130_fd_sc_hd__nor2_1 _29684_ (.A(_03011_),
    .B(_05908_),
    .Y(_00825_));
 sky130_fd_sc_hd__nor2_1 _29685_ (.A(net1401),
    .B(net1141),
    .Y(_00838_));
 sky130_fd_sc_hd__inv_2 _29686_ (.A(_00780_),
    .Y(_00858_));
 sky130_fd_sc_hd__inv_2 _29687_ (.A(_00867_),
    .Y(_03544_));
 sky130_fd_sc_hd__inv_2 _29688_ (.A(_00876_),
    .Y(_03550_));
 sky130_fd_sc_hd__nor2_1 _29689_ (.A(net1401),
    .B(net1140),
    .Y(_00895_));
 sky130_fd_sc_hd__inv_2 _29690_ (.A(_00834_),
    .Y(_00915_));
 sky130_fd_sc_hd__inv_2 _29691_ (.A(_00923_),
    .Y(_03556_));
 sky130_fd_sc_hd__nor2_1 _29692_ (.A(net1694),
    .B(net1266),
    .Y(_00927_));
 sky130_fd_sc_hd__inv_2 _29693_ (.A(_00934_),
    .Y(_03561_));
 sky130_fd_sc_hd__nor2_1 _29694_ (.A(net1401),
    .B(net1138),
    .Y(_00950_));
 sky130_fd_sc_hd__inv_2 _29695_ (.A(_00888_),
    .Y(_00970_));
 sky130_fd_sc_hd__inv_2 _29696_ (.A(_00977_),
    .Y(_03568_));
 sky130_fd_sc_hd__inv_2 _29697_ (.A(_00983_),
    .Y(_03571_));
 sky130_fd_sc_hd__nor2_1 _29698_ (.A(net1156),
    .B(net1718),
    .Y(_00994_));
 sky130_fd_sc_hd__nor2_1 _29699_ (.A(net1401),
    .B(net1136),
    .Y(_01010_));
 sky130_fd_sc_hd__inv_2 _29700_ (.A(_00945_),
    .Y(_01030_));
 sky130_fd_sc_hd__inv_2 _29701_ (.A(_01036_),
    .Y(_03580_));
 sky130_fd_sc_hd__nor2_1 _29702_ (.A(net1694),
    .B(_19946_),
    .Y(_03584_));
 sky130_fd_sc_hd__inv_2 _29703_ (.A(_01041_),
    .Y(_03587_));
 sky130_fd_sc_hd__nor2_1 _29704_ (.A(net1152),
    .B(net1718),
    .Y(_01055_));
 sky130_fd_sc_hd__inv_2 _29705_ (.A(_01005_),
    .Y(_01091_));
 sky130_fd_sc_hd__inv_2 _29706_ (.A(_01097_),
    .Y(_03593_));
 sky130_fd_sc_hd__inv_2 _29707_ (.A(_01102_),
    .Y(_03597_));
 sky130_fd_sc_hd__nor2_1 _29708_ (.A(net1150),
    .B(net1717),
    .Y(_01119_));
 sky130_fd_sc_hd__inv_2 _29709_ (.A(_01066_),
    .Y(_01157_));
 sky130_fd_sc_hd__inv_2 _29710_ (.A(_01163_),
    .Y(_03602_));
 sky130_fd_sc_hd__inv_2 _29711_ (.A(_01130_),
    .Y(_01219_));
 sky130_fd_sc_hd__inv_2 _29712_ (.A(_01225_),
    .Y(_03613_));
 sky130_fd_sc_hd__nor2_1 _29713_ (.A(net1146),
    .B(net1717),
    .Y(_01245_));
 sky130_fd_sc_hd__inv_2 _29714_ (.A(_01284_),
    .Y(_03625_));
 sky130_fd_sc_hd__inv_2 _29715_ (.A(_01255_),
    .Y(_01338_));
 sky130_fd_sc_hd__inv_2 _29716_ (.A(_01280_),
    .Y(_01343_));
 sky130_fd_sc_hd__inv_2 _29717_ (.A(_01349_),
    .Y(_03633_));
 sky130_fd_sc_hd__nor2_1 _29718_ (.A(net1141),
    .B(net1717),
    .Y(_01369_));
 sky130_fd_sc_hd__inv_2 _29719_ (.A(_01311_),
    .Y(_01403_));
 sky130_fd_sc_hd__inv_2 _29720_ (.A(_01409_),
    .Y(_03639_));
 sky130_fd_sc_hd__inv_2 _29721_ (.A(_01379_),
    .Y(_01461_));
 sky130_fd_sc_hd__inv_2 _29722_ (.A(_01467_),
    .Y(_03645_));
 sky130_fd_sc_hd__nor2_1 _29723_ (.A(net1717),
    .B(net1138),
    .Y(_01486_));
 sky130_fd_sc_hd__inv_2 _29724_ (.A(_01436_),
    .Y(_01517_));
 sky130_fd_sc_hd__inv_2 _29725_ (.A(_01523_),
    .Y(_03651_));
 sky130_fd_sc_hd__nor2_1 _29726_ (.A(_20003_),
    .B(net1142),
    .Y(_01538_));
 sky130_fd_sc_hd__nor2_1 _29727_ (.A(net1717),
    .B(net1136),
    .Y(_01545_));
 sky130_fd_sc_hd__nor2_1 _29728_ (.A(net1171),
    .B(net1221),
    .Y(_01565_));
 sky130_fd_sc_hd__inv_2 _29729_ (.A(_01496_),
    .Y(_01575_));
 sky130_fd_sc_hd__inv_2 _29730_ (.A(_01581_),
    .Y(_03657_));
 sky130_fd_sc_hd__nor2_1 _29731_ (.A(net1131),
    .B(net1717),
    .Y(_01600_));
 sky130_fd_sc_hd__inv_2 _29732_ (.A(_01556_),
    .Y(_01629_));
 sky130_fd_sc_hd__inv_2 _29733_ (.A(_01635_),
    .Y(_03663_));
 sky130_fd_sc_hd__nor2_1 _29734_ (.A(net1126),
    .B(net1717),
    .Y(_01654_));
 sky130_fd_sc_hd__inv_2 _29735_ (.A(_01612_),
    .Y(_01681_));
 sky130_fd_sc_hd__inv_2 _29736_ (.A(_01687_),
    .Y(_03669_));
 sky130_fd_sc_hd__nor2_1 _29737_ (.A(net1717),
    .B(net1677),
    .Y(_01706_));
 sky130_fd_sc_hd__inv_2 _29738_ (.A(_02550_),
    .Y(_01734_));
 sky130_fd_sc_hd__inv_2 _29739_ (.A(_02556_),
    .Y(_01783_));
 sky130_fd_sc_hd__inv_2 _29740_ (.A(_03441_),
    .Y(_00450_));
 sky130_fd_sc_hd__inv_2 _29741_ (.A(_03452_),
    .Y(_00479_));
 sky130_fd_sc_hd__inv_2 _29742_ (.A(_03472_),
    .Y(_00558_));
 sky130_fd_sc_hd__inv_2 _29743_ (.A(_03483_),
    .Y(_00604_));
 sky130_fd_sc_hd__inv_2 _29744_ (.A(_03492_),
    .Y(_00654_));
 sky130_fd_sc_hd__inv_2 _29745_ (.A(_03504_),
    .Y(_00702_));
 sky130_fd_sc_hd__inv_2 _29746_ (.A(_03518_),
    .Y(_00751_));
 sky130_fd_sc_hd__inv_2 _29747_ (.A(_03529_),
    .Y(_00806_));
 sky130_fd_sc_hd__inv_2 _29748_ (.A(_03542_),
    .Y(_00863_));
 sky130_fd_sc_hd__inv_2 _29749_ (.A(_03554_),
    .Y(_00920_));
 sky130_fd_sc_hd__inv_2 _29750_ (.A(_03566_),
    .Y(_00974_));
 sky130_fd_sc_hd__inv_2 _29751_ (.A(_03578_),
    .Y(_01033_));
 sky130_fd_sc_hd__inv_2 _29752_ (.A(_03591_),
    .Y(_01094_));
 sky130_fd_sc_hd__inv_2 _29753_ (.A(_03600_),
    .Y(_01160_));
 sky130_fd_sc_hd__inv_2 _29754_ (.A(_03611_),
    .Y(_01222_));
 sky130_fd_sc_hd__inv_2 _29755_ (.A(_03621_),
    .Y(_01235_));
 sky130_fd_sc_hd__inv_2 _29756_ (.A(_03623_),
    .Y(_01281_));
 sky130_fd_sc_hd__inv_2 _29757_ (.A(_03631_),
    .Y(_01290_));
 sky130_fd_sc_hd__inv_2 _29758_ (.A(_03637_),
    .Y(_01406_));
 sky130_fd_sc_hd__inv_2 _29759_ (.A(_03643_),
    .Y(_01464_));
 sky130_fd_sc_hd__inv_2 _29760_ (.A(_03649_),
    .Y(_01520_));
 sky130_fd_sc_hd__inv_2 _29761_ (.A(_03655_),
    .Y(_01578_));
 sky130_fd_sc_hd__inv_2 _29762_ (.A(_03661_),
    .Y(_01632_));
 sky130_fd_sc_hd__inv_2 _29763_ (.A(_03667_),
    .Y(_01684_));
 sky130_fd_sc_hd__inv_2 _29764_ (.A(_02562_),
    .Y(_01831_));
 sky130_fd_sc_hd__inv_2 _29765_ (.A(_02568_),
    .Y(_01884_));
 sky130_fd_sc_hd__inv_2 _29766_ (.A(_02574_),
    .Y(_01937_));
 sky130_fd_sc_hd__inv_2 _29767_ (.A(_02580_),
    .Y(_01985_));
 sky130_fd_sc_hd__inv_2 _29768_ (.A(_02586_),
    .Y(_02032_));
 sky130_fd_sc_hd__inv_2 _29769_ (.A(_02592_),
    .Y(_02078_));
 sky130_fd_sc_hd__inv_2 _29770_ (.A(_02598_),
    .Y(_02117_));
 sky130_fd_sc_hd__inv_2 _29771_ (.A(_02605_),
    .Y(_02147_));
 sky130_fd_sc_hd__inv_2 _29772_ (.A(_02611_),
    .Y(_02180_));
 sky130_fd_sc_hd__inv_2 _29773_ (.A(_02618_),
    .Y(_02207_));
 sky130_fd_sc_hd__inv_2 _29774_ (.A(_02624_),
    .Y(_02241_));
 sky130_fd_sc_hd__inv_2 _29775_ (.A(_02630_),
    .Y(_02280_));
 sky130_fd_sc_hd__inv_2 _29776_ (.A(_02636_),
    .Y(_02314_));
 sky130_fd_sc_hd__inv_2 _29777_ (.A(_02643_),
    .Y(_02341_));
 sky130_fd_sc_hd__inv_2 _29778_ (.A(_02649_),
    .Y(_02371_));
 sky130_fd_sc_hd__inv_2 _29779_ (.A(_02655_),
    .Y(_02401_));
 sky130_fd_sc_hd__inv_2 _29780_ (.A(_02661_),
    .Y(_02426_));
 sky130_fd_sc_hd__inv_2 _29781_ (.A(_02667_),
    .Y(_02451_));
 sky130_fd_sc_hd__inv_2 _29782_ (.A(_02673_),
    .Y(_02472_));
 sky130_fd_sc_hd__inv_2 _29783_ (.A(_02680_),
    .Y(_02487_));
 sky130_fd_sc_hd__inv_2 _29784_ (.A(_02686_),
    .Y(_02506_));
 sky130_fd_sc_hd__inv_2 _29785_ (.A(_02694_),
    .Y(_02535_));
 sky130_fd_sc_hd__inv_2 _29786_ (.A(_03373_),
    .Y(_00202_));
 sky130_fd_sc_hd__inv_2 _29787_ (.A(_03399_),
    .Y(_00265_));
 sky130_fd_sc_hd__inv_2 _29788_ (.A(_03469_),
    .Y(_00560_));
 sky130_fd_sc_hd__inv_2 _29789_ (.A(_03540_),
    .Y(_00862_));
 sky130_fd_sc_hd__inv_2 _29790_ (.A(_03564_),
    .Y(_00947_));
 sky130_fd_sc_hd__inv_2 _29791_ (.A(_03576_),
    .Y(_01007_));
 sky130_fd_sc_hd__inv_2 _29792_ (.A(_03459_),
    .Y(_00559_));
 sky130_fd_sc_hd__inv_2 _29793_ (.A(_03468_),
    .Y(_00605_));
 sky130_fd_sc_hd__inv_2 _29794_ (.A(_03513_),
    .Y(_00779_));
 sky130_fd_sc_hd__inv_2 _29795_ (.A(_03524_),
    .Y(_00833_));
 sky130_fd_sc_hd__inv_2 _29796_ (.A(_03526_),
    .Y(_00861_));
 sky130_fd_sc_hd__inv_2 _29797_ (.A(_03536_),
    .Y(_00887_));
 sky130_fd_sc_hd__inv_2 _29798_ (.A(_03539_),
    .Y(_00918_));
 sky130_fd_sc_hd__inv_2 _29799_ (.A(_03551_),
    .Y(_00944_));
 sky130_fd_sc_hd__inv_2 _29800_ (.A(_03552_),
    .Y(_00946_));
 sky130_fd_sc_hd__inv_2 _29801_ (.A(_03559_),
    .Y(_00990_));
 sky130_fd_sc_hd__inv_2 _29802_ (.A(_03562_),
    .Y(_01004_));
 sky130_fd_sc_hd__inv_2 _29803_ (.A(_03563_),
    .Y(_01006_));
 sky130_fd_sc_hd__inv_2 _29804_ (.A(_03572_),
    .Y(_01048_));
 sky130_fd_sc_hd__inv_2 _29805_ (.A(_03575_),
    .Y(_01067_));
 sky130_fd_sc_hd__inv_2 _29806_ (.A(_03585_),
    .Y(_01106_));
 sky130_fd_sc_hd__inv_2 _29807_ (.A(_03588_),
    .Y(_01114_));
 sky130_fd_sc_hd__inv_2 _29808_ (.A(_03607_),
    .Y(_01234_));
 sky130_fd_sc_hd__inv_2 _29809_ (.A(_03609_),
    .Y(_01242_));
 sky130_fd_sc_hd__inv_2 _29810_ (.A(_03618_),
    .Y(_01289_));
 sky130_fd_sc_hd__inv_2 _29811_ (.A(_03620_),
    .Y(_01294_));
 sky130_fd_sc_hd__o21ai_0 _29812_ (.A1(_20302_),
    .A2(_06036_),
    .B1(net2821),
    .Y(_09354_));
 sky130_fd_sc_hd__nand2_1 _29813_ (.A(_20289_),
    .B(_20291_),
    .Y(_09355_));
 sky130_fd_sc_hd__nand2_1 _29814_ (.A(_09354_),
    .B(_09355_),
    .Y(_09356_));
 sky130_fd_sc_hd__o21ai_0 _29815_ (.A1(_20292_),
    .A2(_20293_),
    .B1(net2821),
    .Y(_09357_));
 sky130_fd_sc_hd__nand2_1 _29816_ (.A(_20299_),
    .B(_20291_),
    .Y(_09358_));
 sky130_fd_sc_hd__nand2_1 _29817_ (.A(_09357_),
    .B(_09358_),
    .Y(_09359_));
 sky130_fd_sc_hd__nand3_1 _29818_ (.A(_09356_),
    .B(_09359_),
    .C(_20307_),
    .Y(_09360_));
 sky130_fd_sc_hd__inv_1 _29819_ (.A(\inst$top.soc.cpu.sink__payload$6[39] ),
    .Y(_09361_));
 sky130_fd_sc_hd__inv_1 _29820_ (.A(\inst$top.soc.cpu.sink__payload$6[63] ),
    .Y(_09362_));
 sky130_fd_sc_hd__nor2_1 _29821_ (.A(_20305_),
    .B(_06036_),
    .Y(_09363_));
 sky130_fd_sc_hd__inv_1 _29822_ (.A(_09363_),
    .Y(_09364_));
 sky130_fd_sc_hd__o22ai_1 _29823_ (.A1(_09361_),
    .A2(_20296_),
    .B1(_09362_),
    .B2(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__a221oi_1 _29824_ (.A1(net2687),
    .A2(_20285_),
    .B1(_09360_),
    .B2(\inst$top.soc.cpu.sink__payload$6[63] ),
    .C1(_09365_),
    .Y(_09366_));
 sky130_fd_sc_hd__inv_2 _29825_ (.A(_09366_),
    .Y(\inst$top.soc.cpu.csrf.d_addr[11] ));
 sky130_fd_sc_hd__o21a_1 _29826_ (.A1(_06037_),
    .A2(_09360_),
    .B1(\inst$top.soc.cpu.sink__payload$6[63] ),
    .X(_09367_));
 sky130_fd_sc_hd__a21oi_1 _29828_ (.A1(\inst$top.soc.cpu.sink__payload$6[44] ),
    .A2(net1191),
    .B1(_09367_),
    .Y(_09369_));
 sky130_fd_sc_hd__inv_2 _29829_ (.A(_09369_),
    .Y(\inst$top.soc.cpu.d_offset[12] ));
 sky130_fd_sc_hd__a21oi_1 _29830_ (.A1(\inst$top.soc.cpu.sink__payload$6[45] ),
    .A2(net1191),
    .B1(_09367_),
    .Y(_09370_));
 sky130_fd_sc_hd__inv_2 _29831_ (.A(_09370_),
    .Y(\inst$top.soc.cpu.d_offset[13] ));
 sky130_fd_sc_hd__a21oi_1 _29833_ (.A1(net2820),
    .A2(net1191),
    .B1(_09367_),
    .Y(_09372_));
 sky130_fd_sc_hd__inv_2 _29834_ (.A(_09372_),
    .Y(\inst$top.soc.cpu.d_offset[14] ));
 sky130_fd_sc_hd__a21oi_1 _29835_ (.A1(net2767),
    .A2(net1191),
    .B1(_09367_),
    .Y(_09373_));
 sky130_fd_sc_hd__inv_2 _29836_ (.A(_09373_),
    .Y(\inst$top.soc.cpu.d_offset[15] ));
 sky130_fd_sc_hd__a21oi_1 _29837_ (.A1(net2724),
    .A2(net1191),
    .B1(_09367_),
    .Y(_09374_));
 sky130_fd_sc_hd__inv_2 _29838_ (.A(_09374_),
    .Y(\inst$top.soc.cpu.d_offset[16] ));
 sky130_fd_sc_hd__a21oi_1 _29839_ (.A1(net2703),
    .A2(net1191),
    .B1(_09367_),
    .Y(_09375_));
 sky130_fd_sc_hd__inv_2 _29840_ (.A(_09375_),
    .Y(\inst$top.soc.cpu.d_offset[17] ));
 sky130_fd_sc_hd__a21oi_1 _29841_ (.A1(net2696),
    .A2(net1191),
    .B1(_09367_),
    .Y(_09376_));
 sky130_fd_sc_hd__inv_2 _29842_ (.A(_09376_),
    .Y(\inst$top.soc.cpu.d_offset[18] ));
 sky130_fd_sc_hd__a21oi_1 _29843_ (.A1(net2690),
    .A2(net1191),
    .B1(_09367_),
    .Y(_09377_));
 sky130_fd_sc_hd__inv_2 _29844_ (.A(_09377_),
    .Y(\inst$top.soc.cpu.d_offset[19] ));
 sky130_fd_sc_hd__inv_1 _29845_ (.A(_06046_),
    .Y(_09378_));
 sky130_fd_sc_hd__nand2_1 _29846_ (.A(_09378_),
    .B(\inst$top.soc.cpu.sink__payload$6[63] ),
    .Y(_09379_));
 sky130_fd_sc_hd__o21ai_1 _29847_ (.A1(net2465),
    .A2(_20311_),
    .B1(_09379_),
    .Y(\inst$top.soc.cpu.d_offset[20] ));
 sky130_fd_sc_hd__o21ai_2 _29848_ (.A1(_20261_),
    .A2(_20311_),
    .B1(_09379_),
    .Y(\inst$top.soc.cpu.d_offset[21] ));
 sky130_fd_sc_hd__o21ai_1 _29849_ (.A1(net2460),
    .A2(_20311_),
    .B1(_09379_),
    .Y(\inst$top.soc.cpu.d_offset[22] ));
 sky130_fd_sc_hd__inv_1 _29850_ (.A(_20311_),
    .Y(_09380_));
 sky130_fd_sc_hd__inv_1 _29851_ (.A(_09379_),
    .Y(_09381_));
 sky130_fd_sc_hd__a21oi_1 _29852_ (.A1(net2597),
    .A2(_09380_),
    .B1(_09381_),
    .Y(_09382_));
 sky130_fd_sc_hd__inv_2 _29853_ (.A(_09382_),
    .Y(\inst$top.soc.cpu.d_offset[23] ));
 sky130_fd_sc_hd__a21oi_1 _29854_ (.A1(net2590),
    .A2(_09380_),
    .B1(_09381_),
    .Y(_09383_));
 sky130_fd_sc_hd__inv_2 _29855_ (.A(_09383_),
    .Y(\inst$top.soc.cpu.d_offset[24] ));
 sky130_fd_sc_hd__a21oi_1 _29856_ (.A1(\inst$top.soc.cpu.sink__payload$6[57] ),
    .A2(_09380_),
    .B1(_09381_),
    .Y(_09384_));
 sky130_fd_sc_hd__inv_2 _29857_ (.A(_09384_),
    .Y(\inst$top.soc.cpu.d_offset[25] ));
 sky130_fd_sc_hd__a21oi_1 _29858_ (.A1(\inst$top.soc.cpu.sink__payload$6[58] ),
    .A2(_09380_),
    .B1(_09381_),
    .Y(_09385_));
 sky130_fd_sc_hd__inv_2 _29859_ (.A(_09385_),
    .Y(\inst$top.soc.cpu.d_offset[26] ));
 sky130_fd_sc_hd__a21oi_1 _29860_ (.A1(\inst$top.soc.cpu.sink__payload$6[59] ),
    .A2(_09380_),
    .B1(_09381_),
    .Y(_09386_));
 sky130_fd_sc_hd__inv_2 _29861_ (.A(_09386_),
    .Y(\inst$top.soc.cpu.d_offset[27] ));
 sky130_fd_sc_hd__a21oi_1 _29862_ (.A1(\inst$top.soc.cpu.sink__payload$6[60] ),
    .A2(_09380_),
    .B1(_09381_),
    .Y(_09387_));
 sky130_fd_sc_hd__inv_2 _29863_ (.A(_09387_),
    .Y(\inst$top.soc.cpu.d_offset[28] ));
 sky130_fd_sc_hd__a21oi_1 _29864_ (.A1(\inst$top.soc.cpu.sink__payload$6[61] ),
    .A2(_09380_),
    .B1(_09381_),
    .Y(_09388_));
 sky130_fd_sc_hd__inv_2 _29865_ (.A(_09388_),
    .Y(\inst$top.soc.cpu.d_offset[29] ));
 sky130_fd_sc_hd__a21oi_1 _29866_ (.A1(\inst$top.soc.cpu.sink__payload$6[62] ),
    .A2(_09380_),
    .B1(_09381_),
    .Y(_09389_));
 sky130_fd_sc_hd__inv_2 _29867_ (.A(_09389_),
    .Y(\inst$top.soc.cpu.d_offset[30] ));
 sky130_fd_sc_hd__nor2_1 _29872_ (.A(\inst$top.soc.cpu.a.source__valid ),
    .B(net666),
    .Y(_09394_));
 sky130_fd_sc_hd__nor2_2 _29873_ (.A(net2938),
    .B(_09394_),
    .Y(_03672_));
 sky130_fd_sc_hd__inv_2 _29880_ (.A(net2957),
    .Y(_09401_));
 sky130_fd_sc_hd__o21ai_0 _29883_ (.A1(\inst$top.soc.cpu.csrf.bank_300_m_select ),
    .A2(net2251),
    .B1(net2085),
    .Y(_09404_));
 sky130_fd_sc_hd__a21oi_1 _29884_ (.A1(_20432_),
    .A2(net2251),
    .B1(_09404_),
    .Y(_03673_));
 sky130_fd_sc_hd__inv_2 _29885_ (.A(net2237),
    .Y(_09405_));
 sky130_fd_sc_hd__nand2_1 _29888_ (.A(net1883),
    .B(\inst$top.soc.cpu.csrf.bank_300_w_select ),
    .Y(_09408_));
 sky130_fd_sc_hd__nand2_1 _29891_ (.A(net2220),
    .B(\inst$top.soc.cpu.csrf.bank_300_m_select ),
    .Y(_09411_));
 sky130_fd_sc_hd__a21oi_1 _29893_ (.A1(_09408_),
    .A2(_09411_),
    .B1(net2957),
    .Y(_03674_));
 sky130_fd_sc_hd__nand2_4 _29894_ (.A(_20356_),
    .B(net792),
    .Y(_09413_));
 sky130_fd_sc_hd__clkinv_1 _29895_ (.A(_20369_),
    .Y(_09414_));
 sky130_fd_sc_hd__nand2_4 _29896_ (.A(net665),
    .B(net755),
    .Y(_09415_));
 sky130_fd_sc_hd__nand2_1 _29899_ (.A(net645),
    .B(\inst$top.soc.cpu.csrf.bank_300_x_select ),
    .Y(_09418_));
 sky130_fd_sc_hd__nand4_1 _29902_ (.A(\inst$top.soc.cpu.csrf.d_addr[9] ),
    .B(\inst$top.soc.cpu.sink__payload$6[60] ),
    .C(_06049_),
    .D(_06051_),
    .Y(_09421_));
 sky130_fd_sc_hd__nor2_1 _29903_ (.A(\inst$top.soc.cpu.csrf.d_addr[11] ),
    .B(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__nand3_1 _29904_ (.A(net664),
    .B(net754),
    .C(_09422_),
    .Y(_09423_));
 sky130_fd_sc_hd__a21oi_4 _29905_ (.A1(_09418_),
    .A2(_09423_),
    .B1(net2953),
    .Y(_03675_));
 sky130_fd_sc_hd__nand2_1 _29909_ (.A(net684),
    .B(net792),
    .Y(_09427_));
 sky130_fd_sc_hd__nand2_1 _29910_ (.A(net1904),
    .B(\inst$top.soc.cpu.d.source__valid ),
    .Y(_09428_));
 sky130_fd_sc_hd__a21oi_4 _29911_ (.A1(_09427_),
    .A2(_09428_),
    .B1(net2954),
    .Y(_03676_));
 sky130_fd_sc_hd__nand2_1 _29912_ (.A(net1159),
    .B(net1158),
    .Y(_09429_));
 sky130_fd_sc_hd__nor2_1 _29913_ (.A(net1351),
    .B(net1356),
    .Y(_09430_));
 sky130_fd_sc_hd__inv_1 _29914_ (.A(_09430_),
    .Y(_09431_));
 sky130_fd_sc_hd__nand3_1 _29915_ (.A(_05900_),
    .B(_02844_),
    .C(net1366),
    .Y(_09432_));
 sky130_fd_sc_hd__nor2_2 _29916_ (.A(_09431_),
    .B(_09432_),
    .Y(_09433_));
 sky130_fd_sc_hd__inv_1 _29917_ (.A(_09433_),
    .Y(_09434_));
 sky130_fd_sc_hd__nor2_1 _29918_ (.A(_09429_),
    .B(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__nor4_1 _29919_ (.A(net1303),
    .B(net1299),
    .C(net1295),
    .D(net1289),
    .Y(_09436_));
 sky130_fd_sc_hd__nor2_1 _29920_ (.A(net1341),
    .B(net1337),
    .Y(_09437_));
 sky130_fd_sc_hd__nor2_1 _29921_ (.A(net1331),
    .B(net1327),
    .Y(_09438_));
 sky130_fd_sc_hd__nand2_1 _29922_ (.A(_09437_),
    .B(_09438_),
    .Y(_09439_));
 sky130_fd_sc_hd__nor2_1 _29923_ (.A(net1312),
    .B(net1308),
    .Y(_09440_));
 sky130_fd_sc_hd__nand3_1 _29924_ (.A(_09440_),
    .B(net1150),
    .C(net1148),
    .Y(_09441_));
 sky130_fd_sc_hd__nor2_1 _29925_ (.A(_09439_),
    .B(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__nor2_1 _29926_ (.A(net1281),
    .B(net1286),
    .Y(_09443_));
 sky130_fd_sc_hd__nand3_1 _29927_ (.A(net1678),
    .B(_09443_),
    .C(net1124),
    .Y(_09444_));
 sky130_fd_sc_hd__inv_1 _29928_ (.A(_09444_),
    .Y(_09445_));
 sky130_fd_sc_hd__nand4_1 _29929_ (.A(_09435_),
    .B(_09436_),
    .C(_09442_),
    .D(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__inv_1 _29930_ (.A(net2842),
    .Y(_09447_));
 sky130_fd_sc_hd__nor2_1 _29931_ (.A(\inst$top.soc.cpu.sink__payload$12[143] ),
    .B(_09447_),
    .Y(_09448_));
 sky130_fd_sc_hd__inv_1 _29932_ (.A(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__nor2_2 _29933_ (.A(_09449_),
    .B(net1222),
    .Y(_09450_));
 sky130_fd_sc_hd__nand2_1 _29935_ (.A(_09446_),
    .B(net1044),
    .Y(_09452_));
 sky130_fd_sc_hd__nand2_1 _29936_ (.A(_09452_),
    .B(net1122),
    .Y(_09453_));
 sky130_fd_sc_hd__nand3_1 _29937_ (.A(_09446_),
    .B(net1272),
    .C(net1044),
    .Y(_09454_));
 sky130_fd_sc_hd__nand2_1 _29938_ (.A(_09453_),
    .B(_09454_),
    .Y(_09455_));
 sky130_fd_sc_hd__nor2_1 _29939_ (.A(net1303),
    .B(net1299),
    .Y(_09456_));
 sky130_fd_sc_hd__nand2_1 _29940_ (.A(_09440_),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__inv_1 _29941_ (.A(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__nor2_1 _29942_ (.A(net1295),
    .B(net1289),
    .Y(_09459_));
 sky130_fd_sc_hd__nand3_1 _29943_ (.A(_09458_),
    .B(_09443_),
    .C(_09459_),
    .Y(_09460_));
 sky130_fd_sc_hd__nand3_1 _29944_ (.A(_09438_),
    .B(net1150),
    .C(net1148),
    .Y(_09461_));
 sky130_fd_sc_hd__nand3_1 _29945_ (.A(_09437_),
    .B(net1159),
    .C(net1158),
    .Y(_09462_));
 sky130_fd_sc_hd__nor2_1 _29946_ (.A(_09461_),
    .B(_09462_),
    .Y(_09463_));
 sky130_fd_sc_hd__nand3b_1 _29947_ (.A_N(_09460_),
    .B(_09433_),
    .C(_09463_),
    .Y(_09464_));
 sky130_fd_sc_hd__nand2_1 _29949_ (.A(_09464_),
    .B(net1043),
    .Y(_09466_));
 sky130_fd_sc_hd__nor2_1 _29950_ (.A(net1272),
    .B(net1276),
    .Y(_09467_));
 sky130_fd_sc_hd__nand2_1 _29951_ (.A(_09467_),
    .B(net1674),
    .Y(_09468_));
 sky130_fd_sc_hd__o21ai_0 _29952_ (.A1(net1260),
    .A2(_09468_),
    .B1(net1042),
    .Y(_09469_));
 sky130_fd_sc_hd__nand2_1 _29953_ (.A(_09466_),
    .B(_09469_),
    .Y(_09470_));
 sky130_fd_sc_hd__nand2_1 _29954_ (.A(_09470_),
    .B(net1253),
    .Y(_09471_));
 sky130_fd_sc_hd__nand3_1 _29955_ (.A(_09466_),
    .B(net1670),
    .C(_09469_),
    .Y(_09472_));
 sky130_fd_sc_hd__nand2_1 _29956_ (.A(_09471_),
    .B(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__nand3_1 _29957_ (.A(net1366),
    .B(net1706),
    .C(net1691),
    .Y(_09474_));
 sky130_fd_sc_hd__nor2_1 _29958_ (.A(net1361),
    .B(net1356),
    .Y(_09475_));
 sky130_fd_sc_hd__nor2_1 _29959_ (.A(net1351),
    .B(net1350),
    .Y(_09476_));
 sky130_fd_sc_hd__nand2_1 _29960_ (.A(_09475_),
    .B(_09476_),
    .Y(_09477_));
 sky130_fd_sc_hd__nor2_1 _29961_ (.A(_09474_),
    .B(_09477_),
    .Y(_09478_));
 sky130_fd_sc_hd__nor2_1 _29962_ (.A(net1299),
    .B(net1295),
    .Y(_09479_));
 sky130_fd_sc_hd__nand3_1 _29963_ (.A(_09479_),
    .B(net1143),
    .C(net1142),
    .Y(_09480_));
 sky130_fd_sc_hd__nor2_1 _29964_ (.A(net1286),
    .B(net1289),
    .Y(_09481_));
 sky130_fd_sc_hd__nand3_1 _29965_ (.A(_09481_),
    .B(net1127),
    .C(net1678),
    .Y(_09482_));
 sky130_fd_sc_hd__nor2_1 _29966_ (.A(_09480_),
    .B(_09482_),
    .Y(_09483_));
 sky130_fd_sc_hd__nor2_1 _29967_ (.A(net1337),
    .B(net1331),
    .Y(_09484_));
 sky130_fd_sc_hd__nor2_1 _29968_ (.A(net1346),
    .B(net1341),
    .Y(_09485_));
 sky130_fd_sc_hd__nand2_1 _29969_ (.A(_09484_),
    .B(_09485_),
    .Y(_09486_));
 sky130_fd_sc_hd__nor2_1 _29970_ (.A(net1327),
    .B(net1322),
    .Y(_09487_));
 sky130_fd_sc_hd__nand3_1 _29971_ (.A(_09487_),
    .B(net1148),
    .C(net1145),
    .Y(_09488_));
 sky130_fd_sc_hd__nor2_1 _29972_ (.A(_09486_),
    .B(_09488_),
    .Y(_09489_));
 sky130_fd_sc_hd__nor2_1 _29973_ (.A(net1253),
    .B(_09468_),
    .Y(_09490_));
 sky130_fd_sc_hd__nand4_1 _29974_ (.A(_09478_),
    .B(_09483_),
    .C(_09489_),
    .D(_09490_),
    .Y(_09491_));
 sky130_fd_sc_hd__nand2_1 _29976_ (.A(_09491_),
    .B(net1042),
    .Y(_09493_));
 sky130_fd_sc_hd__nand2_1 _29977_ (.A(_09493_),
    .B(net1118),
    .Y(_09494_));
 sky130_fd_sc_hd__nand3_1 _29978_ (.A(_09491_),
    .B(net1453),
    .C(net1042),
    .Y(_09495_));
 sky130_fd_sc_hd__nand2_1 _29979_ (.A(_09494_),
    .B(_09495_),
    .Y(_09496_));
 sky130_fd_sc_hd__nand4_1 _29980_ (.A(_09478_),
    .B(_09483_),
    .C(_09467_),
    .D(_09489_),
    .Y(_09497_));
 sky130_fd_sc_hd__nand2_1 _29981_ (.A(_09497_),
    .B(net1042),
    .Y(_09498_));
 sky130_fd_sc_hd__nand2_1 _29982_ (.A(_09498_),
    .B(net1674),
    .Y(_09499_));
 sky130_fd_sc_hd__nand3_1 _29983_ (.A(_09497_),
    .B(net1256),
    .C(net1042),
    .Y(_09500_));
 sky130_fd_sc_hd__nand2_1 _29984_ (.A(_09499_),
    .B(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__nand4_1 _29985_ (.A(_09455_),
    .B(_09473_),
    .C(_09496_),
    .D(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__nor2_1 _29986_ (.A(net1453),
    .B(net1460),
    .Y(_09503_));
 sky130_fd_sc_hd__nand3_1 _29987_ (.A(_09503_),
    .B(net1114),
    .C(net1110),
    .Y(_09504_));
 sky130_fd_sc_hd__nor2_1 _29988_ (.A(_09504_),
    .B(_09491_),
    .Y(_09505_));
 sky130_fd_sc_hd__nor2_1 _29989_ (.A(_09449_),
    .B(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__nor2_1 _29990_ (.A(net1222),
    .B(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__nor2_1 _29991_ (.A(net1260),
    .B(_09468_),
    .Y(_09508_));
 sky130_fd_sc_hd__nand4_1 _29992_ (.A(_09508_),
    .B(net1114),
    .C(net1670),
    .D(_09503_),
    .Y(_09509_));
 sky130_fd_sc_hd__nor2_1 _29993_ (.A(_09460_),
    .B(_09509_),
    .Y(_09510_));
 sky130_fd_sc_hd__inv_1 _29994_ (.A(_09462_),
    .Y(_09511_));
 sky130_fd_sc_hd__nand2_1 _29995_ (.A(_09433_),
    .B(_09511_),
    .Y(_09512_));
 sky130_fd_sc_hd__nor2_1 _29996_ (.A(_09461_),
    .B(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__nand2_1 _29997_ (.A(_09510_),
    .B(_09513_),
    .Y(_09514_));
 sky130_fd_sc_hd__nand2_1 _29998_ (.A(_09514_),
    .B(net1043),
    .Y(_09515_));
 sky130_fd_sc_hd__nand2_1 _29999_ (.A(_09515_),
    .B(net1475),
    .Y(_09516_));
 sky130_fd_sc_hd__nand3_1 _30000_ (.A(_09514_),
    .B(net1110),
    .C(net1043),
    .Y(_09517_));
 sky130_fd_sc_hd__nand2_1 _30001_ (.A(_09516_),
    .B(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__nor2_1 _30002_ (.A(_09507_),
    .B(_09518_),
    .Y(_09519_));
 sky130_fd_sc_hd__nand3_1 _30003_ (.A(_09478_),
    .B(_09483_),
    .C(_09489_),
    .Y(_09520_));
 sky130_fd_sc_hd__nor3_1 _30004_ (.A(net1453),
    .B(net1253),
    .C(_09468_),
    .Y(_09521_));
 sky130_fd_sc_hd__nand3b_1 _30005_ (.A_N(_09520_),
    .B(net1735),
    .C(_09521_),
    .Y(_09522_));
 sky130_fd_sc_hd__nand2_1 _30006_ (.A(_09522_),
    .B(net1042),
    .Y(_09523_));
 sky130_fd_sc_hd__nand2_1 _30007_ (.A(_09523_),
    .B(net1468),
    .Y(_09524_));
 sky130_fd_sc_hd__nand3_1 _30008_ (.A(_09522_),
    .B(net1114),
    .C(net1042),
    .Y(_09525_));
 sky130_fd_sc_hd__nand2_1 _30009_ (.A(_09524_),
    .B(_09525_),
    .Y(_09526_));
 sky130_fd_sc_hd__inv_1 _30010_ (.A(_09526_),
    .Y(_09527_));
 sky130_fd_sc_hd__clkinv_1 _30011_ (.A(net1043),
    .Y(_09528_));
 sky130_fd_sc_hd__nand3_1 _30012_ (.A(_09521_),
    .B(net1678),
    .C(_09443_),
    .Y(_09529_));
 sky130_fd_sc_hd__nand3_1 _30013_ (.A(_09435_),
    .B(_09436_),
    .C(_09442_),
    .Y(_09530_));
 sky130_fd_sc_hd__nor2_1 _30014_ (.A(_09529_),
    .B(_09530_),
    .Y(_09531_));
 sky130_fd_sc_hd__o21ai_0 _30015_ (.A1(_09528_),
    .A2(_09531_),
    .B1(net1735),
    .Y(_09532_));
 sky130_fd_sc_hd__nor2_1 _30016_ (.A(_09528_),
    .B(_09531_),
    .Y(_09533_));
 sky130_fd_sc_hd__nand2_1 _30017_ (.A(_09533_),
    .B(net1460),
    .Y(_09534_));
 sky130_fd_sc_hd__nand2_1 _30018_ (.A(_09532_),
    .B(_09534_),
    .Y(_09535_));
 sky130_fd_sc_hd__nand3_1 _30019_ (.A(_09519_),
    .B(_09527_),
    .C(_09535_),
    .Y(_09536_));
 sky130_fd_sc_hd__nor2_1 _30020_ (.A(_09502_),
    .B(_09536_),
    .Y(_09537_));
 sky130_fd_sc_hd__inv_1 _30021_ (.A(_09474_),
    .Y(_09538_));
 sky130_fd_sc_hd__nand2_1 _30022_ (.A(_09538_),
    .B(_09475_),
    .Y(_09539_));
 sky130_fd_sc_hd__nand2_1 _30023_ (.A(_09539_),
    .B(net1041),
    .Y(_09540_));
 sky130_fd_sc_hd__xor2_1 _30024_ (.A(net1351),
    .B(_09540_),
    .X(_09541_));
 sky130_fd_sc_hd__nand2_1 _30025_ (.A(net1041),
    .B(_09432_),
    .Y(_09542_));
 sky130_fd_sc_hd__xor2_1 _30026_ (.A(net1356),
    .B(_09542_),
    .X(_09543_));
 sky130_fd_sc_hd__nand2_1 _30027_ (.A(_09541_),
    .B(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__nor2_1 _30028_ (.A(_09528_),
    .B(_09433_),
    .Y(_09545_));
 sky130_fd_sc_hd__xor2_1 _30029_ (.A(net1350),
    .B(_09545_),
    .X(_09546_));
 sky130_fd_sc_hd__nor2_1 _30030_ (.A(_09528_),
    .B(_09478_),
    .Y(_09547_));
 sky130_fd_sc_hd__xor2_1 _30031_ (.A(net1346),
    .B(_09547_),
    .X(_09548_));
 sky130_fd_sc_hd__nor2_1 _30032_ (.A(_09546_),
    .B(_09548_),
    .Y(_09549_));
 sky130_fd_sc_hd__inv_1 _30033_ (.A(_02844_),
    .Y(_09550_));
 sky130_fd_sc_hd__nand2_1 _30034_ (.A(net1041),
    .B(_09474_),
    .Y(_09551_));
 sky130_fd_sc_hd__xor2_1 _30035_ (.A(_05900_),
    .B(_09551_),
    .X(_09552_));
 sky130_fd_sc_hd__nor3_1 _30036_ (.A(_09550_),
    .B(net1153),
    .C(_09552_),
    .Y(_09553_));
 sky130_fd_sc_hd__nand3b_1 _30037_ (.A_N(_09544_),
    .B(_09549_),
    .C(_09553_),
    .Y(_09554_));
 sky130_fd_sc_hd__a21oi_1 _30038_ (.A1(_09478_),
    .A2(_09489_),
    .B1(_09528_),
    .Y(_09555_));
 sky130_fd_sc_hd__xor2_2 _30039_ (.A(net1308),
    .B(_09555_),
    .X(_09556_));
 sky130_fd_sc_hd__o21ai_0 _30040_ (.A1(_09528_),
    .A2(_09513_),
    .B1(net1312),
    .Y(_09557_));
 sky130_fd_sc_hd__nor2_1 _30041_ (.A(_09528_),
    .B(_09513_),
    .Y(_09558_));
 sky130_fd_sc_hd__nand2_1 _30042_ (.A(_09558_),
    .B(net1145),
    .Y(_09559_));
 sky130_fd_sc_hd__nand2_1 _30043_ (.A(_09557_),
    .B(_09559_),
    .Y(_09560_));
 sky130_fd_sc_hd__nor2_1 _30044_ (.A(_09556_),
    .B(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__nand4_1 _30045_ (.A(_09487_),
    .B(_09484_),
    .C(_09476_),
    .D(_09485_),
    .Y(_09562_));
 sky130_fd_sc_hd__nor2_1 _30046_ (.A(_09539_),
    .B(_09562_),
    .Y(_09563_));
 sky130_fd_sc_hd__nor2_1 _30047_ (.A(_09528_),
    .B(_09563_),
    .Y(_09564_));
 sky130_fd_sc_hd__xor2_1 _30048_ (.A(net1317),
    .B(_09564_),
    .X(_09565_));
 sky130_fd_sc_hd__nand3_1 _30049_ (.A(_09433_),
    .B(_09511_),
    .C(_09438_),
    .Y(_09566_));
 sky130_fd_sc_hd__nand2_1 _30050_ (.A(_09566_),
    .B(net1043),
    .Y(_09567_));
 sky130_fd_sc_hd__xor2_1 _30051_ (.A(net1150),
    .B(_09567_),
    .X(_09568_));
 sky130_fd_sc_hd__nor2_1 _30052_ (.A(_09565_),
    .B(_09568_),
    .Y(_09569_));
 sky130_fd_sc_hd__nand2_1 _30053_ (.A(_09561_),
    .B(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__nand2_1 _30054_ (.A(_09512_),
    .B(net1044),
    .Y(_09571_));
 sky130_fd_sc_hd__xor2_1 _30055_ (.A(net1156),
    .B(_09571_),
    .X(_09572_));
 sky130_fd_sc_hd__nor2_1 _30056_ (.A(_09486_),
    .B(_09477_),
    .Y(_09573_));
 sky130_fd_sc_hd__nand2_1 _30057_ (.A(_09573_),
    .B(_09538_),
    .Y(_09574_));
 sky130_fd_sc_hd__nand2_1 _30058_ (.A(_09574_),
    .B(net1041),
    .Y(_09575_));
 sky130_fd_sc_hd__xor2_1 _30059_ (.A(net1152),
    .B(_09575_),
    .X(_09576_));
 sky130_fd_sc_hd__nor2_1 _30060_ (.A(_09572_),
    .B(_09576_),
    .Y(_09577_));
 sky130_fd_sc_hd__nor2_1 _30061_ (.A(_09528_),
    .B(_09435_),
    .Y(_09578_));
 sky130_fd_sc_hd__xor2_1 _30062_ (.A(net1157),
    .B(_09578_),
    .X(_09579_));
 sky130_fd_sc_hd__nand2_1 _30063_ (.A(_09478_),
    .B(_09485_),
    .Y(_09580_));
 sky130_fd_sc_hd__nand2_1 _30064_ (.A(_09580_),
    .B(net1041),
    .Y(_09581_));
 sky130_fd_sc_hd__xor2_1 _30065_ (.A(_05907_),
    .B(_09581_),
    .X(_09582_));
 sky130_fd_sc_hd__inv_1 _30066_ (.A(_09582_),
    .Y(_09583_));
 sky130_fd_sc_hd__nand3_1 _30067_ (.A(_09577_),
    .B(_09579_),
    .C(_09583_),
    .Y(_09584_));
 sky130_fd_sc_hd__nor3_1 _30068_ (.A(_09554_),
    .B(_09570_),
    .C(_09584_),
    .Y(_09585_));
 sky130_fd_sc_hd__nand4_1 _30069_ (.A(net1148),
    .B(net1145),
    .C(net1143),
    .D(net1142),
    .Y(_09586_));
 sky130_fd_sc_hd__inv_1 _30070_ (.A(_09586_),
    .Y(_09587_));
 sky130_fd_sc_hd__nand4_1 _30071_ (.A(_09563_),
    .B(_09481_),
    .C(_09479_),
    .D(_09587_),
    .Y(_09588_));
 sky130_fd_sc_hd__nand2_1 _30072_ (.A(_09588_),
    .B(net1041),
    .Y(_09589_));
 sky130_fd_sc_hd__nand2_1 _30073_ (.A(_09589_),
    .B(net1127),
    .Y(_09590_));
 sky130_fd_sc_hd__nand3_1 _30074_ (.A(_09588_),
    .B(net1281),
    .C(net1042),
    .Y(_09591_));
 sky130_fd_sc_hd__nand2_1 _30075_ (.A(_09590_),
    .B(_09591_),
    .Y(_09592_));
 sky130_fd_sc_hd__nand2_1 _30076_ (.A(_09530_),
    .B(net1044),
    .Y(_09593_));
 sky130_fd_sc_hd__nand2_1 _30077_ (.A(_09593_),
    .B(net1130),
    .Y(_09594_));
 sky130_fd_sc_hd__nand3_1 _30078_ (.A(_09530_),
    .B(net1286),
    .C(net1044),
    .Y(_09595_));
 sky130_fd_sc_hd__nand2_1 _30079_ (.A(_09594_),
    .B(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__nand2_1 _30080_ (.A(_09592_),
    .B(_09596_),
    .Y(_09597_));
 sky130_fd_sc_hd__inv_1 _30081_ (.A(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__nand2_1 _30082_ (.A(_09520_),
    .B(net1044),
    .Y(_09599_));
 sky130_fd_sc_hd__xor2_1 _30083_ (.A(net1124),
    .B(_09599_),
    .X(_09600_));
 sky130_fd_sc_hd__xor2_1 _30084_ (.A(net1678),
    .B(_09466_),
    .X(_09601_));
 sky130_fd_sc_hd__nor2_1 _30085_ (.A(_09600_),
    .B(_09601_),
    .Y(_09602_));
 sky130_fd_sc_hd__nand2_1 _30086_ (.A(_09598_),
    .B(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__o21ai_0 _30087_ (.A1(_09441_),
    .A2(_09566_),
    .B1(net1043),
    .Y(_09604_));
 sky130_fd_sc_hd__xor2_2 _30088_ (.A(net1303),
    .B(_09604_),
    .X(_09605_));
 sky130_fd_sc_hd__nand2_1 _30089_ (.A(_09513_),
    .B(_09458_),
    .Y(_09606_));
 sky130_fd_sc_hd__nand2_1 _30090_ (.A(_09606_),
    .B(net1043),
    .Y(_09607_));
 sky130_fd_sc_hd__nand2_1 _30091_ (.A(_09607_),
    .B(net1137),
    .Y(_09608_));
 sky130_fd_sc_hd__nand3_1 _30092_ (.A(_09606_),
    .B(net1295),
    .C(net1043),
    .Y(_09609_));
 sky130_fd_sc_hd__nand2_1 _30093_ (.A(_09608_),
    .B(_09609_),
    .Y(_09610_));
 sky130_fd_sc_hd__nor2_1 _30094_ (.A(_09488_),
    .B(_09480_),
    .Y(_09611_));
 sky130_fd_sc_hd__nand3_1 _30095_ (.A(_09573_),
    .B(_09611_),
    .C(_09538_),
    .Y(_09612_));
 sky130_fd_sc_hd__nand2_1 _30096_ (.A(_09612_),
    .B(net1041),
    .Y(_09613_));
 sky130_fd_sc_hd__xor2_1 _30097_ (.A(net1289),
    .B(_09613_),
    .X(_09614_));
 sky130_fd_sc_hd__nand2_1 _30098_ (.A(_09563_),
    .B(_09587_),
    .Y(_09615_));
 sky130_fd_sc_hd__nand2_1 _30099_ (.A(_09615_),
    .B(net1041),
    .Y(_09616_));
 sky130_fd_sc_hd__nand2_1 _30100_ (.A(_09616_),
    .B(net1139),
    .Y(_09617_));
 sky130_fd_sc_hd__nand3_1 _30101_ (.A(_09615_),
    .B(net1299),
    .C(net1041),
    .Y(_09618_));
 sky130_fd_sc_hd__nand2_1 _30102_ (.A(_09617_),
    .B(_09618_),
    .Y(_09619_));
 sky130_fd_sc_hd__nand4_1 _30103_ (.A(_09605_),
    .B(_09610_),
    .C(_09614_),
    .D(_09619_),
    .Y(_09620_));
 sky130_fd_sc_hd__nor2_1 _30104_ (.A(_09603_),
    .B(_09620_),
    .Y(_09621_));
 sky130_fd_sc_hd__nand3_1 _30105_ (.A(_09537_),
    .B(_09585_),
    .C(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__nand2_1 _30106_ (.A(_03017_),
    .B(net1318),
    .Y(_09623_));
 sky130_fd_sc_hd__nor3_1 _30107_ (.A(net1424),
    .B(net1426),
    .C(_09623_),
    .Y(_09624_));
 sky130_fd_sc_hd__nand2_1 _30108_ (.A(net1722),
    .B(_02983_),
    .Y(_09625_));
 sky130_fd_sc_hd__nand2_1 _30109_ (.A(net1720),
    .B(net1716),
    .Y(_09626_));
 sky130_fd_sc_hd__nor2_1 _30110_ (.A(_09625_),
    .B(_09626_),
    .Y(_09627_));
 sky130_fd_sc_hd__nand2_1 _30111_ (.A(_09624_),
    .B(_09627_),
    .Y(_09628_));
 sky130_fd_sc_hd__nand2_1 _30112_ (.A(_20003_),
    .B(net1437),
    .Y(_09629_));
 sky130_fd_sc_hd__nor3_1 _30113_ (.A(net1447),
    .B(net1443),
    .C(_09629_),
    .Y(_09630_));
 sky130_fd_sc_hd__nor2_1 _30114_ (.A(net1734),
    .B(net1729),
    .Y(_09631_));
 sky130_fd_sc_hd__nor2_1 _30115_ (.A(net1725),
    .B(net1216),
    .Y(_09632_));
 sky130_fd_sc_hd__nand3_1 _30116_ (.A(_09630_),
    .B(_09631_),
    .C(_09632_),
    .Y(_09633_));
 sky130_fd_sc_hd__nor2_1 _30117_ (.A(_09628_),
    .B(_09633_),
    .Y(_09634_));
 sky130_fd_sc_hd__nor2_1 _30118_ (.A(net1394),
    .B(net1389),
    .Y(_09635_));
 sky130_fd_sc_hd__nand2_1 _30119_ (.A(_09635_),
    .B(_02700_),
    .Y(_09636_));
 sky130_fd_sc_hd__nand2_1 _30120_ (.A(_20061_),
    .B(_20734_),
    .Y(_09637_));
 sky130_fd_sc_hd__nand2_1 _30121_ (.A(_20067_),
    .B(net1399),
    .Y(_09638_));
 sky130_fd_sc_hd__nor2_1 _30122_ (.A(_09637_),
    .B(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__inv_1 _30123_ (.A(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__nor2_1 _30124_ (.A(net1398),
    .B(net1397),
    .Y(_09641_));
 sky130_fd_sc_hd__nand3_1 _30125_ (.A(_09641_),
    .B(net1170),
    .C(net1196),
    .Y(_09642_));
 sky130_fd_sc_hd__nor3_1 _30126_ (.A(_09636_),
    .B(_09640_),
    .C(_09642_),
    .Y(_09643_));
 sky130_fd_sc_hd__nand2_1 _30127_ (.A(_09634_),
    .B(_09643_),
    .Y(_09644_));
 sky130_fd_sc_hd__nand2_1 _30128_ (.A(_09644_),
    .B(net1217),
    .Y(_09645_));
 sky130_fd_sc_hd__nand3_1 _30129_ (.A(_09634_),
    .B(net1457),
    .C(_09643_),
    .Y(_09646_));
 sky130_fd_sc_hd__nand2_1 _30130_ (.A(_09645_),
    .B(_09646_),
    .Y(_09647_));
 sky130_fd_sc_hd__nor2_2 _30131_ (.A(_09449_),
    .B(net1739),
    .Y(_09648_));
 sky130_fd_sc_hd__nand2_1 _30134_ (.A(_09647_),
    .B(net1248),
    .Y(_09651_));
 sky130_fd_sc_hd__inv_1 _30135_ (.A(net1247),
    .Y(_09652_));
 sky130_fd_sc_hd__nand2_1 _30136_ (.A(_09652_),
    .B(net1457),
    .Y(_09653_));
 sky130_fd_sc_hd__nand2_1 _30137_ (.A(_09651_),
    .B(_09653_),
    .Y(_09654_));
 sky130_fd_sc_hd__nand3_4 _30138_ (.A(net1181),
    .B(net1697),
    .C(net1682),
    .Y(_09655_));
 sky130_fd_sc_hd__nor2_1 _30139_ (.A(net1203),
    .B(net1403),
    .Y(_09656_));
 sky130_fd_sc_hd__nor2_2 _30140_ (.A(net1398),
    .B(_03045_),
    .Y(_09657_));
 sky130_fd_sc_hd__nand2_1 _30141_ (.A(_09656_),
    .B(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__nor2_1 _30142_ (.A(net1397),
    .B(net1396),
    .Y(_09659_));
 sky130_fd_sc_hd__nand3_2 _30143_ (.A(_09659_),
    .B(net1196),
    .C(net1173),
    .Y(_09660_));
 sky130_fd_sc_hd__nor3_4 _30144_ (.A(_09655_),
    .B(_09658_),
    .C(_09660_),
    .Y(_09661_));
 sky130_fd_sc_hd__nand2_1 _30145_ (.A(net1716),
    .B(net1713),
    .Y(_09662_));
 sky130_fd_sc_hd__nand2_1 _30146_ (.A(net1720),
    .B(net1722),
    .Y(_09663_));
 sky130_fd_sc_hd__nor2_1 _30147_ (.A(_09662_),
    .B(_09663_),
    .Y(_09664_));
 sky130_fd_sc_hd__nand2_1 _30148_ (.A(net1318),
    .B(_20734_),
    .Y(_09665_));
 sky130_fd_sc_hd__nor3_1 _30149_ (.A(net1424),
    .B(net1420),
    .C(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__nand2_1 _30150_ (.A(_09664_),
    .B(_09666_),
    .Y(_09667_));
 sky130_fd_sc_hd__inv_1 _30151_ (.A(_09667_),
    .Y(_09668_));
 sky130_fd_sc_hd__nor2_1 _30152_ (.A(net1443),
    .B(net1210),
    .Y(_09669_));
 sky130_fd_sc_hd__nand3_1 _30153_ (.A(_09669_),
    .B(_20003_),
    .C(_02983_),
    .Y(_09670_));
 sky130_fd_sc_hd__nand4_1 _30154_ (.A(net1265),
    .B(net1268),
    .C(net1450),
    .D(net1213),
    .Y(_09671_));
 sky130_fd_sc_hd__nor2_1 _30155_ (.A(_09670_),
    .B(_09671_),
    .Y(_09672_));
 sky130_fd_sc_hd__nor2_1 _30156_ (.A(net1457),
    .B(net1734),
    .Y(_09673_));
 sky130_fd_sc_hd__nand4_1 _30157_ (.A(_09661_),
    .B(_09668_),
    .C(_09672_),
    .D(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__nand2_1 _30159_ (.A(_09674_),
    .B(net1246),
    .Y(_09676_));
 sky130_fd_sc_hd__nand2_1 _30160_ (.A(_09676_),
    .B(net1218),
    .Y(_09677_));
 sky130_fd_sc_hd__nand3_1 _30161_ (.A(_09674_),
    .B(net1465),
    .C(net1246),
    .Y(_09678_));
 sky130_fd_sc_hd__nand2_1 _30162_ (.A(_09677_),
    .B(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__inv_1 _30163_ (.A(_09679_),
    .Y(_09680_));
 sky130_fd_sc_hd__nor2_1 _30164_ (.A(_09654_),
    .B(_09680_),
    .Y(_09681_));
 sky130_fd_sc_hd__nor3_2 _30165_ (.A(_09670_),
    .B(_09671_),
    .C(_09667_),
    .Y(_09682_));
 sky130_fd_sc_hd__nor2_1 _30166_ (.A(net1473),
    .B(net1465),
    .Y(_09683_));
 sky130_fd_sc_hd__nand4_1 _30167_ (.A(_09682_),
    .B(_09661_),
    .C(_09673_),
    .D(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__a21oi_1 _30168_ (.A1(_09684_),
    .A2(_09448_),
    .B1(net1739),
    .Y(_09685_));
 sky130_fd_sc_hd__nor3_2 _30169_ (.A(net1426),
    .B(net1424),
    .C(_09626_),
    .Y(_09686_));
 sky130_fd_sc_hd__nor2_1 _30170_ (.A(_09629_),
    .B(_09625_),
    .Y(_09687_));
 sky130_fd_sc_hd__nand2_1 _30171_ (.A(_09686_),
    .B(_09687_),
    .Y(_09688_));
 sky130_fd_sc_hd__nand2_1 _30172_ (.A(net1213),
    .B(net1450),
    .Y(_09689_));
 sky130_fd_sc_hd__nor3_1 _30173_ (.A(net1725),
    .B(net1443),
    .C(_09689_),
    .Y(_09690_));
 sky130_fd_sc_hd__nor2_1 _30174_ (.A(net1457),
    .B(net1465),
    .Y(_09691_));
 sky130_fd_sc_hd__nand3_1 _30175_ (.A(_09690_),
    .B(_09631_),
    .C(_09691_),
    .Y(_09692_));
 sky130_fd_sc_hd__nor2_1 _30176_ (.A(_09688_),
    .B(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__nand4_2 _30177_ (.A(_09635_),
    .B(_02700_),
    .C(net1170),
    .D(net1196),
    .Y(_09694_));
 sky130_fd_sc_hd__nor2_1 _30178_ (.A(_09637_),
    .B(_09623_),
    .Y(_09695_));
 sky130_fd_sc_hd__inv_1 _30179_ (.A(_09638_),
    .Y(_09696_));
 sky130_fd_sc_hd__nand3_1 _30180_ (.A(_09695_),
    .B(_09696_),
    .C(_09641_),
    .Y(_09697_));
 sky130_fd_sc_hd__nor2_1 _30181_ (.A(_09694_),
    .B(_09697_),
    .Y(_09698_));
 sky130_fd_sc_hd__nand2_1 _30182_ (.A(_09693_),
    .B(_09698_),
    .Y(_09699_));
 sky130_fd_sc_hd__nand2_1 _30183_ (.A(_09699_),
    .B(net1219),
    .Y(_09700_));
 sky130_fd_sc_hd__nand3_1 _30184_ (.A(_09693_),
    .B(net1473),
    .C(_09698_),
    .Y(_09701_));
 sky130_fd_sc_hd__nand2_1 _30185_ (.A(_09700_),
    .B(_09701_),
    .Y(_09702_));
 sky130_fd_sc_hd__nand2_1 _30186_ (.A(_09702_),
    .B(net1247),
    .Y(_09703_));
 sky130_fd_sc_hd__nand2_1 _30187_ (.A(_09652_),
    .B(net1473),
    .Y(_09704_));
 sky130_fd_sc_hd__nand2_1 _30188_ (.A(_09703_),
    .B(_09704_),
    .Y(_09705_));
 sky130_fd_sc_hd__nor2_1 _30189_ (.A(_09685_),
    .B(_09705_),
    .Y(_09706_));
 sky130_fd_sc_hd__nand2_1 _30190_ (.A(_09681_),
    .B(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__and2_1 _30191_ (.A(_09630_),
    .B(_09627_),
    .X(_09708_));
 sky130_fd_sc_hd__inv_1 _30192_ (.A(_09624_),
    .Y(_09709_));
 sky130_fd_sc_hd__nor2_1 _30193_ (.A(_09640_),
    .B(_09709_),
    .Y(_09710_));
 sky130_fd_sc_hd__inv_1 _30194_ (.A(_09641_),
    .Y(_09711_));
 sky130_fd_sc_hd__nor2_2 _30195_ (.A(_09711_),
    .B(_09694_),
    .Y(_09712_));
 sky130_fd_sc_hd__nand3_1 _30196_ (.A(_09708_),
    .B(_09710_),
    .C(_09712_),
    .Y(_09713_));
 sky130_fd_sc_hd__nand2_1 _30197_ (.A(_09713_),
    .B(net1450),
    .Y(_09714_));
 sky130_fd_sc_hd__nand4_1 _30198_ (.A(_09708_),
    .B(_09710_),
    .C(net1216),
    .D(_09712_),
    .Y(_09715_));
 sky130_fd_sc_hd__nand2_1 _30199_ (.A(_09714_),
    .B(_09715_),
    .Y(_09716_));
 sky130_fd_sc_hd__nand2_1 _30200_ (.A(_09716_),
    .B(net1248),
    .Y(_09717_));
 sky130_fd_sc_hd__nand2_1 _30201_ (.A(_09652_),
    .B(net1216),
    .Y(_09718_));
 sky130_fd_sc_hd__nand2_1 _30202_ (.A(_09717_),
    .B(_09718_),
    .Y(_09719_));
 sky130_fd_sc_hd__nor2_2 _30203_ (.A(_09655_),
    .B(_09660_),
    .Y(_09720_));
 sky130_fd_sc_hd__inv_1 _30204_ (.A(_09665_),
    .Y(_09721_));
 sky130_fd_sc_hd__nand3_1 _30205_ (.A(_09721_),
    .B(_03011_),
    .C(_03017_),
    .Y(_09722_));
 sky130_fd_sc_hd__nor2_1 _30206_ (.A(_09658_),
    .B(_09722_),
    .Y(_09723_));
 sky130_fd_sc_hd__nand2_1 _30207_ (.A(_09720_),
    .B(_09723_),
    .Y(_09724_));
 sky130_fd_sc_hd__nor2_2 _30208_ (.A(_09662_),
    .B(_09724_),
    .Y(_09725_));
 sky130_fd_sc_hd__nor3_1 _30209_ (.A(_09663_),
    .B(_09689_),
    .C(_09670_),
    .Y(_09726_));
 sky130_fd_sc_hd__a21oi_1 _30210_ (.A1(_09725_),
    .A2(_09726_),
    .B1(_09652_),
    .Y(_09727_));
 sky130_fd_sc_hd__xor2_1 _30211_ (.A(net1725),
    .B(_09727_),
    .X(_09728_));
 sky130_fd_sc_hd__nor2_1 _30212_ (.A(_09719_),
    .B(_09728_),
    .Y(_09729_));
 sky130_fd_sc_hd__nand2_1 _30213_ (.A(_09682_),
    .B(_09661_),
    .Y(_09730_));
 sky130_fd_sc_hd__nand2_1 _30214_ (.A(_09730_),
    .B(net1246),
    .Y(_09731_));
 sky130_fd_sc_hd__xor2_1 _30215_ (.A(net1264),
    .B(_09731_),
    .X(_09732_));
 sky130_fd_sc_hd__nor2_1 _30216_ (.A(_09652_),
    .B(_09690_),
    .Y(_09733_));
 sky130_fd_sc_hd__nand2_1 _30217_ (.A(_09712_),
    .B(_09696_),
    .Y(_09734_));
 sky130_fd_sc_hd__nand2_1 _30218_ (.A(_09734_),
    .B(net1248),
    .Y(_09735_));
 sky130_fd_sc_hd__nand2_1 _30219_ (.A(_09686_),
    .B(_09695_),
    .Y(_09736_));
 sky130_fd_sc_hd__nand2_1 _30220_ (.A(_09736_),
    .B(net1249),
    .Y(_09737_));
 sky130_fd_sc_hd__o21ai_0 _30221_ (.A1(_09629_),
    .A2(_09625_),
    .B1(net1249),
    .Y(_09738_));
 sky130_fd_sc_hd__nand3_1 _30222_ (.A(_09735_),
    .B(_09737_),
    .C(_09738_),
    .Y(_09739_));
 sky130_fd_sc_hd__o21ai_1 _30223_ (.A1(_09733_),
    .A2(_09739_),
    .B1(net1265),
    .Y(_09740_));
 sky130_fd_sc_hd__nand2_1 _30224_ (.A(_09735_),
    .B(_09737_),
    .Y(_09741_));
 sky130_fd_sc_hd__clkinv_1 _30225_ (.A(_09741_),
    .Y(_09742_));
 sky130_fd_sc_hd__or2_2 _30226_ (.A(_09652_),
    .B(_09690_),
    .X(_09743_));
 sky130_fd_sc_hd__nand4_1 _30227_ (.A(_09742_),
    .B(net1729),
    .C(_09738_),
    .D(_09743_),
    .Y(_09744_));
 sky130_fd_sc_hd__nand2_1 _30228_ (.A(_09740_),
    .B(_09744_),
    .Y(_09745_));
 sky130_fd_sc_hd__nor2_1 _30229_ (.A(_09732_),
    .B(_09745_),
    .Y(_09746_));
 sky130_fd_sc_hd__nand2_1 _30230_ (.A(_09729_),
    .B(_09746_),
    .Y(_09747_));
 sky130_fd_sc_hd__nor2_2 _30231_ (.A(_09707_),
    .B(_09747_),
    .Y(_09748_));
 sky130_fd_sc_hd__nand2_1 _30232_ (.A(_09636_),
    .B(net1248),
    .Y(_09749_));
 sky130_fd_sc_hd__xor2_1 _30233_ (.A(net1196),
    .B(_09749_),
    .X(_09750_));
 sky130_fd_sc_hd__nor2_1 _30234_ (.A(net1394),
    .B(_09655_),
    .Y(_09751_));
 sky130_fd_sc_hd__a21oi_1 _30235_ (.A1(_09751_),
    .A2(net1196),
    .B1(_09652_),
    .Y(_09752_));
 sky130_fd_sc_hd__xor2_1 _30236_ (.A(net1170),
    .B(_09752_),
    .X(_09753_));
 sky130_fd_sc_hd__inv_1 _30237_ (.A(_09753_),
    .Y(_09754_));
 sky130_fd_sc_hd__nor2_1 _30238_ (.A(_09750_),
    .B(_09754_),
    .Y(_09755_));
 sky130_fd_sc_hd__nand2_1 _30239_ (.A(_09694_),
    .B(net1248),
    .Y(_09756_));
 sky130_fd_sc_hd__xor2_1 _30240_ (.A(net1397),
    .B(_09756_),
    .X(_09757_));
 sky130_fd_sc_hd__inv_1 _30241_ (.A(_02700_),
    .Y(_09758_));
 sky130_fd_sc_hd__nand2_1 _30242_ (.A(_09655_),
    .B(net1248),
    .Y(_09759_));
 sky130_fd_sc_hd__xor2_1 _30243_ (.A(net1394),
    .B(_09759_),
    .X(_09760_));
 sky130_fd_sc_hd__inv_1 _30244_ (.A(_09760_),
    .Y(_09761_));
 sky130_fd_sc_hd__nor3_1 _30245_ (.A(_09758_),
    .B(net1389),
    .C(_09761_),
    .Y(_09762_));
 sky130_fd_sc_hd__o21ai_0 _30246_ (.A1(_09655_),
    .A2(_09660_),
    .B1(net1247),
    .Y(_09763_));
 sky130_fd_sc_hd__xor2_1 _30247_ (.A(net1398),
    .B(_09763_),
    .X(_09764_));
 sky130_fd_sc_hd__nand4_1 _30248_ (.A(_09755_),
    .B(_09757_),
    .C(_09762_),
    .D(_09764_),
    .Y(_09765_));
 sky130_fd_sc_hd__o21ai_0 _30249_ (.A1(_09652_),
    .A2(_09661_),
    .B1(net1411),
    .Y(_09766_));
 sky130_fd_sc_hd__inv_1 _30250_ (.A(_09661_),
    .Y(_09767_));
 sky130_fd_sc_hd__nand3_1 _30251_ (.A(_09767_),
    .B(_20734_),
    .C(net1247),
    .Y(_09768_));
 sky130_fd_sc_hd__nand2_1 _30252_ (.A(_09766_),
    .B(_09768_),
    .Y(_09769_));
 sky130_fd_sc_hd__nand2_1 _30253_ (.A(_09735_),
    .B(_20061_),
    .Y(_09770_));
 sky130_fd_sc_hd__nand3_1 _30254_ (.A(_09734_),
    .B(net1203),
    .C(net1249),
    .Y(_09771_));
 sky130_fd_sc_hd__nand2_1 _30255_ (.A(_09770_),
    .B(_09771_),
    .Y(_09772_));
 sky130_fd_sc_hd__inv_1 _30256_ (.A(_09772_),
    .Y(_09773_));
 sky130_fd_sc_hd__nand2_1 _30257_ (.A(_09720_),
    .B(_09657_),
    .Y(_09774_));
 sky130_fd_sc_hd__nand2_1 _30258_ (.A(_09774_),
    .B(net1247),
    .Y(_09775_));
 sky130_fd_sc_hd__xor2_1 _30259_ (.A(net1403),
    .B(_09775_),
    .X(_09776_));
 sky130_fd_sc_hd__o21ai_0 _30260_ (.A1(_09711_),
    .A2(_09694_),
    .B1(net1248),
    .Y(_09777_));
 sky130_fd_sc_hd__xor2_1 _30261_ (.A(_03045_),
    .B(_09777_),
    .X(_09778_));
 sky130_fd_sc_hd__nand2_1 _30262_ (.A(_09776_),
    .B(_09778_),
    .Y(_09779_));
 sky130_fd_sc_hd__nor3_1 _30263_ (.A(_09769_),
    .B(_09773_),
    .C(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__nor3_1 _30264_ (.A(net1203),
    .B(net1403),
    .C(_09665_),
    .Y(_09781_));
 sky130_fd_sc_hd__nand3_1 _30265_ (.A(_09720_),
    .B(_09657_),
    .C(_09781_),
    .Y(_09782_));
 sky130_fd_sc_hd__nand2_1 _30266_ (.A(_09782_),
    .B(net1246),
    .Y(_09783_));
 sky130_fd_sc_hd__xor2_1 _30267_ (.A(net1420),
    .B(_09783_),
    .X(_09784_));
 sky130_fd_sc_hd__nand2_1 _30268_ (.A(_09712_),
    .B(_09639_),
    .Y(_09785_));
 sky130_fd_sc_hd__nand2_1 _30269_ (.A(_09785_),
    .B(net1249),
    .Y(_09786_));
 sky130_fd_sc_hd__xor2_1 _30270_ (.A(net1415),
    .B(_09786_),
    .X(_09787_));
 sky130_fd_sc_hd__nand2_1 _30271_ (.A(_09784_),
    .B(_09787_),
    .Y(_09788_));
 sky130_fd_sc_hd__nand2_1 _30272_ (.A(_09724_),
    .B(net1246),
    .Y(_09789_));
 sky130_fd_sc_hd__xor2_1 _30273_ (.A(net1713),
    .B(_09789_),
    .X(_09790_));
 sky130_fd_sc_hd__inv_1 _30274_ (.A(_09790_),
    .Y(_09791_));
 sky130_fd_sc_hd__nand3_1 _30275_ (.A(_09712_),
    .B(_09696_),
    .C(_09695_),
    .Y(_09792_));
 sky130_fd_sc_hd__nand2_1 _30276_ (.A(_09792_),
    .B(net1246),
    .Y(_09793_));
 sky130_fd_sc_hd__nand2_1 _30277_ (.A(_09793_),
    .B(_03011_),
    .Y(_09794_));
 sky130_fd_sc_hd__nand3_1 _30278_ (.A(_09792_),
    .B(net1424),
    .C(net1246),
    .Y(_09795_));
 sky130_fd_sc_hd__nand2_1 _30279_ (.A(_09794_),
    .B(_09795_),
    .Y(_09796_));
 sky130_fd_sc_hd__nand2_1 _30280_ (.A(_09791_),
    .B(_09796_),
    .Y(_09797_));
 sky130_fd_sc_hd__nor2_1 _30281_ (.A(_09788_),
    .B(_09797_),
    .Y(_09798_));
 sky130_fd_sc_hd__nand2_1 _30282_ (.A(_09780_),
    .B(_09798_),
    .Y(_09799_));
 sky130_fd_sc_hd__nor2_2 _30283_ (.A(_09765_),
    .B(_09799_),
    .Y(_09800_));
 sky130_fd_sc_hd__xor2_1 _30284_ (.A(_20014_),
    .B(_09741_),
    .X(_09801_));
 sky130_fd_sc_hd__nand2_1 _30285_ (.A(_09661_),
    .B(_09668_),
    .Y(_09802_));
 sky130_fd_sc_hd__nand2_1 _30286_ (.A(_09802_),
    .B(net1246),
    .Y(_09803_));
 sky130_fd_sc_hd__xor2_1 _30287_ (.A(net1435),
    .B(_09803_),
    .X(_09804_));
 sky130_fd_sc_hd__inv_1 _30288_ (.A(_09804_),
    .Y(_09805_));
 sky130_fd_sc_hd__nor2_1 _30289_ (.A(_09801_),
    .B(_09805_),
    .Y(_09806_));
 sky130_fd_sc_hd__o21ai_1 _30290_ (.A1(_09662_),
    .A2(_09724_),
    .B1(net1246),
    .Y(_09807_));
 sky130_fd_sc_hd__xor2_1 _30291_ (.A(net1720),
    .B(_09807_),
    .X(_09808_));
 sky130_fd_sc_hd__nand2_1 _30292_ (.A(_09709_),
    .B(net1249),
    .Y(_09809_));
 sky130_fd_sc_hd__nand2_1 _30293_ (.A(_09786_),
    .B(_09809_),
    .Y(_09810_));
 sky130_fd_sc_hd__xor2_1 _30294_ (.A(_20024_),
    .B(_09810_),
    .X(_09811_));
 sky130_fd_sc_hd__nor2_1 _30295_ (.A(_09808_),
    .B(_09811_),
    .Y(_09812_));
 sky130_fd_sc_hd__nand2_1 _30296_ (.A(_09806_),
    .B(_09812_),
    .Y(_09813_));
 sky130_fd_sc_hd__nor3_1 _30297_ (.A(net1135),
    .B(net1435),
    .C(_09663_),
    .Y(_09814_));
 sky130_fd_sc_hd__nand3_1 _30298_ (.A(_09725_),
    .B(_09814_),
    .C(_09669_),
    .Y(_09815_));
 sky130_fd_sc_hd__nand2_1 _30299_ (.A(_09815_),
    .B(net1247),
    .Y(_09816_));
 sky130_fd_sc_hd__nand2_1 _30300_ (.A(_09816_),
    .B(net1213),
    .Y(_09817_));
 sky130_fd_sc_hd__nand3_1 _30301_ (.A(_09815_),
    .B(net1447),
    .C(net1246),
    .Y(_09818_));
 sky130_fd_sc_hd__nand2_1 _30302_ (.A(_09817_),
    .B(_09818_),
    .Y(_09819_));
 sky130_fd_sc_hd__nand3_1 _30303_ (.A(_09742_),
    .B(net1211),
    .C(_09738_),
    .Y(_09820_));
 sky130_fd_sc_hd__nand2_1 _30304_ (.A(_09739_),
    .B(net1443),
    .Y(_09821_));
 sky130_fd_sc_hd__nand2_1 _30305_ (.A(_09820_),
    .B(_09821_),
    .Y(_09822_));
 sky130_fd_sc_hd__nand2_1 _30306_ (.A(_09819_),
    .B(_09822_),
    .Y(_09823_));
 sky130_fd_sc_hd__inv_1 _30307_ (.A(_09823_),
    .Y(_09824_));
 sky130_fd_sc_hd__nand2_1 _30308_ (.A(_09725_),
    .B(_09814_),
    .Y(_09825_));
 sky130_fd_sc_hd__nand2_1 _30309_ (.A(_09825_),
    .B(net1249),
    .Y(_09826_));
 sky130_fd_sc_hd__nand2_1 _30310_ (.A(_09826_),
    .B(net1210),
    .Y(_09827_));
 sky130_fd_sc_hd__nand3_1 _30311_ (.A(_09825_),
    .B(net1437),
    .C(net1249),
    .Y(_09828_));
 sky130_fd_sc_hd__nand2_1 _30312_ (.A(_09827_),
    .B(_09828_),
    .Y(_09829_));
 sky130_fd_sc_hd__o21ai_0 _30313_ (.A1(_09625_),
    .A2(_09626_),
    .B1(net1249),
    .Y(_09830_));
 sky130_fd_sc_hd__nand3_1 _30314_ (.A(_09786_),
    .B(_09809_),
    .C(_09830_),
    .Y(_09831_));
 sky130_fd_sc_hd__xor2_1 _30315_ (.A(net1135),
    .B(_09831_),
    .X(_09832_));
 sky130_fd_sc_hd__nor2_1 _30316_ (.A(_09829_),
    .B(_09832_),
    .Y(_09833_));
 sky130_fd_sc_hd__nand2_1 _30317_ (.A(_09824_),
    .B(_09833_),
    .Y(_09834_));
 sky130_fd_sc_hd__nor2_2 _30318_ (.A(_09813_),
    .B(_09834_),
    .Y(_09835_));
 sky130_fd_sc_hd__nand3_1 _30319_ (.A(_09748_),
    .B(_09800_),
    .C(_09835_),
    .Y(_09836_));
 sky130_fd_sc_hd__nor2_1 _30320_ (.A(net1903),
    .B(_20231_),
    .Y(_09837_));
 sky130_fd_sc_hd__nand2_1 _30322_ (.A(_09837_),
    .B(net2842),
    .Y(_09839_));
 sky130_fd_sc_hd__inv_1 _30323_ (.A(_09839_),
    .Y(_09840_));
 sky130_fd_sc_hd__nand3_2 _30324_ (.A(_09622_),
    .B(_09836_),
    .C(_09840_),
    .Y(_09841_));
 sky130_fd_sc_hd__inv_2 _30326_ (.A(net615),
    .Y(_09843_));
 sky130_fd_sc_hd__nor2_1 _30327_ (.A(\inst$top.soc.cpu.divider.divisor[0] ),
    .B(_09843_),
    .Y(_09844_));
 sky130_fd_sc_hd__o21ai_1 _30331_ (.A1(net1251),
    .A2(net615),
    .B1(net2116),
    .Y(_09848_));
 sky130_fd_sc_hd__nor2_4 _30332_ (.A(_09844_),
    .B(_09848_),
    .Y(_03677_));
 sky130_fd_sc_hd__o21ai_1 _30334_ (.A1(_09773_),
    .A2(net615),
    .B1(net2116),
    .Y(_09850_));
 sky130_fd_sc_hd__a21oi_4 _30335_ (.A1(_02814_),
    .A2(net614),
    .B1(_09850_),
    .Y(_03678_));
 sky130_fd_sc_hd__o21ai_1 _30336_ (.A1(_09769_),
    .A2(net619),
    .B1(net2117),
    .Y(_09851_));
 sky130_fd_sc_hd__a21oi_4 _30337_ (.A1(_02811_),
    .A2(net619),
    .B1(_09851_),
    .Y(_03679_));
 sky130_fd_sc_hd__inv_1 _30338_ (.A(_09787_),
    .Y(_09852_));
 sky130_fd_sc_hd__o21ai_1 _30340_ (.A1(_09852_),
    .A2(net614),
    .B1(net2117),
    .Y(_09854_));
 sky130_fd_sc_hd__a21oi_4 _30341_ (.A1(_02808_),
    .A2(net613),
    .B1(_09854_),
    .Y(_03680_));
 sky130_fd_sc_hd__inv_1 _30342_ (.A(_09784_),
    .Y(_09855_));
 sky130_fd_sc_hd__o21ai_1 _30343_ (.A1(_09855_),
    .A2(net614),
    .B1(net2103),
    .Y(_09856_));
 sky130_fd_sc_hd__a21oi_4 _30344_ (.A1(_02805_),
    .A2(net613),
    .B1(_09856_),
    .Y(_03681_));
 sky130_fd_sc_hd__inv_1 _30345_ (.A(_09796_),
    .Y(_09857_));
 sky130_fd_sc_hd__o21ai_1 _30346_ (.A1(_09857_),
    .A2(net614),
    .B1(net2103),
    .Y(_09858_));
 sky130_fd_sc_hd__a21oi_4 _30347_ (.A1(_02802_),
    .A2(net613),
    .B1(_09858_),
    .Y(_03682_));
 sky130_fd_sc_hd__o21ai_1 _30348_ (.A1(_09790_),
    .A2(net615),
    .B1(net2116),
    .Y(_09859_));
 sky130_fd_sc_hd__a21oi_4 _30349_ (.A1(_02799_),
    .A2(net615),
    .B1(_09859_),
    .Y(_03683_));
 sky130_fd_sc_hd__o21ai_1 _30350_ (.A1(_09811_),
    .A2(net617),
    .B1(net2115),
    .Y(_09860_));
 sky130_fd_sc_hd__a21oi_4 _30351_ (.A1(_02796_),
    .A2(net614),
    .B1(_09860_),
    .Y(_03684_));
 sky130_fd_sc_hd__o21ai_1 _30353_ (.A1(_09808_),
    .A2(net617),
    .B1(net2115),
    .Y(_09862_));
 sky130_fd_sc_hd__a21oi_4 _30354_ (.A1(_02793_),
    .A2(net613),
    .B1(_09862_),
    .Y(_03685_));
 sky130_fd_sc_hd__o21ai_1 _30355_ (.A1(_09801_),
    .A2(net613),
    .B1(net2103),
    .Y(_09863_));
 sky130_fd_sc_hd__a21oi_4 _30356_ (.A1(_02790_),
    .A2(net613),
    .B1(_09863_),
    .Y(_03686_));
 sky130_fd_sc_hd__o21ai_1 _30357_ (.A1(_09805_),
    .A2(net613),
    .B1(net2103),
    .Y(_09864_));
 sky130_fd_sc_hd__a21oi_4 _30358_ (.A1(_02787_),
    .A2(net613),
    .B1(_09864_),
    .Y(_03687_));
 sky130_fd_sc_hd__nand2_1 _30359_ (.A(net1248),
    .B(_02701_),
    .Y(_09865_));
 sky130_fd_sc_hd__o21ai_0 _30360_ (.A1(net1697),
    .A2(net1248),
    .B1(_09865_),
    .Y(_09866_));
 sky130_fd_sc_hd__nand2_1 _30361_ (.A(_09843_),
    .B(_09866_),
    .Y(_09867_));
 sky130_fd_sc_hd__nand2_1 _30362_ (.A(net615),
    .B(\inst$top.soc.cpu.divider.divisor[1] ),
    .Y(_09868_));
 sky130_fd_sc_hd__a21oi_4 _30363_ (.A1(_09867_),
    .A2(_09868_),
    .B1(net2977),
    .Y(_03688_));
 sky130_fd_sc_hd__o21ai_1 _30365_ (.A1(_09832_),
    .A2(net616),
    .B1(net2115),
    .Y(_09870_));
 sky130_fd_sc_hd__a21oi_4 _30366_ (.A1(_02784_),
    .A2(net614),
    .B1(_09870_),
    .Y(_03689_));
 sky130_fd_sc_hd__o21ai_1 _30367_ (.A1(_09829_),
    .A2(net616),
    .B1(net2115),
    .Y(_09871_));
 sky130_fd_sc_hd__a21oi_4 _30368_ (.A1(_02781_),
    .A2(net614),
    .B1(_09871_),
    .Y(_03690_));
 sky130_fd_sc_hd__inv_1 _30369_ (.A(_09822_),
    .Y(_09872_));
 sky130_fd_sc_hd__o21ai_1 _30371_ (.A1(_09872_),
    .A2(net616),
    .B1(net2115),
    .Y(_09874_));
 sky130_fd_sc_hd__a21oi_4 _30372_ (.A1(_02778_),
    .A2(net619),
    .B1(_09874_),
    .Y(_03691_));
 sky130_fd_sc_hd__inv_1 _30373_ (.A(_09819_),
    .Y(_09875_));
 sky130_fd_sc_hd__o21ai_1 _30374_ (.A1(_09875_),
    .A2(net617),
    .B1(net2115),
    .Y(_09876_));
 sky130_fd_sc_hd__a21oi_4 _30375_ (.A1(_02775_),
    .A2(net616),
    .B1(_09876_),
    .Y(_03692_));
 sky130_fd_sc_hd__o21ai_1 _30376_ (.A1(_09719_),
    .A2(net617),
    .B1(net2116),
    .Y(_09877_));
 sky130_fd_sc_hd__a21oi_4 _30377_ (.A1(_02772_),
    .A2(net617),
    .B1(_09877_),
    .Y(_03693_));
 sky130_fd_sc_hd__o21ai_1 _30378_ (.A1(_09728_),
    .A2(net617),
    .B1(net2116),
    .Y(_09878_));
 sky130_fd_sc_hd__a21oi_4 _30379_ (.A1(_02769_),
    .A2(net617),
    .B1(_09878_),
    .Y(_03694_));
 sky130_fd_sc_hd__o21ai_1 _30380_ (.A1(_09745_),
    .A2(net616),
    .B1(net2115),
    .Y(_09879_));
 sky130_fd_sc_hd__a21oi_4 _30381_ (.A1(_02766_),
    .A2(net619),
    .B1(_09879_),
    .Y(_03695_));
 sky130_fd_sc_hd__o21ai_1 _30384_ (.A1(_09732_),
    .A2(net616),
    .B1(net2116),
    .Y(_09882_));
 sky130_fd_sc_hd__a21oi_4 _30385_ (.A1(_02763_),
    .A2(net619),
    .B1(_09882_),
    .Y(_03696_));
 sky130_fd_sc_hd__o21ai_1 _30386_ (.A1(_09654_),
    .A2(net616),
    .B1(net2115),
    .Y(_09883_));
 sky130_fd_sc_hd__a21oi_4 _30387_ (.A1(_02760_),
    .A2(net616),
    .B1(_09883_),
    .Y(_03697_));
 sky130_fd_sc_hd__o21ai_1 _30388_ (.A1(_09680_),
    .A2(net616),
    .B1(net2115),
    .Y(_09884_));
 sky130_fd_sc_hd__a21oi_4 _30389_ (.A1(_02757_),
    .A2(net616),
    .B1(_09884_),
    .Y(_03698_));
 sky130_fd_sc_hd__nand2_1 _30391_ (.A(net1248),
    .B(_09758_),
    .Y(_09886_));
 sky130_fd_sc_hd__xor2_1 _30392_ (.A(net1181),
    .B(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__o21ai_1 _30393_ (.A1(_09887_),
    .A2(net618),
    .B1(net2116),
    .Y(_09888_));
 sky130_fd_sc_hd__a21oi_4 _30394_ (.A1(_02838_),
    .A2(net618),
    .B1(_09888_),
    .Y(_03699_));
 sky130_fd_sc_hd__o21ai_1 _30395_ (.A1(_09705_),
    .A2(net617),
    .B1(net2115),
    .Y(_09889_));
 sky130_fd_sc_hd__a21oi_4 _30396_ (.A1(_02754_),
    .A2(net617),
    .B1(_09889_),
    .Y(_03700_));
 sky130_fd_sc_hd__nand2_1 _30397_ (.A(_09843_),
    .B(_09685_),
    .Y(_09890_));
 sky130_fd_sc_hd__nand2_1 _30398_ (.A(net618),
    .B(\inst$top.soc.cpu.divider.divisor[31] ),
    .Y(_09891_));
 sky130_fd_sc_hd__a21oi_4 _30399_ (.A1(_09890_),
    .A2(_09891_),
    .B1(net2977),
    .Y(_03701_));
 sky130_fd_sc_hd__o21ai_1 _30400_ (.A1(_09761_),
    .A2(net611),
    .B1(net2103),
    .Y(_09892_));
 sky130_fd_sc_hd__a21oi_4 _30401_ (.A1(_02835_),
    .A2(net612),
    .B1(_09892_),
    .Y(_03702_));
 sky130_fd_sc_hd__o21ai_1 _30402_ (.A1(_09750_),
    .A2(net615),
    .B1(net2116),
    .Y(_09893_));
 sky130_fd_sc_hd__a21oi_4 _30403_ (.A1(_02832_),
    .A2(net615),
    .B1(_09893_),
    .Y(_03703_));
 sky130_fd_sc_hd__o21ai_1 _30404_ (.A1(_09754_),
    .A2(net615),
    .B1(net2116),
    .Y(_09894_));
 sky130_fd_sc_hd__a21oi_4 _30405_ (.A1(_02829_),
    .A2(net615),
    .B1(_09894_),
    .Y(_03704_));
 sky130_fd_sc_hd__inv_1 _30406_ (.A(_09757_),
    .Y(_09895_));
 sky130_fd_sc_hd__o21ai_1 _30407_ (.A1(_09895_),
    .A2(net614),
    .B1(net2117),
    .Y(_09896_));
 sky130_fd_sc_hd__a21oi_4 _30408_ (.A1(_02826_),
    .A2(net614),
    .B1(_09896_),
    .Y(_03705_));
 sky130_fd_sc_hd__inv_1 _30409_ (.A(_09764_),
    .Y(_09897_));
 sky130_fd_sc_hd__o21ai_1 _30410_ (.A1(_09897_),
    .A2(net611),
    .B1(net2103),
    .Y(_09898_));
 sky130_fd_sc_hd__a21oi_4 _30411_ (.A1(_02823_),
    .A2(net612),
    .B1(_09898_),
    .Y(_03706_));
 sky130_fd_sc_hd__inv_1 _30412_ (.A(_09778_),
    .Y(_09899_));
 sky130_fd_sc_hd__o21ai_1 _30414_ (.A1(_09899_),
    .A2(net612),
    .B1(net2118),
    .Y(_09901_));
 sky130_fd_sc_hd__a21oi_4 _30415_ (.A1(_02820_),
    .A2(net612),
    .B1(_09901_),
    .Y(_03707_));
 sky130_fd_sc_hd__inv_1 _30416_ (.A(_09776_),
    .Y(_09902_));
 sky130_fd_sc_hd__o21ai_1 _30417_ (.A1(_09902_),
    .A2(net611),
    .B1(net2103),
    .Y(_09903_));
 sky130_fd_sc_hd__a21oi_4 _30418_ (.A1(_02817_),
    .A2(net612),
    .B1(_09903_),
    .Y(_03708_));
 sky130_fd_sc_hd__nor2_1 _30419_ (.A(\inst$top.soc.cpu.divider.timer[2] ),
    .B(\inst$top.soc.cpu.divider.timer[3] ),
    .Y(_09904_));
 sky130_fd_sc_hd__nand2_1 _30420_ (.A(_09904_),
    .B(_02859_),
    .Y(_09905_));
 sky130_fd_sc_hd__nor3_1 _30421_ (.A(\inst$top.soc.cpu.divider.timer[5] ),
    .B(\inst$top.soc.cpu.divider.timer[4] ),
    .C(_09905_),
    .Y(_09906_));
 sky130_fd_sc_hd__inv_1 _30422_ (.A(net1664),
    .Y(_09907_));
 sky130_fd_sc_hd__nand2_1 _30424_ (.A(net1245),
    .B(net2927),
    .Y(_09909_));
 sky130_fd_sc_hd__a21oi_4 _30427_ (.A1(net611),
    .A2(net1104),
    .B1(net2967),
    .Y(_03709_));
 sky130_fd_sc_hd__clkinv_1 _30428_ (.A(\inst$top.soc.cpu.sink__payload$12[144] ),
    .Y(_09912_));
 sky130_fd_sc_hd__o21ai_0 _30431_ (.A1(net2922),
    .A2(_09840_),
    .B1(net2112),
    .Y(_09915_));
 sky130_fd_sc_hd__a21oi_1 _30432_ (.A1(_09912_),
    .A2(_09840_),
    .B1(_09915_),
    .Y(_03710_));
 sky130_fd_sc_hd__inv_1 _30433_ (.A(_02922_),
    .Y(_09916_));
 sky130_fd_sc_hd__nor2_1 _30434_ (.A(\inst$top.soc.cpu.sink__payload$12[144] ),
    .B(\inst$top.soc.cpu.sink__payload$12[143] ),
    .Y(_09917_));
 sky130_fd_sc_hd__a32oi_1 _30435_ (.A1(\inst$top.soc.cpu.d.sink__payload.csr_fmt_i ),
    .A2(_09916_),
    .A3(_09917_),
    .B1(net1044),
    .B2(\inst$top.soc.cpu.sink__payload$12[144] ),
    .Y(_09918_));
 sky130_fd_sc_hd__o21ai_0 _30436_ (.A1(\inst$top.soc.cpu.divider.m_negative ),
    .A2(_09840_),
    .B1(net2112),
    .Y(_09919_));
 sky130_fd_sc_hd__a21oi_1 _30437_ (.A1(_09840_),
    .A2(_09918_),
    .B1(_09919_),
    .Y(_03711_));
 sky130_fd_sc_hd__inv_2 _30438_ (.A(net2931),
    .Y(_09920_));
 sky130_fd_sc_hd__nand3_1 _30440_ (.A(_09622_),
    .B(net2024),
    .C(_03082_),
    .Y(_09922_));
 sky130_fd_sc_hd__nor2_1 _30441_ (.A(net2026),
    .B(net1245),
    .Y(_09923_));
 sky130_fd_sc_hd__inv_1 _30443_ (.A(net1100),
    .Y(_09925_));
 sky130_fd_sc_hd__nand2_1 _30444_ (.A(_09839_),
    .B(net2023),
    .Y(_09926_));
 sky130_fd_sc_hd__o21ai_1 _30445_ (.A1(\inst$top.soc.cpu.divider.m_negative ),
    .A2(_09925_),
    .B1(_09926_),
    .Y(_09927_));
 sky130_fd_sc_hd__nor2_1 _30446_ (.A(net1102),
    .B(net749),
    .Y(_09928_));
 sky130_fd_sc_hd__nand4_4 _30447_ (.A(_09748_),
    .B(_09835_),
    .C(net2023),
    .D(_09800_),
    .Y(_09929_));
 sky130_fd_sc_hd__inv_1 _30448_ (.A(\inst$top.soc.cpu.divider.remainder[31] ),
    .Y(_09930_));
 sky130_fd_sc_hd__nand2_1 _30449_ (.A(_02825_),
    .B(_02828_),
    .Y(_09931_));
 sky130_fd_sc_hd__nand2_1 _30450_ (.A(_02837_),
    .B(_02840_),
    .Y(_09932_));
 sky130_fd_sc_hd__nand2_1 _30451_ (.A(_02831_),
    .B(_02834_),
    .Y(_09933_));
 sky130_fd_sc_hd__nor2_1 _30452_ (.A(_09932_),
    .B(_09933_),
    .Y(_09934_));
 sky130_fd_sc_hd__a21oi_1 _30453_ (.A1(_02837_),
    .A2(_02839_),
    .B1(_02836_),
    .Y(_09935_));
 sky130_fd_sc_hd__a21oi_1 _30454_ (.A1(_02831_),
    .A2(_02833_),
    .B1(_02830_),
    .Y(_09936_));
 sky130_fd_sc_hd__o21ai_0 _30455_ (.A1(_09933_),
    .A2(_09935_),
    .B1(_09936_),
    .Y(_09937_));
 sky130_fd_sc_hd__a21oi_1 _30456_ (.A1(_02543_),
    .A2(_09934_),
    .B1(_09937_),
    .Y(_09938_));
 sky130_fd_sc_hd__a21oi_1 _30457_ (.A1(_02825_),
    .A2(_02827_),
    .B1(_02824_),
    .Y(_09939_));
 sky130_fd_sc_hd__o21ai_0 _30458_ (.A1(_09931_),
    .A2(_09938_),
    .B1(_09939_),
    .Y(_09940_));
 sky130_fd_sc_hd__nand2_1 _30459_ (.A(_02813_),
    .B(_02816_),
    .Y(_09941_));
 sky130_fd_sc_hd__nand2_1 _30460_ (.A(_02819_),
    .B(_02822_),
    .Y(_09942_));
 sky130_fd_sc_hd__nand2_1 _30461_ (.A(_02801_),
    .B(_02804_),
    .Y(_09943_));
 sky130_fd_sc_hd__inv_1 _30462_ (.A(_09943_),
    .Y(_09944_));
 sky130_fd_sc_hd__nand2_1 _30463_ (.A(_02807_),
    .B(_02810_),
    .Y(_09945_));
 sky130_fd_sc_hd__inv_1 _30464_ (.A(_09945_),
    .Y(_09946_));
 sky130_fd_sc_hd__nand2_1 _30465_ (.A(_09944_),
    .B(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__nor3_1 _30466_ (.A(_09941_),
    .B(_09942_),
    .C(_09947_),
    .Y(_09948_));
 sky130_fd_sc_hd__nand2_1 _30467_ (.A(_02777_),
    .B(_02780_),
    .Y(_09949_));
 sky130_fd_sc_hd__nand2_1 _30468_ (.A(_02783_),
    .B(_02786_),
    .Y(_09950_));
 sky130_fd_sc_hd__nand2_1 _30469_ (.A(_02789_),
    .B(_02792_),
    .Y(_09951_));
 sky130_fd_sc_hd__nand2_1 _30470_ (.A(_02795_),
    .B(_02798_),
    .Y(_09952_));
 sky130_fd_sc_hd__nor4_1 _30471_ (.A(_09949_),
    .B(_09950_),
    .C(_09951_),
    .D(_09952_),
    .Y(_09953_));
 sky130_fd_sc_hd__nand3_1 _30472_ (.A(_09940_),
    .B(_09948_),
    .C(_09953_),
    .Y(_09954_));
 sky130_fd_sc_hd__a21oi_1 _30473_ (.A1(_02795_),
    .A2(_02797_),
    .B1(_02794_),
    .Y(_09955_));
 sky130_fd_sc_hd__a21oi_1 _30474_ (.A1(_02789_),
    .A2(_02791_),
    .B1(_02788_),
    .Y(_09956_));
 sky130_fd_sc_hd__o21ai_0 _30475_ (.A1(_09951_),
    .A2(_09955_),
    .B1(_09956_),
    .Y(_09957_));
 sky130_fd_sc_hd__nor2_1 _30476_ (.A(_09949_),
    .B(_09950_),
    .Y(_09958_));
 sky130_fd_sc_hd__a21oi_1 _30477_ (.A1(_02783_),
    .A2(_02785_),
    .B1(_02782_),
    .Y(_09959_));
 sky130_fd_sc_hd__a21oi_1 _30478_ (.A1(_02777_),
    .A2(_02779_),
    .B1(_02776_),
    .Y(_09960_));
 sky130_fd_sc_hd__o21ai_0 _30479_ (.A1(_09949_),
    .A2(_09959_),
    .B1(_09960_),
    .Y(_09961_));
 sky130_fd_sc_hd__a21oi_1 _30480_ (.A1(_09957_),
    .A2(_09958_),
    .B1(_09961_),
    .Y(_09962_));
 sky130_fd_sc_hd__a21oi_1 _30481_ (.A1(_02819_),
    .A2(_02821_),
    .B1(_02818_),
    .Y(_09963_));
 sky130_fd_sc_hd__inv_1 _30482_ (.A(_09963_),
    .Y(_09964_));
 sky130_fd_sc_hd__inv_1 _30483_ (.A(_09941_),
    .Y(_09965_));
 sky130_fd_sc_hd__a21oi_1 _30484_ (.A1(_02813_),
    .A2(_02815_),
    .B1(_02812_),
    .Y(_09966_));
 sky130_fd_sc_hd__inv_1 _30485_ (.A(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__a21oi_1 _30486_ (.A1(_09964_),
    .A2(_09965_),
    .B1(_09967_),
    .Y(_09968_));
 sky130_fd_sc_hd__a21oi_1 _30487_ (.A1(_02801_),
    .A2(_02803_),
    .B1(_02800_),
    .Y(_09969_));
 sky130_fd_sc_hd__nand2_1 _30488_ (.A(_02807_),
    .B(_02809_),
    .Y(_09970_));
 sky130_fd_sc_hd__inv_1 _30489_ (.A(_02806_),
    .Y(_09971_));
 sky130_fd_sc_hd__nand2_1 _30490_ (.A(_09970_),
    .B(_09971_),
    .Y(_09972_));
 sky130_fd_sc_hd__nand2_1 _30491_ (.A(_09972_),
    .B(_09944_),
    .Y(_09973_));
 sky130_fd_sc_hd__o211ai_1 _30492_ (.A1(_09947_),
    .A2(_09968_),
    .B1(_09969_),
    .C1(_09973_),
    .Y(_09974_));
 sky130_fd_sc_hd__nand2_1 _30493_ (.A(_09974_),
    .B(_09953_),
    .Y(_09975_));
 sky130_fd_sc_hd__nand3_1 _30494_ (.A(_09954_),
    .B(_09962_),
    .C(_09975_),
    .Y(_09976_));
 sky130_fd_sc_hd__nand2_1 _30495_ (.A(_02765_),
    .B(_02768_),
    .Y(_09977_));
 sky130_fd_sc_hd__nand2_1 _30496_ (.A(_02771_),
    .B(_02774_),
    .Y(_09978_));
 sky130_fd_sc_hd__nor2_1 _30497_ (.A(_09977_),
    .B(_09978_),
    .Y(_09979_));
 sky130_fd_sc_hd__a21oi_1 _30498_ (.A1(_02771_),
    .A2(_02773_),
    .B1(_02770_),
    .Y(_09980_));
 sky130_fd_sc_hd__a21oi_1 _30499_ (.A1(_02765_),
    .A2(_02767_),
    .B1(_02764_),
    .Y(_09981_));
 sky130_fd_sc_hd__o21ai_0 _30500_ (.A1(_09977_),
    .A2(_09980_),
    .B1(_09981_),
    .Y(_09982_));
 sky130_fd_sc_hd__a21o_1 _30501_ (.A1(_09976_),
    .A2(_09979_),
    .B1(_09982_),
    .X(_09983_));
 sky130_fd_sc_hd__inv_1 _30502_ (.A(_02753_),
    .Y(_09984_));
 sky130_fd_sc_hd__inv_1 _30503_ (.A(_02756_),
    .Y(_09985_));
 sky130_fd_sc_hd__nand2_1 _30504_ (.A(_02759_),
    .B(_02762_),
    .Y(_09986_));
 sky130_fd_sc_hd__nor3_1 _30505_ (.A(_09984_),
    .B(_09985_),
    .C(_09986_),
    .Y(_09987_));
 sky130_fd_sc_hd__a21oi_1 _30506_ (.A1(_02759_),
    .A2(_02761_),
    .B1(_02758_),
    .Y(_09988_));
 sky130_fd_sc_hd__a21oi_1 _30507_ (.A1(_02753_),
    .A2(_02755_),
    .B1(_02752_),
    .Y(_09989_));
 sky130_fd_sc_hd__o31ai_1 _30508_ (.A1(_09984_),
    .A2(_09985_),
    .A3(_09988_),
    .B1(_09989_),
    .Y(_09990_));
 sky130_fd_sc_hd__a21oi_1 _30509_ (.A1(_09983_),
    .A2(_09987_),
    .B1(_09990_),
    .Y(_09991_));
 sky130_fd_sc_hd__xor2_1 _30510_ (.A(_09930_),
    .B(_09991_),
    .X(_09992_));
 sky130_fd_sc_hd__inv_2 _30511_ (.A(net1104),
    .Y(_09993_));
 sky130_fd_sc_hd__nand2_1 _30513_ (.A(net856),
    .B(net1036),
    .Y(_09995_));
 sky130_fd_sc_hd__nand4_1 _30514_ (.A(_09922_),
    .B(_09928_),
    .C(_09929_),
    .D(_09995_),
    .Y(_09996_));
 sky130_fd_sc_hd__inv_1 _30515_ (.A(_09928_),
    .Y(_09997_));
 sky130_fd_sc_hd__a21oi_1 _30518_ (.A1(_09997_),
    .A2(_02846_),
    .B1(net2977),
    .Y(_10000_));
 sky130_fd_sc_hd__nand2_1 _30519_ (.A(_09996_),
    .B(_10000_),
    .Y(_10001_));
 sky130_fd_sc_hd__inv_2 _30520_ (.A(_10001_),
    .Y(_03712_));
 sky130_fd_sc_hd__nand2_1 _30522_ (.A(_09572_),
    .B(net2024),
    .Y(_10003_));
 sky130_fd_sc_hd__inv_1 _30523_ (.A(\inst$top.soc.cpu.divider.quotient[6] ),
    .Y(_10004_));
 sky130_fd_sc_hd__inv_1 _30524_ (.A(\inst$top.soc.cpu.divider.quotient[7] ),
    .Y(_10005_));
 sky130_fd_sc_hd__inv_1 _30525_ (.A(\inst$top.soc.cpu.divider.quotient[8] ),
    .Y(_10006_));
 sky130_fd_sc_hd__inv_1 _30526_ (.A(\inst$top.soc.cpu.divider.quotient[9] ),
    .Y(_10007_));
 sky130_fd_sc_hd__nand4_1 _30527_ (.A(_10004_),
    .B(_10005_),
    .C(_10006_),
    .D(_10007_),
    .Y(_10008_));
 sky130_fd_sc_hd__inv_1 _30528_ (.A(\inst$top.soc.cpu.divider.quotient[2] ),
    .Y(_10009_));
 sky130_fd_sc_hd__inv_1 _30529_ (.A(\inst$top.soc.cpu.divider.quotient[3] ),
    .Y(_10010_));
 sky130_fd_sc_hd__nand3_1 _30530_ (.A(_10009_),
    .B(_10010_),
    .C(_02848_),
    .Y(_10011_));
 sky130_fd_sc_hd__nor3_1 _30531_ (.A(\inst$top.soc.cpu.divider.quotient[4] ),
    .B(\inst$top.soc.cpu.divider.quotient[5] ),
    .C(_10011_),
    .Y(_10012_));
 sky130_fd_sc_hd__inv_1 _30532_ (.A(_10012_),
    .Y(_10013_));
 sky130_fd_sc_hd__nor2_1 _30533_ (.A(_10008_),
    .B(_10013_),
    .Y(_10014_));
 sky130_fd_sc_hd__inv_1 _30534_ (.A(_10014_),
    .Y(_10015_));
 sky130_fd_sc_hd__nand2_1 _30535_ (.A(_10015_),
    .B(\inst$top.soc.cpu.divider.quotient[10] ),
    .Y(_10016_));
 sky130_fd_sc_hd__inv_1 _30536_ (.A(\inst$top.soc.cpu.divider.quotient[10] ),
    .Y(_10017_));
 sky130_fd_sc_hd__nand2_1 _30537_ (.A(_10014_),
    .B(_10017_),
    .Y(_10018_));
 sky130_fd_sc_hd__a32oi_1 _30540_ (.A1(_10016_),
    .A2(_10018_),
    .A3(net1103),
    .B1(\inst$top.soc.cpu.divider.quotient[9] ),
    .B2(net1035),
    .Y(_10021_));
 sky130_fd_sc_hd__nand2_1 _30541_ (.A(_10003_),
    .B(_10021_),
    .Y(_10022_));
 sky130_fd_sc_hd__inv_1 _30542_ (.A(net749),
    .Y(_10023_));
 sky130_fd_sc_hd__nand2_2 _30543_ (.A(_09929_),
    .B(net725),
    .Y(_10024_));
 sky130_fd_sc_hd__a21oi_1 _30548_ (.A1(net744),
    .A2(_10017_),
    .B1(net2974),
    .Y(_10029_));
 sky130_fd_sc_hd__o21ai_1 _30549_ (.A1(_10022_),
    .A2(net609),
    .B1(_10029_),
    .Y(_10030_));
 sky130_fd_sc_hd__inv_2 _30550_ (.A(_10030_),
    .Y(_03713_));
 sky130_fd_sc_hd__inv_2 _30555_ (.A(net609),
    .Y(_10035_));
 sky130_fd_sc_hd__inv_1 _30556_ (.A(\inst$top.soc.cpu.divider.quotient[4] ),
    .Y(_10036_));
 sky130_fd_sc_hd__nand2_1 _30557_ (.A(_10010_),
    .B(_10036_),
    .Y(_10037_));
 sky130_fd_sc_hd__nand3_1 _30558_ (.A(_02847_),
    .B(_10009_),
    .C(_02846_),
    .Y(_10038_));
 sky130_fd_sc_hd__nor2_1 _30559_ (.A(_10037_),
    .B(_10038_),
    .Y(_10039_));
 sky130_fd_sc_hd__inv_1 _30560_ (.A(\inst$top.soc.cpu.divider.quotient[5] ),
    .Y(_10040_));
 sky130_fd_sc_hd__nand2_1 _30561_ (.A(_10039_),
    .B(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__nor2_1 _30562_ (.A(\inst$top.soc.cpu.divider.quotient[6] ),
    .B(_10041_),
    .Y(_10042_));
 sky130_fd_sc_hd__nand3_1 _30563_ (.A(_10042_),
    .B(_10005_),
    .C(_10006_),
    .Y(_10043_));
 sky130_fd_sc_hd__nor2_1 _30564_ (.A(\inst$top.soc.cpu.divider.quotient[9] ),
    .B(_10043_),
    .Y(_10044_));
 sky130_fd_sc_hd__inv_1 _30565_ (.A(\inst$top.soc.cpu.divider.quotient[11] ),
    .Y(_10045_));
 sky130_fd_sc_hd__a21oi_1 _30566_ (.A1(_10044_),
    .A2(_10017_),
    .B1(_10045_),
    .Y(_10046_));
 sky130_fd_sc_hd__nand3_1 _30567_ (.A(_10044_),
    .B(_10017_),
    .C(_10045_),
    .Y(_10047_));
 sky130_fd_sc_hd__nand2_1 _30568_ (.A(_10047_),
    .B(net1103),
    .Y(_10048_));
 sky130_fd_sc_hd__o22ai_1 _30569_ (.A1(_10017_),
    .A2(net1105),
    .B1(_10046_),
    .B2(_10048_),
    .Y(_10049_));
 sky130_fd_sc_hd__a21oi_1 _30570_ (.A1(_09576_),
    .A2(net2026),
    .B1(_10049_),
    .Y(_10050_));
 sky130_fd_sc_hd__nand2_1 _30571_ (.A(_10035_),
    .B(_10050_),
    .Y(_10051_));
 sky130_fd_sc_hd__o211ai_1 _30572_ (.A1(\inst$top.soc.cpu.divider.quotient[11] ),
    .A2(net723),
    .B1(net2117),
    .C1(_10051_),
    .Y(_10052_));
 sky130_fd_sc_hd__inv_2 _30573_ (.A(_10052_),
    .Y(_03714_));
 sky130_fd_sc_hd__nor3_1 _30574_ (.A(\inst$top.soc.cpu.divider.quotient[11] ),
    .B(\inst$top.soc.cpu.divider.quotient[12] ),
    .C(_10018_),
    .Y(_10053_));
 sky130_fd_sc_hd__o21ai_0 _30575_ (.A1(\inst$top.soc.cpu.divider.quotient[11] ),
    .A2(_10018_),
    .B1(\inst$top.soc.cpu.divider.quotient[12] ),
    .Y(_10054_));
 sky130_fd_sc_hd__nand2_1 _30576_ (.A(_10054_),
    .B(net1100),
    .Y(_10055_));
 sky130_fd_sc_hd__nand2_1 _30577_ (.A(_09568_),
    .B(net2026),
    .Y(_10056_));
 sky130_fd_sc_hd__o221ai_1 _30578_ (.A1(_10045_),
    .A2(_09909_),
    .B1(_10053_),
    .B2(_10055_),
    .C1(_10056_),
    .Y(_10057_));
 sky130_fd_sc_hd__inv_1 _30579_ (.A(\inst$top.soc.cpu.divider.quotient[12] ),
    .Y(_10058_));
 sky130_fd_sc_hd__a21oi_1 _30580_ (.A1(net744),
    .A2(_10058_),
    .B1(net2971),
    .Y(_10059_));
 sky130_fd_sc_hd__o21ai_1 _30581_ (.A1(_10057_),
    .A2(net609),
    .B1(_10059_),
    .Y(_10060_));
 sky130_fd_sc_hd__inv_2 _30582_ (.A(_10060_),
    .Y(_03715_));
 sky130_fd_sc_hd__nand4_1 _30583_ (.A(_10044_),
    .B(_10017_),
    .C(_10045_),
    .D(_10058_),
    .Y(_10061_));
 sky130_fd_sc_hd__nor2_1 _30584_ (.A(\inst$top.soc.cpu.divider.quotient[13] ),
    .B(_10061_),
    .Y(_10062_));
 sky130_fd_sc_hd__nand2_1 _30585_ (.A(_10061_),
    .B(\inst$top.soc.cpu.divider.quotient[13] ),
    .Y(_10063_));
 sky130_fd_sc_hd__nand2_1 _30586_ (.A(_10063_),
    .B(net1100),
    .Y(_10064_));
 sky130_fd_sc_hd__o22ai_1 _30587_ (.A1(_10058_),
    .A2(net1105),
    .B1(_10062_),
    .B2(_10064_),
    .Y(_10065_));
 sky130_fd_sc_hd__a21oi_1 _30588_ (.A1(_09565_),
    .A2(net2026),
    .B1(_10065_),
    .Y(_10066_));
 sky130_fd_sc_hd__nand2_1 _30589_ (.A(_10035_),
    .B(_10066_),
    .Y(_10067_));
 sky130_fd_sc_hd__o211ai_1 _30590_ (.A1(\inst$top.soc.cpu.divider.quotient[13] ),
    .A2(net723),
    .B1(net2100),
    .C1(_10067_),
    .Y(_10068_));
 sky130_fd_sc_hd__inv_2 _30591_ (.A(_10068_),
    .Y(_03716_));
 sky130_fd_sc_hd__nand2_1 _30592_ (.A(_09560_),
    .B(net2026),
    .Y(_10069_));
 sky130_fd_sc_hd__nor4_1 _30593_ (.A(\inst$top.soc.cpu.divider.quotient[10] ),
    .B(\inst$top.soc.cpu.divider.quotient[11] ),
    .C(\inst$top.soc.cpu.divider.quotient[12] ),
    .D(\inst$top.soc.cpu.divider.quotient[13] ),
    .Y(_10070_));
 sky130_fd_sc_hd__inv_1 _30594_ (.A(_10070_),
    .Y(_10071_));
 sky130_fd_sc_hd__o21ai_0 _30595_ (.A1(_10071_),
    .A2(_10015_),
    .B1(\inst$top.soc.cpu.divider.quotient[14] ),
    .Y(_10072_));
 sky130_fd_sc_hd__nor2_1 _30596_ (.A(_10071_),
    .B(_10015_),
    .Y(_10073_));
 sky130_fd_sc_hd__inv_1 _30597_ (.A(\inst$top.soc.cpu.divider.quotient[14] ),
    .Y(_10074_));
 sky130_fd_sc_hd__nand2_1 _30598_ (.A(_10073_),
    .B(_10074_),
    .Y(_10075_));
 sky130_fd_sc_hd__a32oi_1 _30599_ (.A1(_10072_),
    .A2(_10075_),
    .A3(net1100),
    .B1(\inst$top.soc.cpu.divider.quotient[13] ),
    .B2(net1035),
    .Y(_10076_));
 sky130_fd_sc_hd__nand2_1 _30600_ (.A(_10069_),
    .B(_10076_),
    .Y(_10077_));
 sky130_fd_sc_hd__a21oi_1 _30602_ (.A1(net744),
    .A2(_10074_),
    .B1(net2967),
    .Y(_10079_));
 sky130_fd_sc_hd__o21ai_1 _30603_ (.A1(_10077_),
    .A2(net609),
    .B1(_10079_),
    .Y(_10080_));
 sky130_fd_sc_hd__inv_2 _30604_ (.A(_10080_),
    .Y(_03717_));
 sky130_fd_sc_hd__nand2_1 _30606_ (.A(_10062_),
    .B(_10074_),
    .Y(_10082_));
 sky130_fd_sc_hd__nor2_1 _30607_ (.A(\inst$top.soc.cpu.divider.quotient[15] ),
    .B(_10082_),
    .Y(_10083_));
 sky130_fd_sc_hd__nand2_1 _30608_ (.A(_10082_),
    .B(\inst$top.soc.cpu.divider.quotient[15] ),
    .Y(_10084_));
 sky130_fd_sc_hd__nand2_1 _30609_ (.A(_10084_),
    .B(net1100),
    .Y(_10085_));
 sky130_fd_sc_hd__o22ai_1 _30610_ (.A1(_10074_),
    .A2(net1105),
    .B1(_10083_),
    .B2(_10085_),
    .Y(_10086_));
 sky130_fd_sc_hd__a21oi_1 _30611_ (.A1(net2026),
    .A2(_09556_),
    .B1(_10086_),
    .Y(_10087_));
 sky130_fd_sc_hd__nand2_1 _30612_ (.A(_10035_),
    .B(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__o211ai_1 _30613_ (.A1(\inst$top.soc.cpu.divider.quotient[15] ),
    .A2(net723),
    .B1(net2100),
    .C1(_10088_),
    .Y(_10089_));
 sky130_fd_sc_hd__inv_2 _30614_ (.A(_10089_),
    .Y(_03718_));
 sky130_fd_sc_hd__nand2_1 _30616_ (.A(_10012_),
    .B(_10004_),
    .Y(_10091_));
 sky130_fd_sc_hd__nor2_1 _30617_ (.A(\inst$top.soc.cpu.divider.quotient[7] ),
    .B(_10091_),
    .Y(_10092_));
 sky130_fd_sc_hd__nor4_1 _30618_ (.A(\inst$top.soc.cpu.divider.quotient[8] ),
    .B(\inst$top.soc.cpu.divider.quotient[9] ),
    .C(\inst$top.soc.cpu.divider.quotient[10] ),
    .D(\inst$top.soc.cpu.divider.quotient[11] ),
    .Y(_10093_));
 sky130_fd_sc_hd__nor4_1 _30619_ (.A(\inst$top.soc.cpu.divider.quotient[12] ),
    .B(\inst$top.soc.cpu.divider.quotient[13] ),
    .C(\inst$top.soc.cpu.divider.quotient[14] ),
    .D(\inst$top.soc.cpu.divider.quotient[15] ),
    .Y(_10094_));
 sky130_fd_sc_hd__nand3_1 _30620_ (.A(_10092_),
    .B(_10093_),
    .C(_10094_),
    .Y(_10095_));
 sky130_fd_sc_hd__inv_1 _30621_ (.A(_10095_),
    .Y(_10096_));
 sky130_fd_sc_hd__inv_1 _30622_ (.A(\inst$top.soc.cpu.divider.quotient[16] ),
    .Y(_10097_));
 sky130_fd_sc_hd__nand2_1 _30623_ (.A(_10096_),
    .B(_10097_),
    .Y(_10098_));
 sky130_fd_sc_hd__nand2_1 _30624_ (.A(_10095_),
    .B(\inst$top.soc.cpu.divider.quotient[16] ),
    .Y(_10099_));
 sky130_fd_sc_hd__a32oi_1 _30625_ (.A1(_10098_),
    .A2(_10099_),
    .A3(net1100),
    .B1(\inst$top.soc.cpu.divider.quotient[15] ),
    .B2(net1035),
    .Y(_10100_));
 sky130_fd_sc_hd__o21ai_0 _30626_ (.A1(net2925),
    .A2(_09605_),
    .B1(_10100_),
    .Y(_10101_));
 sky130_fd_sc_hd__a21oi_1 _30627_ (.A1(net744),
    .A2(_10097_),
    .B1(net2966),
    .Y(_10102_));
 sky130_fd_sc_hd__o21ai_1 _30628_ (.A1(_10101_),
    .A2(net609),
    .B1(_10102_),
    .Y(_10103_));
 sky130_fd_sc_hd__inv_2 _30629_ (.A(_10103_),
    .Y(_03719_));
 sky130_fd_sc_hd__nand2_1 _30630_ (.A(_10083_),
    .B(_10097_),
    .Y(_10104_));
 sky130_fd_sc_hd__nand2_1 _30631_ (.A(_10104_),
    .B(\inst$top.soc.cpu.divider.quotient[17] ),
    .Y(_10105_));
 sky130_fd_sc_hd__inv_1 _30633_ (.A(\inst$top.soc.cpu.divider.quotient[17] ),
    .Y(_10107_));
 sky130_fd_sc_hd__nand3_1 _30634_ (.A(_10083_),
    .B(_10097_),
    .C(_10107_),
    .Y(_10108_));
 sky130_fd_sc_hd__nand3_1 _30635_ (.A(_10105_),
    .B(net1100),
    .C(_10108_),
    .Y(_10109_));
 sky130_fd_sc_hd__nand2_1 _30637_ (.A(net1035),
    .B(\inst$top.soc.cpu.divider.quotient[16] ),
    .Y(_10111_));
 sky130_fd_sc_hd__nand3_1 _30638_ (.A(_09617_),
    .B(net2023),
    .C(_09618_),
    .Y(_10112_));
 sky130_fd_sc_hd__nand3_1 _30639_ (.A(_10109_),
    .B(_10111_),
    .C(_10112_),
    .Y(_10113_));
 sky130_fd_sc_hd__a21oi_1 _30640_ (.A1(net744),
    .A2(_10107_),
    .B1(net2964),
    .Y(_10114_));
 sky130_fd_sc_hd__o21ai_1 _30641_ (.A1(_10113_),
    .A2(net609),
    .B1(_10114_),
    .Y(_10115_));
 sky130_fd_sc_hd__inv_2 _30642_ (.A(_10115_),
    .Y(_03720_));
 sky130_fd_sc_hd__nor4_1 _30643_ (.A(\inst$top.soc.cpu.divider.quotient[14] ),
    .B(\inst$top.soc.cpu.divider.quotient[15] ),
    .C(\inst$top.soc.cpu.divider.quotient[16] ),
    .D(\inst$top.soc.cpu.divider.quotient[17] ),
    .Y(_10116_));
 sky130_fd_sc_hd__nand2_1 _30644_ (.A(_10073_),
    .B(_10116_),
    .Y(_10117_));
 sky130_fd_sc_hd__nand2_1 _30645_ (.A(_10117_),
    .B(\inst$top.soc.cpu.divider.quotient[18] ),
    .Y(_10118_));
 sky130_fd_sc_hd__inv_1 _30646_ (.A(\inst$top.soc.cpu.divider.quotient[18] ),
    .Y(_10119_));
 sky130_fd_sc_hd__nand3_1 _30647_ (.A(_10073_),
    .B(_10119_),
    .C(_10116_),
    .Y(_10120_));
 sky130_fd_sc_hd__a32oi_1 _30648_ (.A1(_10118_),
    .A2(_10120_),
    .A3(net1100),
    .B1(\inst$top.soc.cpu.divider.quotient[17] ),
    .B2(net1035),
    .Y(_10121_));
 sky130_fd_sc_hd__o21ai_0 _30649_ (.A1(net2931),
    .A2(_09610_),
    .B1(_10121_),
    .Y(_10122_));
 sky130_fd_sc_hd__a21oi_1 _30652_ (.A1(net744),
    .A2(_10119_),
    .B1(net2966),
    .Y(_10125_));
 sky130_fd_sc_hd__o21ai_1 _30653_ (.A1(_10122_),
    .A2(net609),
    .B1(_10125_),
    .Y(_10126_));
 sky130_fd_sc_hd__inv_2 _30654_ (.A(_10126_),
    .Y(_03721_));
 sky130_fd_sc_hd__inv_1 _30656_ (.A(\inst$top.soc.cpu.divider.quotient[19] ),
    .Y(_10128_));
 sky130_fd_sc_hd__nor2_1 _30657_ (.A(\inst$top.soc.cpu.divider.quotient[15] ),
    .B(\inst$top.soc.cpu.divider.quotient[16] ),
    .Y(_10129_));
 sky130_fd_sc_hd__nand3_1 _30658_ (.A(_10129_),
    .B(_10107_),
    .C(_10119_),
    .Y(_10130_));
 sky130_fd_sc_hd__nor2_1 _30659_ (.A(_10130_),
    .B(_10082_),
    .Y(_10131_));
 sky130_fd_sc_hd__a21oi_1 _30660_ (.A1(_10131_),
    .A2(_10128_),
    .B1(_09925_),
    .Y(_10132_));
 sky130_fd_sc_hd__o21ai_0 _30661_ (.A1(_10128_),
    .A2(_10131_),
    .B1(_10132_),
    .Y(_10133_));
 sky130_fd_sc_hd__o221ai_1 _30662_ (.A1(net2925),
    .A2(_09614_),
    .B1(_10119_),
    .B2(_09909_),
    .C1(_10133_),
    .Y(_10134_));
 sky130_fd_sc_hd__a21oi_1 _30663_ (.A1(net744),
    .A2(_10128_),
    .B1(net2972),
    .Y(_10135_));
 sky130_fd_sc_hd__o21ai_1 _30664_ (.A1(_10134_),
    .A2(net609),
    .B1(_10135_),
    .Y(_10136_));
 sky130_fd_sc_hd__inv_2 _30665_ (.A(_10136_),
    .Y(_03722_));
 sky130_fd_sc_hd__nand2_1 _30666_ (.A(net1043),
    .B(_02845_),
    .Y(_10137_));
 sky130_fd_sc_hd__o21ai_0 _30667_ (.A1(net1706),
    .A2(net1043),
    .B1(_10137_),
    .Y(_10138_));
 sky130_fd_sc_hd__nand3_1 _30668_ (.A(_09622_),
    .B(net2024),
    .C(_10138_),
    .Y(_10139_));
 sky130_fd_sc_hd__a22oi_1 _30670_ (.A1(net1102),
    .A2(_02849_),
    .B1(net1037),
    .B2(\inst$top.soc.cpu.divider.quotient[0] ),
    .Y(_10141_));
 sky130_fd_sc_hd__nand4_1 _30671_ (.A(_10139_),
    .B(net726),
    .C(_09929_),
    .D(_10141_),
    .Y(_10142_));
 sky130_fd_sc_hd__a21oi_1 _30674_ (.A1(net748),
    .A2(_02847_),
    .B1(net2977),
    .Y(_10145_));
 sky130_fd_sc_hd__nand2_1 _30675_ (.A(_10142_),
    .B(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__inv_2 _30676_ (.A(_10146_),
    .Y(_03723_));
 sky130_fd_sc_hd__nor4_1 _30678_ (.A(\inst$top.soc.cpu.divider.quotient[16] ),
    .B(\inst$top.soc.cpu.divider.quotient[17] ),
    .C(\inst$top.soc.cpu.divider.quotient[18] ),
    .D(\inst$top.soc.cpu.divider.quotient[19] ),
    .Y(_10148_));
 sky130_fd_sc_hd__nand2_1 _30679_ (.A(_10096_),
    .B(_10148_),
    .Y(_10149_));
 sky130_fd_sc_hd__xor2_1 _30680_ (.A(\inst$top.soc.cpu.divider.quotient[20] ),
    .B(_10149_),
    .X(_10150_));
 sky130_fd_sc_hd__a22oi_1 _30681_ (.A1(\inst$top.soc.cpu.divider.quotient[19] ),
    .A2(net1036),
    .B1(_10150_),
    .B2(net1101),
    .Y(_10151_));
 sky130_fd_sc_hd__o21ai_0 _30682_ (.A1(net2925),
    .A2(_09596_),
    .B1(_10151_),
    .Y(_10152_));
 sky130_fd_sc_hd__inv_1 _30683_ (.A(\inst$top.soc.cpu.divider.quotient[20] ),
    .Y(_10153_));
 sky130_fd_sc_hd__a21oi_1 _30684_ (.A1(net747),
    .A2(_10153_),
    .B1(net2972),
    .Y(_10154_));
 sky130_fd_sc_hd__o21ai_1 _30685_ (.A1(_10152_),
    .A2(net610),
    .B1(_10154_),
    .Y(_10155_));
 sky130_fd_sc_hd__inv_2 _30686_ (.A(_10155_),
    .Y(_03724_));
 sky130_fd_sc_hd__nand2_1 _30687_ (.A(_10131_),
    .B(_10128_),
    .Y(_10156_));
 sky130_fd_sc_hd__o21ai_0 _30688_ (.A1(\inst$top.soc.cpu.divider.quotient[20] ),
    .A2(_10156_),
    .B1(\inst$top.soc.cpu.divider.quotient[21] ),
    .Y(_10157_));
 sky130_fd_sc_hd__inv_1 _30689_ (.A(\inst$top.soc.cpu.divider.quotient[21] ),
    .Y(_10158_));
 sky130_fd_sc_hd__nand4_1 _30690_ (.A(_10131_),
    .B(_10128_),
    .C(_10153_),
    .D(_10158_),
    .Y(_10159_));
 sky130_fd_sc_hd__o22ai_1 _30691_ (.A1(_10153_),
    .A2(net1105),
    .B1(net2928),
    .B2(_09592_),
    .Y(_10160_));
 sky130_fd_sc_hd__a31oi_1 _30692_ (.A1(_10157_),
    .A2(_10159_),
    .A3(net1101),
    .B1(_10160_),
    .Y(_10161_));
 sky130_fd_sc_hd__nand2_1 _30693_ (.A(_10035_),
    .B(_10161_),
    .Y(_10162_));
 sky130_fd_sc_hd__o211ai_1 _30694_ (.A1(\inst$top.soc.cpu.divider.quotient[21] ),
    .A2(net725),
    .B1(net2110),
    .C1(_10162_),
    .Y(_10163_));
 sky130_fd_sc_hd__inv_2 _30695_ (.A(_10163_),
    .Y(_03725_));
 sky130_fd_sc_hd__nand2_1 _30696_ (.A(_09601_),
    .B(net2023),
    .Y(_10164_));
 sky130_fd_sc_hd__nor2_1 _30697_ (.A(\inst$top.soc.cpu.divider.quotient[20] ),
    .B(\inst$top.soc.cpu.divider.quotient[21] ),
    .Y(_10165_));
 sky130_fd_sc_hd__nand3_1 _30698_ (.A(_10165_),
    .B(_10119_),
    .C(_10128_),
    .Y(_10166_));
 sky130_fd_sc_hd__o21ai_0 _30699_ (.A1(_10166_),
    .A2(_10117_),
    .B1(\inst$top.soc.cpu.divider.quotient[22] ),
    .Y(_10167_));
 sky130_fd_sc_hd__nor2_1 _30700_ (.A(_10166_),
    .B(_10117_),
    .Y(_10168_));
 sky130_fd_sc_hd__inv_1 _30701_ (.A(\inst$top.soc.cpu.divider.quotient[22] ),
    .Y(_10169_));
 sky130_fd_sc_hd__nand2_1 _30702_ (.A(_10168_),
    .B(_10169_),
    .Y(_10170_));
 sky130_fd_sc_hd__a32oi_1 _30703_ (.A1(_10167_),
    .A2(_10170_),
    .A3(net1101),
    .B1(\inst$top.soc.cpu.divider.quotient[21] ),
    .B2(net1036),
    .Y(_10171_));
 sky130_fd_sc_hd__nand2_1 _30704_ (.A(_10164_),
    .B(_10171_),
    .Y(_10172_));
 sky130_fd_sc_hd__a21oi_1 _30705_ (.A1(net747),
    .A2(_10169_),
    .B1(net2972),
    .Y(_10173_));
 sky130_fd_sc_hd__o21ai_1 _30706_ (.A1(_10172_),
    .A2(net610),
    .B1(_10173_),
    .Y(_10174_));
 sky130_fd_sc_hd__inv_2 _30707_ (.A(_10174_),
    .Y(_03726_));
 sky130_fd_sc_hd__o21ai_0 _30708_ (.A1(\inst$top.soc.cpu.divider.quotient[22] ),
    .A2(_10159_),
    .B1(\inst$top.soc.cpu.divider.quotient[23] ),
    .Y(_10175_));
 sky130_fd_sc_hd__inv_1 _30709_ (.A(\inst$top.soc.cpu.divider.quotient[23] ),
    .Y(_10176_));
 sky130_fd_sc_hd__nand4_1 _30710_ (.A(_10128_),
    .B(_10153_),
    .C(_10158_),
    .D(_10169_),
    .Y(_10177_));
 sky130_fd_sc_hd__inv_1 _30711_ (.A(_10177_),
    .Y(_10178_));
 sky130_fd_sc_hd__nand3_1 _30712_ (.A(_10131_),
    .B(_10176_),
    .C(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__nand3_1 _30713_ (.A(_10175_),
    .B(net1101),
    .C(_10179_),
    .Y(_10180_));
 sky130_fd_sc_hd__nand2_1 _30714_ (.A(net1036),
    .B(\inst$top.soc.cpu.divider.quotient[22] ),
    .Y(_10181_));
 sky130_fd_sc_hd__nand2_1 _30715_ (.A(_09600_),
    .B(net2023),
    .Y(_10182_));
 sky130_fd_sc_hd__nand4_1 _30716_ (.A(_09929_),
    .B(_10180_),
    .C(_10181_),
    .D(_10182_),
    .Y(_10183_));
 sky130_fd_sc_hd__a21oi_1 _30717_ (.A1(net747),
    .A2(_10176_),
    .B1(net2972),
    .Y(_10184_));
 sky130_fd_sc_hd__o21ai_0 _30718_ (.A1(net747),
    .A2(_10183_),
    .B1(_10184_),
    .Y(_10185_));
 sky130_fd_sc_hd__inv_2 _30719_ (.A(_10185_),
    .Y(_03727_));
 sky130_fd_sc_hd__inv_1 _30720_ (.A(\inst$top.soc.cpu.divider.quotient[24] ),
    .Y(_10186_));
 sky130_fd_sc_hd__nand3_1 _30721_ (.A(_10165_),
    .B(_10169_),
    .C(_10176_),
    .Y(_10187_));
 sky130_fd_sc_hd__nor2_1 _30722_ (.A(_10187_),
    .B(_10149_),
    .Y(_10188_));
 sky130_fd_sc_hd__xor2_1 _30723_ (.A(_10186_),
    .B(_10188_),
    .X(_10189_));
 sky130_fd_sc_hd__a22oi_1 _30724_ (.A1(\inst$top.soc.cpu.divider.quotient[23] ),
    .A2(net1036),
    .B1(_10189_),
    .B2(net1101),
    .Y(_10190_));
 sky130_fd_sc_hd__o211ai_1 _30725_ (.A1(net2930),
    .A2(_09455_),
    .B1(_10190_),
    .C1(_09929_),
    .Y(_10191_));
 sky130_fd_sc_hd__a21oi_1 _30726_ (.A1(net747),
    .A2(_10186_),
    .B1(net2972),
    .Y(_10192_));
 sky130_fd_sc_hd__o21ai_0 _30727_ (.A1(net747),
    .A2(_10191_),
    .B1(_10192_),
    .Y(_10193_));
 sky130_fd_sc_hd__inv_2 _30728_ (.A(_10193_),
    .Y(_03728_));
 sky130_fd_sc_hd__inv_1 _30730_ (.A(\inst$top.soc.cpu.divider.quotient[25] ),
    .Y(_10195_));
 sky130_fd_sc_hd__nor2_1 _30731_ (.A(\inst$top.soc.cpu.divider.quotient[24] ),
    .B(_10179_),
    .Y(_10196_));
 sky130_fd_sc_hd__xor2_1 _30732_ (.A(_10195_),
    .B(_10196_),
    .X(_10197_));
 sky130_fd_sc_hd__a22oi_1 _30733_ (.A1(\inst$top.soc.cpu.divider.quotient[24] ),
    .A2(net1037),
    .B1(_10197_),
    .B2(net1101),
    .Y(_10198_));
 sky130_fd_sc_hd__nand3_1 _30734_ (.A(_09499_),
    .B(net2023),
    .C(_09500_),
    .Y(_10199_));
 sky130_fd_sc_hd__nand3_1 _30735_ (.A(_10198_),
    .B(_09929_),
    .C(_10199_),
    .Y(_10200_));
 sky130_fd_sc_hd__a21oi_1 _30736_ (.A1(net748),
    .A2(_10195_),
    .B1(net2973),
    .Y(_10201_));
 sky130_fd_sc_hd__o21ai_0 _30737_ (.A1(net748),
    .A2(_10200_),
    .B1(_10201_),
    .Y(_10202_));
 sky130_fd_sc_hd__inv_2 _30738_ (.A(_10202_),
    .Y(_03729_));
 sky130_fd_sc_hd__nor4_1 _30739_ (.A(\inst$top.soc.cpu.divider.quotient[22] ),
    .B(\inst$top.soc.cpu.divider.quotient[23] ),
    .C(\inst$top.soc.cpu.divider.quotient[24] ),
    .D(\inst$top.soc.cpu.divider.quotient[25] ),
    .Y(_10203_));
 sky130_fd_sc_hd__nand2_1 _30740_ (.A(_10168_),
    .B(_10203_),
    .Y(_10204_));
 sky130_fd_sc_hd__xor2_1 _30741_ (.A(\inst$top.soc.cpu.divider.quotient[26] ),
    .B(_10204_),
    .X(_10205_));
 sky130_fd_sc_hd__a22oi_1 _30742_ (.A1(\inst$top.soc.cpu.divider.quotient[25] ),
    .A2(net1036),
    .B1(_10205_),
    .B2(net1101),
    .Y(_10206_));
 sky130_fd_sc_hd__o211ai_1 _30743_ (.A1(net2930),
    .A2(_09473_),
    .B1(_10206_),
    .C1(_09929_),
    .Y(_10207_));
 sky130_fd_sc_hd__inv_1 _30745_ (.A(\inst$top.soc.cpu.divider.quotient[26] ),
    .Y(_10209_));
 sky130_fd_sc_hd__a21oi_1 _30746_ (.A1(net747),
    .A2(_10209_),
    .B1(net2972),
    .Y(_10210_));
 sky130_fd_sc_hd__o21ai_0 _30747_ (.A1(net747),
    .A2(_10207_),
    .B1(_10210_),
    .Y(_10211_));
 sky130_fd_sc_hd__inv_2 _30748_ (.A(_10211_),
    .Y(_03730_));
 sky130_fd_sc_hd__nor4_1 _30749_ (.A(\inst$top.soc.cpu.divider.quotient[23] ),
    .B(\inst$top.soc.cpu.divider.quotient[24] ),
    .C(\inst$top.soc.cpu.divider.quotient[25] ),
    .D(\inst$top.soc.cpu.divider.quotient[26] ),
    .Y(_10212_));
 sky130_fd_sc_hd__nand3_1 _30750_ (.A(_10131_),
    .B(_10178_),
    .C(_10212_),
    .Y(_10213_));
 sky130_fd_sc_hd__inv_1 _30751_ (.A(_10213_),
    .Y(_10214_));
 sky130_fd_sc_hd__inv_1 _30752_ (.A(\inst$top.soc.cpu.divider.quotient[27] ),
    .Y(_10215_));
 sky130_fd_sc_hd__nand2_1 _30753_ (.A(_10214_),
    .B(_10215_),
    .Y(_10216_));
 sky130_fd_sc_hd__nand2_1 _30754_ (.A(_10213_),
    .B(\inst$top.soc.cpu.divider.quotient[27] ),
    .Y(_10217_));
 sky130_fd_sc_hd__nand3_1 _30755_ (.A(_10216_),
    .B(net1102),
    .C(_10217_),
    .Y(_10218_));
 sky130_fd_sc_hd__nand2_1 _30756_ (.A(net1037),
    .B(\inst$top.soc.cpu.divider.quotient[26] ),
    .Y(_10219_));
 sky130_fd_sc_hd__nand3_1 _30757_ (.A(_09494_),
    .B(net2023),
    .C(_09495_),
    .Y(_10220_));
 sky130_fd_sc_hd__nand4_1 _30758_ (.A(_10035_),
    .B(_10218_),
    .C(_10219_),
    .D(_10220_),
    .Y(_10221_));
 sky130_fd_sc_hd__a21oi_1 _30759_ (.A1(net748),
    .A2(_10215_),
    .B1(net2972),
    .Y(_10222_));
 sky130_fd_sc_hd__nand2_1 _30760_ (.A(_10221_),
    .B(_10222_),
    .Y(_10223_));
 sky130_fd_sc_hd__inv_2 _30761_ (.A(_10223_),
    .Y(_03731_));
 sky130_fd_sc_hd__inv_1 _30762_ (.A(\inst$top.soc.cpu.divider.quotient[28] ),
    .Y(_10224_));
 sky130_fd_sc_hd__nand4_1 _30763_ (.A(_10203_),
    .B(_10209_),
    .C(_10215_),
    .D(_10165_),
    .Y(_10225_));
 sky130_fd_sc_hd__nor2_1 _30764_ (.A(_10225_),
    .B(_10149_),
    .Y(_10226_));
 sky130_fd_sc_hd__xor2_1 _30765_ (.A(_10224_),
    .B(_10226_),
    .X(_10227_));
 sky130_fd_sc_hd__a22oi_1 _30766_ (.A1(\inst$top.soc.cpu.divider.quotient[27] ),
    .A2(net1036),
    .B1(_10227_),
    .B2(net1101),
    .Y(_10228_));
 sky130_fd_sc_hd__o211ai_1 _30767_ (.A1(net2930),
    .A2(_09535_),
    .B1(_10228_),
    .C1(_09929_),
    .Y(_10229_));
 sky130_fd_sc_hd__a21oi_1 _30768_ (.A1(net748),
    .A2(_10224_),
    .B1(net2973),
    .Y(_10230_));
 sky130_fd_sc_hd__o21ai_0 _30769_ (.A1(net748),
    .A2(_10229_),
    .B1(_10230_),
    .Y(_10231_));
 sky130_fd_sc_hd__inv_2 _30770_ (.A(_10231_),
    .Y(_03732_));
 sky130_fd_sc_hd__o21ai_0 _30771_ (.A1(\inst$top.soc.cpu.divider.quotient[28] ),
    .A2(_10216_),
    .B1(\inst$top.soc.cpu.divider.quotient[29] ),
    .Y(_10232_));
 sky130_fd_sc_hd__inv_1 _30772_ (.A(\inst$top.soc.cpu.divider.quotient[29] ),
    .Y(_10233_));
 sky130_fd_sc_hd__nand4_1 _30773_ (.A(_10214_),
    .B(_10215_),
    .C(_10224_),
    .D(_10233_),
    .Y(_10234_));
 sky130_fd_sc_hd__nand3_1 _30774_ (.A(_10232_),
    .B(net1102),
    .C(_10234_),
    .Y(_10235_));
 sky130_fd_sc_hd__nand2_1 _30775_ (.A(net1037),
    .B(\inst$top.soc.cpu.divider.quotient[28] ),
    .Y(_10236_));
 sky130_fd_sc_hd__nand2_1 _30776_ (.A(_09526_),
    .B(net2023),
    .Y(_10237_));
 sky130_fd_sc_hd__nand4_1 _30777_ (.A(_10035_),
    .B(_10235_),
    .C(_10236_),
    .D(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__a21oi_1 _30778_ (.A1(net747),
    .A2(_10233_),
    .B1(net2972),
    .Y(_10239_));
 sky130_fd_sc_hd__nand2_1 _30779_ (.A(_10238_),
    .B(_10239_),
    .Y(_10240_));
 sky130_fd_sc_hd__inv_2 _30780_ (.A(_10240_),
    .Y(_03733_));
 sky130_fd_sc_hd__xor2_1 _30781_ (.A(\inst$top.soc.cpu.divider.quotient[2] ),
    .B(_02848_),
    .X(_10241_));
 sky130_fd_sc_hd__nand2_1 _30782_ (.A(net1041),
    .B(_09550_),
    .Y(_10242_));
 sky130_fd_sc_hd__xor2_1 _30783_ (.A(net1366),
    .B(_10242_),
    .X(_10243_));
 sky130_fd_sc_hd__nand2_1 _30784_ (.A(_10243_),
    .B(net2024),
    .Y(_10244_));
 sky130_fd_sc_hd__o221ai_1 _30785_ (.A1(_02847_),
    .A2(net1105),
    .B1(_09925_),
    .B2(_10241_),
    .C1(_10244_),
    .Y(_10245_));
 sky130_fd_sc_hd__a21oi_1 _30786_ (.A1(net748),
    .A2(_10009_),
    .B1(net2975),
    .Y(_10246_));
 sky130_fd_sc_hd__o21ai_1 _30787_ (.A1(_10245_),
    .A2(net610),
    .B1(_10246_),
    .Y(_10247_));
 sky130_fd_sc_hd__inv_2 _30788_ (.A(_10247_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand2_1 _30789_ (.A(_09518_),
    .B(net2023),
    .Y(_10248_));
 sky130_fd_sc_hd__inv_1 _30790_ (.A(\inst$top.soc.cpu.divider.quotient[30] ),
    .Y(_10249_));
 sky130_fd_sc_hd__nor2_1 _30791_ (.A(\inst$top.soc.cpu.divider.quotient[27] ),
    .B(\inst$top.soc.cpu.divider.quotient[28] ),
    .Y(_10250_));
 sky130_fd_sc_hd__nand3_1 _30792_ (.A(_10250_),
    .B(_10209_),
    .C(_10233_),
    .Y(_10251_));
 sky130_fd_sc_hd__nor2_1 _30793_ (.A(_10251_),
    .B(_10204_),
    .Y(_10252_));
 sky130_fd_sc_hd__xor2_1 _30794_ (.A(_10249_),
    .B(_10252_),
    .X(_10253_));
 sky130_fd_sc_hd__a22oi_1 _30795_ (.A1(\inst$top.soc.cpu.divider.quotient[29] ),
    .A2(net1037),
    .B1(_10253_),
    .B2(net1101),
    .Y(_10254_));
 sky130_fd_sc_hd__nand4_1 _30796_ (.A(_09929_),
    .B(net726),
    .C(_10248_),
    .D(_10254_),
    .Y(_10255_));
 sky130_fd_sc_hd__o211ai_1 _30797_ (.A1(\inst$top.soc.cpu.divider.quotient[30] ),
    .A2(net726),
    .B1(net2112),
    .C1(_10255_),
    .Y(_10256_));
 sky130_fd_sc_hd__inv_2 _30798_ (.A(_10256_),
    .Y(_03735_));
 sky130_fd_sc_hd__nand3_1 _30799_ (.A(_10250_),
    .B(_10233_),
    .C(_10249_),
    .Y(_10257_));
 sky130_fd_sc_hd__nor2_1 _30800_ (.A(_10257_),
    .B(_10213_),
    .Y(_10258_));
 sky130_fd_sc_hd__a21oi_1 _30801_ (.A1(_10258_),
    .A2(_02850_),
    .B1(_09925_),
    .Y(_10259_));
 sky130_fd_sc_hd__o21ai_0 _30802_ (.A1(_02850_),
    .A2(_10258_),
    .B1(_10259_),
    .Y(_10260_));
 sky130_fd_sc_hd__nand2_1 _30803_ (.A(net1037),
    .B(\inst$top.soc.cpu.divider.quotient[30] ),
    .Y(_10261_));
 sky130_fd_sc_hd__nand2_1 _30804_ (.A(_09507_),
    .B(net2023),
    .Y(_10262_));
 sky130_fd_sc_hd__nand4_1 _30805_ (.A(_10035_),
    .B(_10260_),
    .C(_10261_),
    .D(_10262_),
    .Y(_10263_));
 sky130_fd_sc_hd__a21oi_1 _30806_ (.A1(net747),
    .A2(_02850_),
    .B1(net2972),
    .Y(_10264_));
 sky130_fd_sc_hd__nand2_1 _30807_ (.A(_10263_),
    .B(_10264_),
    .Y(_10265_));
 sky130_fd_sc_hd__inv_2 _30808_ (.A(_10265_),
    .Y(_03736_));
 sky130_fd_sc_hd__xor2_1 _30809_ (.A(_10010_),
    .B(_10038_),
    .X(_10266_));
 sky130_fd_sc_hd__o22ai_1 _30810_ (.A1(_10009_),
    .A2(net1105),
    .B1(_10266_),
    .B2(_09925_),
    .Y(_10267_));
 sky130_fd_sc_hd__a21oi_1 _30811_ (.A1(_09552_),
    .A2(net2025),
    .B1(_10267_),
    .Y(_10268_));
 sky130_fd_sc_hd__nand2_1 _30812_ (.A(_10035_),
    .B(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__o211ai_1 _30813_ (.A1(\inst$top.soc.cpu.divider.quotient[3] ),
    .A2(net726),
    .B1(net2117),
    .C1(_10269_),
    .Y(_10270_));
 sky130_fd_sc_hd__inv_2 _30814_ (.A(_10270_),
    .Y(_03737_));
 sky130_fd_sc_hd__xor2_1 _30815_ (.A(\inst$top.soc.cpu.divider.quotient[4] ),
    .B(_10011_),
    .X(_10271_));
 sky130_fd_sc_hd__a22oi_1 _30816_ (.A1(net1102),
    .A2(_10271_),
    .B1(net1036),
    .B2(\inst$top.soc.cpu.divider.quotient[3] ),
    .Y(_10272_));
 sky130_fd_sc_hd__o21ai_0 _30817_ (.A1(net2928),
    .A2(_09543_),
    .B1(_10272_),
    .Y(_10273_));
 sky130_fd_sc_hd__a21oi_1 _30819_ (.A1(net748),
    .A2(_10036_),
    .B1(net2975),
    .Y(_10275_));
 sky130_fd_sc_hd__o21ai_0 _30820_ (.A1(_10273_),
    .A2(net609),
    .B1(_10275_),
    .Y(_10276_));
 sky130_fd_sc_hd__inv_2 _30821_ (.A(_10276_),
    .Y(_03738_));
 sky130_fd_sc_hd__o21ai_0 _30822_ (.A1(_10037_),
    .A2(_10038_),
    .B1(\inst$top.soc.cpu.divider.quotient[5] ),
    .Y(_10277_));
 sky130_fd_sc_hd__a32oi_1 _30823_ (.A1(net1101),
    .A2(_10041_),
    .A3(_10277_),
    .B1(\inst$top.soc.cpu.divider.quotient[4] ),
    .B2(net1036),
    .Y(_10278_));
 sky130_fd_sc_hd__o21ai_0 _30824_ (.A1(net2928),
    .A2(_09541_),
    .B1(_10278_),
    .Y(_10279_));
 sky130_fd_sc_hd__a21oi_1 _30825_ (.A1(net748),
    .A2(_10040_),
    .B1(net2975),
    .Y(_10280_));
 sky130_fd_sc_hd__o21ai_0 _30826_ (.A1(_10279_),
    .A2(net610),
    .B1(_10280_),
    .Y(_10281_));
 sky130_fd_sc_hd__inv_2 _30827_ (.A(_10281_),
    .Y(_03739_));
 sky130_fd_sc_hd__nand2_1 _30828_ (.A(_09546_),
    .B(net2024),
    .Y(_10282_));
 sky130_fd_sc_hd__nand2_1 _30829_ (.A(_10013_),
    .B(\inst$top.soc.cpu.divider.quotient[6] ),
    .Y(_10283_));
 sky130_fd_sc_hd__a32oi_1 _30830_ (.A1(net1100),
    .A2(_10283_),
    .A3(_10091_),
    .B1(\inst$top.soc.cpu.divider.quotient[5] ),
    .B2(net1036),
    .Y(_10284_));
 sky130_fd_sc_hd__nand2_1 _30831_ (.A(_10282_),
    .B(_10284_),
    .Y(_10285_));
 sky130_fd_sc_hd__a21oi_1 _30832_ (.A1(net746),
    .A2(_10004_),
    .B1(net2974),
    .Y(_10286_));
 sky130_fd_sc_hd__o21ai_0 _30833_ (.A1(_10285_),
    .A2(net610),
    .B1(_10286_),
    .Y(_10287_));
 sky130_fd_sc_hd__inv_2 _30834_ (.A(_10287_),
    .Y(_03740_));
 sky130_fd_sc_hd__xor2_1 _30835_ (.A(\inst$top.soc.cpu.divider.quotient[7] ),
    .B(_10042_),
    .X(_10288_));
 sky130_fd_sc_hd__o22ai_1 _30836_ (.A1(_10004_),
    .A2(net1105),
    .B1(_09925_),
    .B2(_10288_),
    .Y(_10289_));
 sky130_fd_sc_hd__a21oi_1 _30837_ (.A1(_09548_),
    .A2(net2025),
    .B1(_10289_),
    .Y(_10290_));
 sky130_fd_sc_hd__nand2_1 _30838_ (.A(_10035_),
    .B(_10290_),
    .Y(_10291_));
 sky130_fd_sc_hd__o211ai_1 _30839_ (.A1(\inst$top.soc.cpu.divider.quotient[7] ),
    .A2(net725),
    .B1(net2114),
    .C1(_10291_),
    .Y(_10292_));
 sky130_fd_sc_hd__inv_2 _30840_ (.A(_10292_),
    .Y(_03741_));
 sky130_fd_sc_hd__a21oi_1 _30841_ (.A1(_10092_),
    .A2(_10006_),
    .B1(_09925_),
    .Y(_10293_));
 sky130_fd_sc_hd__o21ai_0 _30842_ (.A1(_10006_),
    .A2(_10092_),
    .B1(_10293_),
    .Y(_10294_));
 sky130_fd_sc_hd__o221ai_1 _30843_ (.A1(_10005_),
    .A2(net1105),
    .B1(net2925),
    .B2(_09579_),
    .C1(_10294_),
    .Y(_10295_));
 sky130_fd_sc_hd__a21oi_1 _30844_ (.A1(net746),
    .A2(_10006_),
    .B1(net2974),
    .Y(_10296_));
 sky130_fd_sc_hd__o21ai_0 _30845_ (.A1(_10295_),
    .A2(net610),
    .B1(_10296_),
    .Y(_10297_));
 sky130_fd_sc_hd__inv_2 _30846_ (.A(_10297_),
    .Y(_03742_));
 sky130_fd_sc_hd__xor2_1 _30847_ (.A(\inst$top.soc.cpu.divider.quotient[9] ),
    .B(_10043_),
    .X(_10298_));
 sky130_fd_sc_hd__a22oi_1 _30848_ (.A1(\inst$top.soc.cpu.divider.quotient[8] ),
    .A2(net1035),
    .B1(_10298_),
    .B2(net1100),
    .Y(_10299_));
 sky130_fd_sc_hd__o21ai_0 _30849_ (.A1(net2925),
    .A2(_09583_),
    .B1(_10299_),
    .Y(_10300_));
 sky130_fd_sc_hd__a21oi_1 _30850_ (.A1(net746),
    .A2(_10007_),
    .B1(net2974),
    .Y(_10301_));
 sky130_fd_sc_hd__o21ai_0 _30851_ (.A1(_10300_),
    .A2(net609),
    .B1(_10301_),
    .Y(_10302_));
 sky130_fd_sc_hd__inv_2 _30852_ (.A(_10302_),
    .Y(_03743_));
 sky130_fd_sc_hd__inv_2 _30853_ (.A(_09929_),
    .Y(_10303_));
 sky130_fd_sc_hd__nand2_1 _30855_ (.A(net606),
    .B(_03082_),
    .Y(_10305_));
 sky130_fd_sc_hd__or2_2 _30856_ (.A(_02852_),
    .B(_09995_),
    .X(_10306_));
 sky130_fd_sc_hd__nor2_1 _30857_ (.A(net1105),
    .B(net856),
    .Y(_10307_));
 sky130_fd_sc_hd__nand2_1 _30859_ (.A(net836),
    .B(\inst$top.soc.cpu.divider.quotient[31] ),
    .Y(_10309_));
 sky130_fd_sc_hd__nand4_1 _30860_ (.A(_10305_),
    .B(_10306_),
    .C(_09928_),
    .D(_10309_),
    .Y(_10310_));
 sky130_fd_sc_hd__a21oi_1 _30861_ (.A1(_09997_),
    .A2(_02853_),
    .B1(net2977),
    .Y(_10311_));
 sky130_fd_sc_hd__nand2_1 _30862_ (.A(_10310_),
    .B(_10311_),
    .Y(_10312_));
 sky130_fd_sc_hd__inv_2 _30863_ (.A(_10312_),
    .Y(_03744_));
 sky130_fd_sc_hd__a31oi_1 _30866_ (.A1(_09940_),
    .A2(_02819_),
    .A3(_02822_),
    .B1(_09964_),
    .Y(_10315_));
 sky130_fd_sc_hd__xnor2_1 _30867_ (.A(_02816_),
    .B(_10315_),
    .Y(_10316_));
 sky130_fd_sc_hd__nand3_1 _30868_ (.A(net854),
    .B(net1032),
    .C(_10316_),
    .Y(_10317_));
 sky130_fd_sc_hd__xor2_1 _30869_ (.A(\inst$top.soc.cpu.divider.remainder[31] ),
    .B(_09991_),
    .X(_10318_));
 sky130_fd_sc_hd__nand3_1 _30872_ (.A(net852),
    .B(\inst$top.soc.cpu.divider.remainder[9] ),
    .C(net1032),
    .Y(_10321_));
 sky130_fd_sc_hd__inv_1 _30873_ (.A(\inst$top.soc.cpu.divider.remainder[6] ),
    .Y(_10322_));
 sky130_fd_sc_hd__inv_1 _30874_ (.A(\inst$top.soc.cpu.divider.remainder[7] ),
    .Y(_10323_));
 sky130_fd_sc_hd__inv_1 _30875_ (.A(\inst$top.soc.cpu.divider.remainder[8] ),
    .Y(_10324_));
 sky130_fd_sc_hd__inv_1 _30876_ (.A(\inst$top.soc.cpu.divider.remainder[9] ),
    .Y(_10325_));
 sky130_fd_sc_hd__nand4_1 _30877_ (.A(_10322_),
    .B(_10323_),
    .C(_10324_),
    .D(_10325_),
    .Y(_10326_));
 sky130_fd_sc_hd__nor2_1 _30878_ (.A(\inst$top.soc.cpu.divider.remainder[4] ),
    .B(\inst$top.soc.cpu.divider.remainder[5] ),
    .Y(_10327_));
 sky130_fd_sc_hd__inv_1 _30879_ (.A(\inst$top.soc.cpu.divider.remainder[2] ),
    .Y(_10328_));
 sky130_fd_sc_hd__inv_1 _30880_ (.A(\inst$top.soc.cpu.divider.remainder[3] ),
    .Y(_10329_));
 sky130_fd_sc_hd__nand4_1 _30881_ (.A(_10327_),
    .B(_10328_),
    .C(_10329_),
    .D(_02855_),
    .Y(_10330_));
 sky130_fd_sc_hd__nor2_1 _30882_ (.A(_10326_),
    .B(_10330_),
    .Y(_10331_));
 sky130_fd_sc_hd__nor2_1 _30883_ (.A(\inst$top.soc.cpu.divider.remainder[10] ),
    .B(_10331_),
    .Y(_10332_));
 sky130_fd_sc_hd__inv_1 _30884_ (.A(\inst$top.soc.cpu.divider.remainder[10] ),
    .Y(_10333_));
 sky130_fd_sc_hd__nor3_1 _30885_ (.A(_10333_),
    .B(_10326_),
    .C(_10330_),
    .Y(_10334_));
 sky130_fd_sc_hd__o21ai_0 _30887_ (.A1(_10332_),
    .A2(_10334_),
    .B1(net1665),
    .Y(_10336_));
 sky130_fd_sc_hd__nand3_1 _30888_ (.A(_10317_),
    .B(_10321_),
    .C(_10336_),
    .Y(_10337_));
 sky130_fd_sc_hd__nand2_1 _30890_ (.A(_10337_),
    .B(net2926),
    .Y(_10339_));
 sky130_fd_sc_hd__nand2_1 _30891_ (.A(net606),
    .B(net1331),
    .Y(_10340_));
 sky130_fd_sc_hd__nand3_1 _30892_ (.A(_10339_),
    .B(_10340_),
    .C(net724),
    .Y(_10341_));
 sky130_fd_sc_hd__a21oi_1 _30893_ (.A1(net745),
    .A2(_10333_),
    .B1(net2974),
    .Y(_10342_));
 sky130_fd_sc_hd__nand2_1 _30894_ (.A(_10341_),
    .B(_10342_),
    .Y(_10343_));
 sky130_fd_sc_hd__inv_2 _30895_ (.A(_10343_),
    .Y(_03745_));
 sky130_fd_sc_hd__nand2_1 _30896_ (.A(net835),
    .B(\inst$top.soc.cpu.divider.remainder[10] ),
    .Y(_10344_));
 sky130_fd_sc_hd__inv_1 _30898_ (.A(_02822_),
    .Y(_10346_));
 sky130_fd_sc_hd__nand2_1 _30899_ (.A(_02828_),
    .B(_02831_),
    .Y(_10347_));
 sky130_fd_sc_hd__a21oi_1 _30900_ (.A1(_02834_),
    .A2(_02836_),
    .B1(_02833_),
    .Y(_10348_));
 sky130_fd_sc_hd__a21oi_1 _30901_ (.A1(_02828_),
    .A2(_02830_),
    .B1(_02827_),
    .Y(_10349_));
 sky130_fd_sc_hd__o21a_1 _30902_ (.A1(_10347_),
    .A2(_10348_),
    .B1(_10349_),
    .X(_10350_));
 sky130_fd_sc_hd__inv_1 _30903_ (.A(_02834_),
    .Y(_10351_));
 sky130_fd_sc_hd__inv_1 _30904_ (.A(_02837_),
    .Y(_10352_));
 sky130_fd_sc_hd__nor3_1 _30905_ (.A(_10351_),
    .B(_10352_),
    .C(_10347_),
    .Y(_10353_));
 sky130_fd_sc_hd__a21oi_1 _30906_ (.A1(_02840_),
    .A2(_02841_),
    .B1(_02839_),
    .Y(_10354_));
 sky130_fd_sc_hd__nand3_1 _30907_ (.A(_02542_),
    .B(_02840_),
    .C(_02842_),
    .Y(_10355_));
 sky130_fd_sc_hd__nand2_1 _30908_ (.A(_10354_),
    .B(_10355_),
    .Y(_10356_));
 sky130_fd_sc_hd__nand2_1 _30909_ (.A(_10353_),
    .B(_10356_),
    .Y(_10357_));
 sky130_fd_sc_hd__nand2_1 _30910_ (.A(_10350_),
    .B(_10357_),
    .Y(_10358_));
 sky130_fd_sc_hd__a21oi_1 _30911_ (.A1(_10358_),
    .A2(_02825_),
    .B1(_02824_),
    .Y(_10359_));
 sky130_fd_sc_hd__o21bai_1 _30912_ (.A1(_10346_),
    .A2(_10359_),
    .B1_N(_02821_),
    .Y(_10360_));
 sky130_fd_sc_hd__nand2_1 _30913_ (.A(_02816_),
    .B(_02819_),
    .Y(_10361_));
 sky130_fd_sc_hd__inv_1 _30914_ (.A(_10361_),
    .Y(_10362_));
 sky130_fd_sc_hd__nand2_1 _30915_ (.A(_10360_),
    .B(_10362_),
    .Y(_10363_));
 sky130_fd_sc_hd__a21oi_1 _30916_ (.A1(_02816_),
    .A2(_02818_),
    .B1(_02815_),
    .Y(_10364_));
 sky130_fd_sc_hd__nand2_1 _30917_ (.A(_10363_),
    .B(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__xor2_1 _30918_ (.A(_02813_),
    .B(_10365_),
    .X(_10366_));
 sky130_fd_sc_hd__nand3_1 _30919_ (.A(net854),
    .B(net1032),
    .C(_10366_),
    .Y(_10367_));
 sky130_fd_sc_hd__nor3_1 _30920_ (.A(\inst$top.soc.cpu.divider.remainder[1] ),
    .B(\inst$top.soc.cpu.divider.remainder[2] ),
    .C(\inst$top.soc.cpu.divider.remainder[0] ),
    .Y(_10368_));
 sky130_fd_sc_hd__inv_1 _30921_ (.A(\inst$top.soc.cpu.divider.remainder[4] ),
    .Y(_10369_));
 sky130_fd_sc_hd__nand3_1 _30922_ (.A(_10368_),
    .B(_10329_),
    .C(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__nor3_1 _30923_ (.A(\inst$top.soc.cpu.divider.remainder[5] ),
    .B(\inst$top.soc.cpu.divider.remainder[6] ),
    .C(_10370_),
    .Y(_10371_));
 sky130_fd_sc_hd__nor2_1 _30924_ (.A(\inst$top.soc.cpu.divider.remainder[7] ),
    .B(\inst$top.soc.cpu.divider.remainder[8] ),
    .Y(_10372_));
 sky130_fd_sc_hd__nand4_1 _30925_ (.A(_10371_),
    .B(_10325_),
    .C(_10333_),
    .D(_10372_),
    .Y(_10373_));
 sky130_fd_sc_hd__inv_1 _30926_ (.A(_10373_),
    .Y(_10374_));
 sky130_fd_sc_hd__inv_1 _30927_ (.A(\inst$top.soc.cpu.divider.remainder[11] ),
    .Y(_10375_));
 sky130_fd_sc_hd__nand2_1 _30928_ (.A(_10374_),
    .B(_10375_),
    .Y(_10376_));
 sky130_fd_sc_hd__nand2_1 _30929_ (.A(_10373_),
    .B(\inst$top.soc.cpu.divider.remainder[11] ),
    .Y(_10377_));
 sky130_fd_sc_hd__nand3_1 _30930_ (.A(_10376_),
    .B(net1665),
    .C(_10377_),
    .Y(_10378_));
 sky130_fd_sc_hd__nand3_1 _30931_ (.A(_10344_),
    .B(_10367_),
    .C(_10378_),
    .Y(_10379_));
 sky130_fd_sc_hd__nand2_1 _30932_ (.A(_10379_),
    .B(net2926),
    .Y(_10380_));
 sky130_fd_sc_hd__nand2_1 _30934_ (.A(net606),
    .B(net1327),
    .Y(_10382_));
 sky130_fd_sc_hd__nand3_1 _30935_ (.A(_10380_),
    .B(net723),
    .C(_10382_),
    .Y(_10383_));
 sky130_fd_sc_hd__a21oi_1 _30937_ (.A1(net746),
    .A2(_10375_),
    .B1(net2974),
    .Y(_10385_));
 sky130_fd_sc_hd__nand2_1 _30938_ (.A(_10383_),
    .B(_10385_),
    .Y(_10386_));
 sky130_fd_sc_hd__inv_2 _30939_ (.A(_10386_),
    .Y(_03746_));
 sky130_fd_sc_hd__o21ai_0 _30940_ (.A1(_09941_),
    .A2(_10315_),
    .B1(_09966_),
    .Y(_10387_));
 sky130_fd_sc_hd__xor2_1 _30941_ (.A(_02810_),
    .B(_10387_),
    .X(_10388_));
 sky130_fd_sc_hd__nand3_1 _30942_ (.A(net854),
    .B(net1032),
    .C(_10388_),
    .Y(_10389_));
 sky130_fd_sc_hd__nand3_1 _30943_ (.A(net852),
    .B(\inst$top.soc.cpu.divider.remainder[11] ),
    .C(net1032),
    .Y(_10390_));
 sky130_fd_sc_hd__nor3_1 _30944_ (.A(\inst$top.soc.cpu.divider.remainder[6] ),
    .B(\inst$top.soc.cpu.divider.remainder[7] ),
    .C(_10330_),
    .Y(_10391_));
 sky130_fd_sc_hd__nor4_1 _30945_ (.A(\inst$top.soc.cpu.divider.remainder[8] ),
    .B(\inst$top.soc.cpu.divider.remainder[9] ),
    .C(\inst$top.soc.cpu.divider.remainder[10] ),
    .D(\inst$top.soc.cpu.divider.remainder[11] ),
    .Y(_10392_));
 sky130_fd_sc_hd__nand2_1 _30946_ (.A(_10391_),
    .B(_10392_),
    .Y(_10393_));
 sky130_fd_sc_hd__a21oi_1 _30947_ (.A1(_10393_),
    .A2(\inst$top.soc.cpu.divider.remainder[12] ),
    .B1(net1245),
    .Y(_10394_));
 sky130_fd_sc_hd__o21ai_0 _30948_ (.A1(\inst$top.soc.cpu.divider.remainder[12] ),
    .A2(_10393_),
    .B1(_10394_),
    .Y(_10395_));
 sky130_fd_sc_hd__nand3_1 _30949_ (.A(_10389_),
    .B(_10390_),
    .C(_10395_),
    .Y(_10396_));
 sky130_fd_sc_hd__nand2_1 _30950_ (.A(_10396_),
    .B(net2927),
    .Y(_10397_));
 sky130_fd_sc_hd__nand2_1 _30951_ (.A(net605),
    .B(net1322),
    .Y(_10398_));
 sky130_fd_sc_hd__nand3_1 _30952_ (.A(_10397_),
    .B(_10398_),
    .C(net723),
    .Y(_10399_));
 sky130_fd_sc_hd__inv_1 _30953_ (.A(\inst$top.soc.cpu.divider.remainder[12] ),
    .Y(_10400_));
 sky130_fd_sc_hd__a21oi_1 _30954_ (.A1(net744),
    .A2(_10400_),
    .B1(net2967),
    .Y(_10401_));
 sky130_fd_sc_hd__nand2_1 _30955_ (.A(_10399_),
    .B(_10401_),
    .Y(_10402_));
 sky130_fd_sc_hd__inv_2 _30956_ (.A(_10402_),
    .Y(_03747_));
 sky130_fd_sc_hd__nand2_1 _30957_ (.A(net835),
    .B(\inst$top.soc.cpu.divider.remainder[12] ),
    .Y(_10403_));
 sky130_fd_sc_hd__nand3_1 _30958_ (.A(_10365_),
    .B(_02810_),
    .C(_02813_),
    .Y(_10404_));
 sky130_fd_sc_hd__a21oi_1 _30959_ (.A1(_02810_),
    .A2(_02812_),
    .B1(_02809_),
    .Y(_10405_));
 sky130_fd_sc_hd__nand2_1 _30960_ (.A(_10404_),
    .B(_10405_),
    .Y(_10406_));
 sky130_fd_sc_hd__xor2_1 _30961_ (.A(_02807_),
    .B(_10406_),
    .X(_10407_));
 sky130_fd_sc_hd__nand3_1 _30962_ (.A(net854),
    .B(net1033),
    .C(_10407_),
    .Y(_10408_));
 sky130_fd_sc_hd__o21ai_0 _30963_ (.A1(\inst$top.soc.cpu.divider.remainder[12] ),
    .A2(_10376_),
    .B1(\inst$top.soc.cpu.divider.remainder[13] ),
    .Y(_10409_));
 sky130_fd_sc_hd__nor2_1 _30964_ (.A(\inst$top.soc.cpu.divider.remainder[12] ),
    .B(_10376_),
    .Y(_10410_));
 sky130_fd_sc_hd__inv_1 _30965_ (.A(\inst$top.soc.cpu.divider.remainder[13] ),
    .Y(_10411_));
 sky130_fd_sc_hd__nand2_1 _30966_ (.A(_10410_),
    .B(_10411_),
    .Y(_10412_));
 sky130_fd_sc_hd__nand3_1 _30967_ (.A(_10409_),
    .B(_10412_),
    .C(net1665),
    .Y(_10413_));
 sky130_fd_sc_hd__nand3_1 _30968_ (.A(_10403_),
    .B(_10408_),
    .C(_10413_),
    .Y(_10414_));
 sky130_fd_sc_hd__nand2_1 _30969_ (.A(_10414_),
    .B(net2926),
    .Y(_10415_));
 sky130_fd_sc_hd__nand2_1 _30970_ (.A(net605),
    .B(net1317),
    .Y(_10416_));
 sky130_fd_sc_hd__nand3_1 _30971_ (.A(_10415_),
    .B(net723),
    .C(_10416_),
    .Y(_10417_));
 sky130_fd_sc_hd__a21oi_1 _30973_ (.A1(net745),
    .A2(_10411_),
    .B1(net2975),
    .Y(_10419_));
 sky130_fd_sc_hd__nand2_1 _30974_ (.A(_10417_),
    .B(_10419_),
    .Y(_10420_));
 sky130_fd_sc_hd__inv_2 _30975_ (.A(_10420_),
    .Y(_03748_));
 sky130_fd_sc_hd__inv_1 _30976_ (.A(_09938_),
    .Y(_10421_));
 sky130_fd_sc_hd__nand2_1 _30977_ (.A(_09946_),
    .B(_09965_),
    .Y(_10422_));
 sky130_fd_sc_hd__nor3_1 _30978_ (.A(_09931_),
    .B(_09942_),
    .C(_10422_),
    .Y(_10423_));
 sky130_fd_sc_hd__nor2_1 _30979_ (.A(_09942_),
    .B(_09939_),
    .Y(_10424_));
 sky130_fd_sc_hd__nor2_1 _30980_ (.A(_09964_),
    .B(_10424_),
    .Y(_10425_));
 sky130_fd_sc_hd__a21oi_1 _30981_ (.A1(_09967_),
    .A2(_09946_),
    .B1(_09972_),
    .Y(_10426_));
 sky130_fd_sc_hd__o21ai_0 _30982_ (.A1(_10422_),
    .A2(_10425_),
    .B1(_10426_),
    .Y(_10427_));
 sky130_fd_sc_hd__a21oi_1 _30983_ (.A1(_10421_),
    .A2(_10423_),
    .B1(_10427_),
    .Y(_10428_));
 sky130_fd_sc_hd__xnor2_1 _30984_ (.A(_02804_),
    .B(_10428_),
    .Y(_10429_));
 sky130_fd_sc_hd__nand3_1 _30985_ (.A(net854),
    .B(net1033),
    .C(_10429_),
    .Y(_10430_));
 sky130_fd_sc_hd__nand3_1 _30986_ (.A(net852),
    .B(\inst$top.soc.cpu.divider.remainder[13] ),
    .C(net1035),
    .Y(_10431_));
 sky130_fd_sc_hd__nor4_1 _30987_ (.A(\inst$top.soc.cpu.divider.remainder[10] ),
    .B(\inst$top.soc.cpu.divider.remainder[11] ),
    .C(\inst$top.soc.cpu.divider.remainder[12] ),
    .D(\inst$top.soc.cpu.divider.remainder[13] ),
    .Y(_10432_));
 sky130_fd_sc_hd__nand2_1 _30988_ (.A(_10432_),
    .B(_10331_),
    .Y(_10433_));
 sky130_fd_sc_hd__a21oi_1 _30989_ (.A1(_10433_),
    .A2(\inst$top.soc.cpu.divider.remainder[14] ),
    .B1(net1245),
    .Y(_10434_));
 sky130_fd_sc_hd__o21ai_0 _30990_ (.A1(\inst$top.soc.cpu.divider.remainder[14] ),
    .A2(_10433_),
    .B1(_10434_),
    .Y(_10435_));
 sky130_fd_sc_hd__nand3_1 _30991_ (.A(_10430_),
    .B(_10431_),
    .C(_10435_),
    .Y(_10436_));
 sky130_fd_sc_hd__nand2_1 _30992_ (.A(_10436_),
    .B(net2925),
    .Y(_10437_));
 sky130_fd_sc_hd__nand2_1 _30993_ (.A(net605),
    .B(net1312),
    .Y(_10438_));
 sky130_fd_sc_hd__nand3_1 _30994_ (.A(_10437_),
    .B(_10438_),
    .C(net724),
    .Y(_10439_));
 sky130_fd_sc_hd__inv_1 _30995_ (.A(\inst$top.soc.cpu.divider.remainder[14] ),
    .Y(_10440_));
 sky130_fd_sc_hd__a21oi_1 _30996_ (.A1(net745),
    .A2(_10440_),
    .B1(net2975),
    .Y(_10441_));
 sky130_fd_sc_hd__nand2_1 _30997_ (.A(_10439_),
    .B(_10441_),
    .Y(_10442_));
 sky130_fd_sc_hd__inv_2 _30998_ (.A(_10442_),
    .Y(_03749_));
 sky130_fd_sc_hd__nand2_1 _30999_ (.A(net835),
    .B(\inst$top.soc.cpu.divider.remainder[14] ),
    .Y(_10443_));
 sky130_fd_sc_hd__inv_1 _31000_ (.A(_02825_),
    .Y(_10444_));
 sky130_fd_sc_hd__nor3_1 _31001_ (.A(_10346_),
    .B(_10444_),
    .C(_10361_),
    .Y(_10445_));
 sky130_fd_sc_hd__nand2_1 _31002_ (.A(_02810_),
    .B(_02813_),
    .Y(_10446_));
 sky130_fd_sc_hd__nand2_1 _31003_ (.A(_02804_),
    .B(_02807_),
    .Y(_10447_));
 sky130_fd_sc_hd__nor2_1 _31004_ (.A(_10446_),
    .B(_10447_),
    .Y(_10448_));
 sky130_fd_sc_hd__nand3_1 _31005_ (.A(_10358_),
    .B(_10445_),
    .C(_10448_),
    .Y(_10449_));
 sky130_fd_sc_hd__a21oi_1 _31006_ (.A1(_02822_),
    .A2(_02824_),
    .B1(_02821_),
    .Y(_10450_));
 sky130_fd_sc_hd__o21ai_0 _31007_ (.A1(_10361_),
    .A2(_10450_),
    .B1(_10364_),
    .Y(_10451_));
 sky130_fd_sc_hd__a21oi_1 _31008_ (.A1(_02804_),
    .A2(_02806_),
    .B1(_02803_),
    .Y(_10452_));
 sky130_fd_sc_hd__o21ai_0 _31009_ (.A1(_10447_),
    .A2(_10405_),
    .B1(_10452_),
    .Y(_10453_));
 sky130_fd_sc_hd__a21oi_1 _31010_ (.A1(_10451_),
    .A2(_10448_),
    .B1(_10453_),
    .Y(_10454_));
 sky130_fd_sc_hd__nand2_1 _31011_ (.A(_10449_),
    .B(_10454_),
    .Y(_10455_));
 sky130_fd_sc_hd__xor2_1 _31012_ (.A(_02801_),
    .B(_10455_),
    .X(_10456_));
 sky130_fd_sc_hd__nand3_1 _31013_ (.A(net854),
    .B(net1033),
    .C(_10456_),
    .Y(_10457_));
 sky130_fd_sc_hd__nand3_1 _31014_ (.A(_10410_),
    .B(_10411_),
    .C(_10440_),
    .Y(_10458_));
 sky130_fd_sc_hd__inv_1 _31015_ (.A(_10458_),
    .Y(_10459_));
 sky130_fd_sc_hd__inv_1 _31016_ (.A(\inst$top.soc.cpu.divider.remainder[15] ),
    .Y(_10460_));
 sky130_fd_sc_hd__nand2_1 _31017_ (.A(_10459_),
    .B(_10460_),
    .Y(_10461_));
 sky130_fd_sc_hd__nand2_1 _31018_ (.A(_10458_),
    .B(\inst$top.soc.cpu.divider.remainder[15] ),
    .Y(_10462_));
 sky130_fd_sc_hd__nand3_1 _31019_ (.A(_10461_),
    .B(net1665),
    .C(_10462_),
    .Y(_10463_));
 sky130_fd_sc_hd__nand3_1 _31020_ (.A(_10443_),
    .B(_10457_),
    .C(_10463_),
    .Y(_10464_));
 sky130_fd_sc_hd__nand2_1 _31021_ (.A(_10464_),
    .B(net2925),
    .Y(_10465_));
 sky130_fd_sc_hd__nand2_1 _31022_ (.A(net605),
    .B(net1308),
    .Y(_10466_));
 sky130_fd_sc_hd__nand3_1 _31023_ (.A(_10465_),
    .B(net723),
    .C(_10466_),
    .Y(_10467_));
 sky130_fd_sc_hd__a21oi_1 _31024_ (.A1(net745),
    .A2(_10460_),
    .B1(net2975),
    .Y(_10468_));
 sky130_fd_sc_hd__nand2_1 _31025_ (.A(_10467_),
    .B(_10468_),
    .Y(_10469_));
 sky130_fd_sc_hd__inv_2 _31026_ (.A(_10469_),
    .Y(_03750_));
 sky130_fd_sc_hd__a21oi_1 _31027_ (.A1(_09940_),
    .A2(_09948_),
    .B1(_09974_),
    .Y(_10470_));
 sky130_fd_sc_hd__xnor2_1 _31028_ (.A(_02798_),
    .B(_10470_),
    .Y(_10471_));
 sky130_fd_sc_hd__nand3_1 _31029_ (.A(net854),
    .B(net1033),
    .C(_10471_),
    .Y(_10472_));
 sky130_fd_sc_hd__nand3_1 _31030_ (.A(net852),
    .B(\inst$top.soc.cpu.divider.remainder[15] ),
    .C(net1033),
    .Y(_10473_));
 sky130_fd_sc_hd__nor4_1 _31031_ (.A(\inst$top.soc.cpu.divider.remainder[12] ),
    .B(\inst$top.soc.cpu.divider.remainder[13] ),
    .C(\inst$top.soc.cpu.divider.remainder[14] ),
    .D(\inst$top.soc.cpu.divider.remainder[15] ),
    .Y(_10474_));
 sky130_fd_sc_hd__inv_1 _31032_ (.A(_10474_),
    .Y(_10475_));
 sky130_fd_sc_hd__nor2_1 _31033_ (.A(_10475_),
    .B(_10393_),
    .Y(_10476_));
 sky130_fd_sc_hd__inv_1 _31034_ (.A(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__a21oi_1 _31035_ (.A1(_10477_),
    .A2(\inst$top.soc.cpu.divider.remainder[16] ),
    .B1(net1245),
    .Y(_10478_));
 sky130_fd_sc_hd__o21ai_0 _31036_ (.A1(\inst$top.soc.cpu.divider.remainder[16] ),
    .A2(_10477_),
    .B1(_10478_),
    .Y(_10479_));
 sky130_fd_sc_hd__nand3_1 _31037_ (.A(_10472_),
    .B(_10473_),
    .C(_10479_),
    .Y(_10480_));
 sky130_fd_sc_hd__nand2_1 _31038_ (.A(_10480_),
    .B(net2925),
    .Y(_10481_));
 sky130_fd_sc_hd__nand2_1 _31039_ (.A(net606),
    .B(net1303),
    .Y(_10482_));
 sky130_fd_sc_hd__nand3_1 _31040_ (.A(_10481_),
    .B(_10482_),
    .C(net724),
    .Y(_10483_));
 sky130_fd_sc_hd__inv_1 _31041_ (.A(\inst$top.soc.cpu.divider.remainder[16] ),
    .Y(_10484_));
 sky130_fd_sc_hd__a21oi_1 _31042_ (.A1(net745),
    .A2(_10484_),
    .B1(net2974),
    .Y(_10485_));
 sky130_fd_sc_hd__nand2_1 _31043_ (.A(_10483_),
    .B(_10485_),
    .Y(_10486_));
 sky130_fd_sc_hd__inv_2 _31044_ (.A(_10486_),
    .Y(_03751_));
 sky130_fd_sc_hd__nand2_1 _31045_ (.A(net835),
    .B(\inst$top.soc.cpu.divider.remainder[16] ),
    .Y(_10487_));
 sky130_fd_sc_hd__nand2_1 _31046_ (.A(_02798_),
    .B(_02801_),
    .Y(_10488_));
 sky130_fd_sc_hd__inv_1 _31047_ (.A(_10488_),
    .Y(_10489_));
 sky130_fd_sc_hd__a21oi_1 _31048_ (.A1(_02798_),
    .A2(_02800_),
    .B1(_02797_),
    .Y(_10490_));
 sky130_fd_sc_hd__inv_1 _31049_ (.A(_10490_),
    .Y(_10491_));
 sky130_fd_sc_hd__a21oi_1 _31050_ (.A1(_10455_),
    .A2(_10489_),
    .B1(_10491_),
    .Y(_10492_));
 sky130_fd_sc_hd__xnor2_1 _31051_ (.A(_02795_),
    .B(_10492_),
    .Y(_10493_));
 sky130_fd_sc_hd__nand3_1 _31052_ (.A(net855),
    .B(net1034),
    .C(_10493_),
    .Y(_10494_));
 sky130_fd_sc_hd__nand3_1 _31053_ (.A(_10459_),
    .B(_10460_),
    .C(_10484_),
    .Y(_10495_));
 sky130_fd_sc_hd__inv_1 _31054_ (.A(_10495_),
    .Y(_10496_));
 sky130_fd_sc_hd__inv_1 _31055_ (.A(\inst$top.soc.cpu.divider.remainder[17] ),
    .Y(_10497_));
 sky130_fd_sc_hd__nand2_1 _31056_ (.A(_10496_),
    .B(_10497_),
    .Y(_10498_));
 sky130_fd_sc_hd__nand2_1 _31057_ (.A(_10495_),
    .B(\inst$top.soc.cpu.divider.remainder[17] ),
    .Y(_10499_));
 sky130_fd_sc_hd__nand3_1 _31058_ (.A(_10498_),
    .B(net1665),
    .C(_10499_),
    .Y(_10500_));
 sky130_fd_sc_hd__nand3_1 _31059_ (.A(_10487_),
    .B(_10494_),
    .C(_10500_),
    .Y(_10501_));
 sky130_fd_sc_hd__nand2_1 _31061_ (.A(_10501_),
    .B(net2926),
    .Y(_10503_));
 sky130_fd_sc_hd__nand2_1 _31063_ (.A(net607),
    .B(net1299),
    .Y(_10505_));
 sky130_fd_sc_hd__nand3_1 _31064_ (.A(_10503_),
    .B(net723),
    .C(_10505_),
    .Y(_10506_));
 sky130_fd_sc_hd__a21oi_1 _31065_ (.A1(net745),
    .A2(_10497_),
    .B1(net2976),
    .Y(_10507_));
 sky130_fd_sc_hd__nand2_1 _31066_ (.A(_10506_),
    .B(_10507_),
    .Y(_10508_));
 sky130_fd_sc_hd__inv_2 _31067_ (.A(_10508_),
    .Y(_03752_));
 sky130_fd_sc_hd__o21ai_1 _31068_ (.A1(net1295),
    .A2(net749),
    .B1(net610),
    .Y(_10509_));
 sky130_fd_sc_hd__nand2_1 _31069_ (.A(net835),
    .B(\inst$top.soc.cpu.divider.remainder[17] ),
    .Y(_10510_));
 sky130_fd_sc_hd__nor2_1 _31070_ (.A(_09952_),
    .B(_10428_),
    .Y(_10511_));
 sky130_fd_sc_hd__o21ai_0 _31071_ (.A1(_09952_),
    .A2(_09969_),
    .B1(_09955_),
    .Y(_10512_));
 sky130_fd_sc_hd__a21oi_1 _31072_ (.A1(_10511_),
    .A2(_09944_),
    .B1(_10512_),
    .Y(_10513_));
 sky130_fd_sc_hd__xor2_1 _31073_ (.A(_02792_),
    .B(_10513_),
    .X(_10514_));
 sky130_fd_sc_hd__nand3b_1 _31074_ (.A_N(_10514_),
    .B(net855),
    .C(net1034),
    .Y(_10515_));
 sky130_fd_sc_hd__inv_1 _31075_ (.A(\inst$top.soc.cpu.divider.remainder[18] ),
    .Y(_10516_));
 sky130_fd_sc_hd__nand2_1 _31076_ (.A(_10484_),
    .B(_10497_),
    .Y(_10517_));
 sky130_fd_sc_hd__nor4_1 _31077_ (.A(\inst$top.soc.cpu.divider.remainder[14] ),
    .B(\inst$top.soc.cpu.divider.remainder[15] ),
    .C(_10517_),
    .D(_10433_),
    .Y(_10518_));
 sky130_fd_sc_hd__xor2_1 _31078_ (.A(_10516_),
    .B(_10518_),
    .X(_10519_));
 sky130_fd_sc_hd__nand2_1 _31079_ (.A(_10519_),
    .B(net1665),
    .Y(_10520_));
 sky130_fd_sc_hd__nand3_1 _31080_ (.A(_10510_),
    .B(_10515_),
    .C(_10520_),
    .Y(_10521_));
 sky130_fd_sc_hd__nand2_1 _31081_ (.A(_10521_),
    .B(net2928),
    .Y(_10522_));
 sky130_fd_sc_hd__o21ai_0 _31082_ (.A1(\inst$top.soc.cpu.divider.remainder[18] ),
    .A2(net725),
    .B1(net2117),
    .Y(_10523_));
 sky130_fd_sc_hd__a21oi_4 _31083_ (.A1(_10509_),
    .A2(_10522_),
    .B1(_10523_),
    .Y(_03753_));
 sky130_fd_sc_hd__nand2_1 _31084_ (.A(_02792_),
    .B(_02795_),
    .Y(_10524_));
 sky130_fd_sc_hd__a21oi_1 _31085_ (.A1(_02792_),
    .A2(_02794_),
    .B1(_02791_),
    .Y(_10525_));
 sky130_fd_sc_hd__o21ai_0 _31086_ (.A1(_10524_),
    .A2(_10492_),
    .B1(_10525_),
    .Y(_10526_));
 sky130_fd_sc_hd__xor2_1 _31087_ (.A(_02789_),
    .B(_10526_),
    .X(_10527_));
 sky130_fd_sc_hd__nand3_1 _31088_ (.A(net855),
    .B(net1034),
    .C(_10527_),
    .Y(_10528_));
 sky130_fd_sc_hd__nand3_1 _31089_ (.A(net853),
    .B(\inst$top.soc.cpu.divider.remainder[18] ),
    .C(net1040),
    .Y(_10529_));
 sky130_fd_sc_hd__inv_1 _31090_ (.A(\inst$top.soc.cpu.divider.remainder[19] ),
    .Y(_10530_));
 sky130_fd_sc_hd__nand4_1 _31091_ (.A(_10460_),
    .B(_10484_),
    .C(_10497_),
    .D(_10516_),
    .Y(_10531_));
 sky130_fd_sc_hd__nor2_1 _31092_ (.A(_10531_),
    .B(_10458_),
    .Y(_10532_));
 sky130_fd_sc_hd__xor2_1 _31093_ (.A(_10530_),
    .B(_10532_),
    .X(_10533_));
 sky130_fd_sc_hd__nand2_1 _31095_ (.A(_10533_),
    .B(net1664),
    .Y(_10535_));
 sky130_fd_sc_hd__nand3_1 _31096_ (.A(_10528_),
    .B(_10529_),
    .C(_10535_),
    .Y(_10536_));
 sky130_fd_sc_hd__nand2_1 _31097_ (.A(_10536_),
    .B(net2926),
    .Y(_10537_));
 sky130_fd_sc_hd__nand2_1 _31098_ (.A(net605),
    .B(net1289),
    .Y(_10538_));
 sky130_fd_sc_hd__nand3_1 _31099_ (.A(_10537_),
    .B(_10538_),
    .C(net724),
    .Y(_10539_));
 sky130_fd_sc_hd__a21oi_1 _31100_ (.A1(net745),
    .A2(_10530_),
    .B1(net2976),
    .Y(_10540_));
 sky130_fd_sc_hd__nand2_1 _31101_ (.A(_10539_),
    .B(_10540_),
    .Y(_10541_));
 sky130_fd_sc_hd__inv_2 _31102_ (.A(_10541_),
    .Y(_03754_));
 sky130_fd_sc_hd__nand2_1 _31103_ (.A(net606),
    .B(net1262),
    .Y(_10542_));
 sky130_fd_sc_hd__nand2_1 _31104_ (.A(net836),
    .B(\inst$top.soc.cpu.divider.remainder[0] ),
    .Y(_10543_));
 sky130_fd_sc_hd__nand3_1 _31105_ (.A(net856),
    .B(_02544_),
    .C(net1039),
    .Y(_10544_));
 sky130_fd_sc_hd__a21oi_1 _31106_ (.A1(_02856_),
    .A2(net1102),
    .B1(net749),
    .Y(_10545_));
 sky130_fd_sc_hd__nand4_1 _31107_ (.A(_10542_),
    .B(_10543_),
    .C(_10544_),
    .D(_10545_),
    .Y(_10546_));
 sky130_fd_sc_hd__a21oi_1 _31108_ (.A1(net749),
    .A2(_02854_),
    .B1(net2975),
    .Y(_10547_));
 sky130_fd_sc_hd__nand2_1 _31109_ (.A(_10546_),
    .B(_10547_),
    .Y(_10548_));
 sky130_fd_sc_hd__inv_2 _31110_ (.A(_10548_),
    .Y(_03755_));
 sky130_fd_sc_hd__o21ai_0 _31112_ (.A1(_09951_),
    .A2(_10513_),
    .B1(_09956_),
    .Y(_10550_));
 sky130_fd_sc_hd__xor2_1 _31113_ (.A(_02786_),
    .B(_10550_),
    .X(_10551_));
 sky130_fd_sc_hd__nand3_1 _31114_ (.A(net855),
    .B(_10551_),
    .C(net1034),
    .Y(_10552_));
 sky130_fd_sc_hd__nand3_1 _31115_ (.A(net853),
    .B(\inst$top.soc.cpu.divider.remainder[19] ),
    .C(net1034),
    .Y(_10553_));
 sky130_fd_sc_hd__nor3_1 _31116_ (.A(\inst$top.soc.cpu.divider.remainder[18] ),
    .B(\inst$top.soc.cpu.divider.remainder[19] ),
    .C(_10517_),
    .Y(_10554_));
 sky130_fd_sc_hd__nand2_1 _31117_ (.A(_10476_),
    .B(_10554_),
    .Y(_10555_));
 sky130_fd_sc_hd__xor2_1 _31118_ (.A(\inst$top.soc.cpu.divider.remainder[20] ),
    .B(_10555_),
    .X(_10556_));
 sky130_fd_sc_hd__nand2_1 _31119_ (.A(_10556_),
    .B(net1665),
    .Y(_10557_));
 sky130_fd_sc_hd__nand3_1 _31120_ (.A(_10552_),
    .B(_10553_),
    .C(_10557_),
    .Y(_10558_));
 sky130_fd_sc_hd__nand2_1 _31121_ (.A(_10558_),
    .B(net2926),
    .Y(_10559_));
 sky130_fd_sc_hd__nand2_1 _31122_ (.A(net605),
    .B(net1286),
    .Y(_10560_));
 sky130_fd_sc_hd__nand3_1 _31123_ (.A(_10559_),
    .B(_10560_),
    .C(net725),
    .Y(_10561_));
 sky130_fd_sc_hd__inv_1 _31124_ (.A(\inst$top.soc.cpu.divider.remainder[20] ),
    .Y(_10562_));
 sky130_fd_sc_hd__a21oi_1 _31125_ (.A1(net751),
    .A2(_10562_),
    .B1(net2976),
    .Y(_10563_));
 sky130_fd_sc_hd__nand2_1 _31126_ (.A(_10561_),
    .B(_10563_),
    .Y(_10564_));
 sky130_fd_sc_hd__inv_2 _31127_ (.A(_10564_),
    .Y(_03756_));
 sky130_fd_sc_hd__nand2_1 _31128_ (.A(net606),
    .B(net1281),
    .Y(_10565_));
 sky130_fd_sc_hd__nor4_1 _31129_ (.A(\inst$top.soc.cpu.divider.remainder[17] ),
    .B(\inst$top.soc.cpu.divider.remainder[18] ),
    .C(\inst$top.soc.cpu.divider.remainder[19] ),
    .D(\inst$top.soc.cpu.divider.remainder[20] ),
    .Y(_10566_));
 sky130_fd_sc_hd__inv_1 _31130_ (.A(_10566_),
    .Y(_10567_));
 sky130_fd_sc_hd__o21ai_0 _31131_ (.A1(_10567_),
    .A2(_10495_),
    .B1(\inst$top.soc.cpu.divider.remainder[21] ),
    .Y(_10568_));
 sky130_fd_sc_hd__inv_1 _31132_ (.A(\inst$top.soc.cpu.divider.remainder[21] ),
    .Y(_10569_));
 sky130_fd_sc_hd__nand3_1 _31133_ (.A(_10496_),
    .B(_10569_),
    .C(_10566_),
    .Y(_10570_));
 sky130_fd_sc_hd__a31oi_1 _31134_ (.A1(_10568_),
    .A2(_10570_),
    .A3(net1103),
    .B1(net745),
    .Y(_10571_));
 sky130_fd_sc_hd__nand2_1 _31135_ (.A(_02786_),
    .B(_02789_),
    .Y(_10572_));
 sky130_fd_sc_hd__inv_1 _31136_ (.A(_10572_),
    .Y(_10573_));
 sky130_fd_sc_hd__a21oi_1 _31137_ (.A1(_02786_),
    .A2(_02788_),
    .B1(_02785_),
    .Y(_10574_));
 sky130_fd_sc_hd__a21boi_0 _31138_ (.A1(_10526_),
    .A2(_10573_),
    .B1_N(_10574_),
    .Y(_10575_));
 sky130_fd_sc_hd__xnor2_1 _31139_ (.A(_02783_),
    .B(_10575_),
    .Y(_10576_));
 sky130_fd_sc_hd__nand3_1 _31140_ (.A(net855),
    .B(net1034),
    .C(_10576_),
    .Y(_10577_));
 sky130_fd_sc_hd__nand2_1 _31141_ (.A(net835),
    .B(\inst$top.soc.cpu.divider.remainder[20] ),
    .Y(_10578_));
 sky130_fd_sc_hd__nand4_1 _31142_ (.A(_10565_),
    .B(_10571_),
    .C(_10577_),
    .D(_10578_),
    .Y(_10579_));
 sky130_fd_sc_hd__a21oi_1 _31144_ (.A1(net746),
    .A2(_10569_),
    .B1(net2974),
    .Y(_10581_));
 sky130_fd_sc_hd__nand2_1 _31145_ (.A(_10579_),
    .B(_10581_),
    .Y(_10582_));
 sky130_fd_sc_hd__inv_2 _31146_ (.A(_10582_),
    .Y(_03757_));
 sky130_fd_sc_hd__nor4_1 _31147_ (.A(_09950_),
    .B(_09951_),
    .C(_09943_),
    .D(_09952_),
    .Y(_10583_));
 sky130_fd_sc_hd__nand3_1 _31148_ (.A(_10421_),
    .B(_10423_),
    .C(_10583_),
    .Y(_10584_));
 sky130_fd_sc_hd__nor2_1 _31149_ (.A(_09950_),
    .B(_09951_),
    .Y(_10585_));
 sky130_fd_sc_hd__o21ai_0 _31150_ (.A1(_09950_),
    .A2(_09956_),
    .B1(_09959_),
    .Y(_10586_));
 sky130_fd_sc_hd__a21oi_1 _31151_ (.A1(_10512_),
    .A2(_10585_),
    .B1(_10586_),
    .Y(_10587_));
 sky130_fd_sc_hd__nand2_1 _31152_ (.A(_10427_),
    .B(_10583_),
    .Y(_10588_));
 sky130_fd_sc_hd__nand3_1 _31153_ (.A(_10584_),
    .B(_10587_),
    .C(_10588_),
    .Y(_10589_));
 sky130_fd_sc_hd__xor2_1 _31154_ (.A(_02780_),
    .B(_10589_),
    .X(_10590_));
 sky130_fd_sc_hd__nand3_1 _31155_ (.A(net856),
    .B(net1038),
    .C(_10590_),
    .Y(_10591_));
 sky130_fd_sc_hd__nand3_1 _31156_ (.A(net853),
    .B(\inst$top.soc.cpu.divider.remainder[21] ),
    .C(net1038),
    .Y(_10592_));
 sky130_fd_sc_hd__nor2_1 _31157_ (.A(\inst$top.soc.cpu.divider.remainder[20] ),
    .B(\inst$top.soc.cpu.divider.remainder[21] ),
    .Y(_10593_));
 sky130_fd_sc_hd__nand4_1 _31158_ (.A(_10518_),
    .B(_10516_),
    .C(_10530_),
    .D(_10593_),
    .Y(_10594_));
 sky130_fd_sc_hd__xor2_1 _31159_ (.A(\inst$top.soc.cpu.divider.remainder[22] ),
    .B(_10594_),
    .X(_10595_));
 sky130_fd_sc_hd__nand2_1 _31160_ (.A(_10595_),
    .B(net1664),
    .Y(_10596_));
 sky130_fd_sc_hd__nand3_1 _31161_ (.A(_10591_),
    .B(_10592_),
    .C(_10596_),
    .Y(_10597_));
 sky130_fd_sc_hd__nand2_1 _31162_ (.A(_10597_),
    .B(net2928),
    .Y(_10598_));
 sky130_fd_sc_hd__nand2_1 _31163_ (.A(net608),
    .B(net1260),
    .Y(_10599_));
 sky130_fd_sc_hd__nand3_1 _31164_ (.A(_10598_),
    .B(_10599_),
    .C(net725),
    .Y(_10600_));
 sky130_fd_sc_hd__inv_1 _31165_ (.A(\inst$top.soc.cpu.divider.remainder[22] ),
    .Y(_10601_));
 sky130_fd_sc_hd__a21oi_1 _31166_ (.A1(net751),
    .A2(_10601_),
    .B1(net2975),
    .Y(_10602_));
 sky130_fd_sc_hd__nand2_1 _31167_ (.A(_10600_),
    .B(_10602_),
    .Y(_10603_));
 sky130_fd_sc_hd__inv_2 _31168_ (.A(_10603_),
    .Y(_03758_));
 sky130_fd_sc_hd__nand2_1 _31169_ (.A(net836),
    .B(\inst$top.soc.cpu.divider.remainder[22] ),
    .Y(_10604_));
 sky130_fd_sc_hd__nand2_1 _31170_ (.A(_02780_),
    .B(_02783_),
    .Y(_10605_));
 sky130_fd_sc_hd__nor2_1 _31171_ (.A(_10572_),
    .B(_10605_),
    .Y(_10606_));
 sky130_fd_sc_hd__a21oi_1 _31172_ (.A1(_02780_),
    .A2(_02782_),
    .B1(_02779_),
    .Y(_10607_));
 sky130_fd_sc_hd__o21ai_0 _31173_ (.A1(_10605_),
    .A2(_10574_),
    .B1(_10607_),
    .Y(_10608_));
 sky130_fd_sc_hd__a21oi_1 _31174_ (.A1(_10526_),
    .A2(_10606_),
    .B1(_10608_),
    .Y(_10609_));
 sky130_fd_sc_hd__xnor2_1 _31175_ (.A(_02777_),
    .B(_10609_),
    .Y(_10610_));
 sky130_fd_sc_hd__nand3_1 _31176_ (.A(net856),
    .B(_10610_),
    .C(net1038),
    .Y(_10611_));
 sky130_fd_sc_hd__nor2_1 _31177_ (.A(\inst$top.soc.cpu.divider.remainder[21] ),
    .B(\inst$top.soc.cpu.divider.remainder[22] ),
    .Y(_10612_));
 sky130_fd_sc_hd__nand3_1 _31178_ (.A(_10612_),
    .B(_10530_),
    .C(_10562_),
    .Y(_10613_));
 sky130_fd_sc_hd__inv_1 _31179_ (.A(_10613_),
    .Y(_10614_));
 sky130_fd_sc_hd__nand2_1 _31180_ (.A(_10532_),
    .B(_10614_),
    .Y(_10615_));
 sky130_fd_sc_hd__a21oi_1 _31181_ (.A1(_10615_),
    .A2(\inst$top.soc.cpu.divider.remainder[23] ),
    .B1(_09907_),
    .Y(_10616_));
 sky130_fd_sc_hd__o21ai_0 _31182_ (.A1(\inst$top.soc.cpu.divider.remainder[23] ),
    .A2(_10615_),
    .B1(_10616_),
    .Y(_10617_));
 sky130_fd_sc_hd__nand3_1 _31183_ (.A(_10604_),
    .B(_10611_),
    .C(_10617_),
    .Y(_10618_));
 sky130_fd_sc_hd__nand2_1 _31184_ (.A(_10618_),
    .B(net2928),
    .Y(_10619_));
 sky130_fd_sc_hd__nand2_1 _31185_ (.A(net607),
    .B(net1276),
    .Y(_10620_));
 sky130_fd_sc_hd__nand3_1 _31186_ (.A(_10619_),
    .B(net725),
    .C(_10620_),
    .Y(_10621_));
 sky130_fd_sc_hd__inv_1 _31187_ (.A(\inst$top.soc.cpu.divider.remainder[23] ),
    .Y(_10622_));
 sky130_fd_sc_hd__a21oi_1 _31189_ (.A1(net751),
    .A2(_10622_),
    .B1(net2976),
    .Y(_10624_));
 sky130_fd_sc_hd__nand2_1 _31190_ (.A(_10621_),
    .B(_10624_),
    .Y(_10625_));
 sky130_fd_sc_hd__inv_2 _31191_ (.A(_10625_),
    .Y(_03759_));
 sky130_fd_sc_hd__xor2_1 _31192_ (.A(_02774_),
    .B(_09976_),
    .X(_10626_));
 sky130_fd_sc_hd__nand3_1 _31193_ (.A(net856),
    .B(net1038),
    .C(_10626_),
    .Y(_10627_));
 sky130_fd_sc_hd__nand3_1 _31194_ (.A(net853),
    .B(\inst$top.soc.cpu.divider.remainder[23] ),
    .C(net1038),
    .Y(_10628_));
 sky130_fd_sc_hd__nand3_1 _31195_ (.A(_10593_),
    .B(_10601_),
    .C(_10622_),
    .Y(_10629_));
 sky130_fd_sc_hd__nor2_1 _31196_ (.A(_10629_),
    .B(_10555_),
    .Y(_10630_));
 sky130_fd_sc_hd__inv_1 _31197_ (.A(_10630_),
    .Y(_10631_));
 sky130_fd_sc_hd__a21oi_1 _31198_ (.A1(_10631_),
    .A2(\inst$top.soc.cpu.divider.remainder[24] ),
    .B1(net1245),
    .Y(_10632_));
 sky130_fd_sc_hd__o21ai_0 _31199_ (.A1(\inst$top.soc.cpu.divider.remainder[24] ),
    .A2(_10631_),
    .B1(_10632_),
    .Y(_10633_));
 sky130_fd_sc_hd__nand3_1 _31200_ (.A(_10627_),
    .B(_10628_),
    .C(_10633_),
    .Y(_10634_));
 sky130_fd_sc_hd__nand2_1 _31201_ (.A(_10634_),
    .B(net2928),
    .Y(_10635_));
 sky130_fd_sc_hd__nand2_1 _31202_ (.A(net607),
    .B(net1272),
    .Y(_10636_));
 sky130_fd_sc_hd__nand3_1 _31203_ (.A(_10635_),
    .B(_10636_),
    .C(net726),
    .Y(_10637_));
 sky130_fd_sc_hd__inv_1 _31204_ (.A(\inst$top.soc.cpu.divider.remainder[24] ),
    .Y(_10638_));
 sky130_fd_sc_hd__a21oi_1 _31205_ (.A1(net750),
    .A2(_10638_),
    .B1(net2976),
    .Y(_10639_));
 sky130_fd_sc_hd__nand2_1 _31206_ (.A(_10637_),
    .B(_10639_),
    .Y(_10640_));
 sky130_fd_sc_hd__inv_2 _31207_ (.A(_10640_),
    .Y(_03760_));
 sky130_fd_sc_hd__a21oi_1 _31208_ (.A1(net607),
    .A2(net1256),
    .B1(net749),
    .Y(_10641_));
 sky130_fd_sc_hd__nand2_1 _31209_ (.A(_02774_),
    .B(_02777_),
    .Y(_10642_));
 sky130_fd_sc_hd__a21oi_1 _31210_ (.A1(_02774_),
    .A2(_02776_),
    .B1(_02773_),
    .Y(_10643_));
 sky130_fd_sc_hd__o21ai_0 _31211_ (.A1(_10642_),
    .A2(_10609_),
    .B1(_10643_),
    .Y(_10644_));
 sky130_fd_sc_hd__xor2_1 _31212_ (.A(_02771_),
    .B(_10644_),
    .X(_10645_));
 sky130_fd_sc_hd__nand3_1 _31213_ (.A(_10645_),
    .B(net856),
    .C(net1038),
    .Y(_10646_));
 sky130_fd_sc_hd__nand3_1 _31214_ (.A(net853),
    .B(\inst$top.soc.cpu.divider.remainder[24] ),
    .C(net1038),
    .Y(_10647_));
 sky130_fd_sc_hd__nor2_1 _31215_ (.A(\inst$top.soc.cpu.divider.remainder[23] ),
    .B(_10615_),
    .Y(_10648_));
 sky130_fd_sc_hd__nand2_1 _31216_ (.A(_10648_),
    .B(_10638_),
    .Y(_10649_));
 sky130_fd_sc_hd__a21oi_1 _31217_ (.A1(_10649_),
    .A2(\inst$top.soc.cpu.divider.remainder[25] ),
    .B1(net1245),
    .Y(_10650_));
 sky130_fd_sc_hd__o21ai_0 _31218_ (.A1(\inst$top.soc.cpu.divider.remainder[25] ),
    .A2(_10649_),
    .B1(_10650_),
    .Y(_10651_));
 sky130_fd_sc_hd__nand3_1 _31219_ (.A(_10646_),
    .B(_10647_),
    .C(_10651_),
    .Y(_10652_));
 sky130_fd_sc_hd__nand2_1 _31220_ (.A(_10652_),
    .B(net2929),
    .Y(_10653_));
 sky130_fd_sc_hd__nand2_1 _31221_ (.A(_10641_),
    .B(_10653_),
    .Y(_10654_));
 sky130_fd_sc_hd__inv_1 _31222_ (.A(\inst$top.soc.cpu.divider.remainder[25] ),
    .Y(_10655_));
 sky130_fd_sc_hd__a21oi_1 _31223_ (.A1(net750),
    .A2(_10655_),
    .B1(net2978),
    .Y(_10656_));
 sky130_fd_sc_hd__nand2_1 _31224_ (.A(_10654_),
    .B(_10656_),
    .Y(_10657_));
 sky130_fd_sc_hd__inv_2 _31225_ (.A(_10657_),
    .Y(_03761_));
 sky130_fd_sc_hd__nor2_1 _31226_ (.A(_09978_),
    .B(_09949_),
    .Y(_10658_));
 sky130_fd_sc_hd__nand2_1 _31227_ (.A(_10589_),
    .B(_10658_),
    .Y(_10659_));
 sky130_fd_sc_hd__o211ai_1 _31228_ (.A1(_09978_),
    .A2(_09960_),
    .B1(_09980_),
    .C1(_10659_),
    .Y(_10660_));
 sky130_fd_sc_hd__xor2_1 _31229_ (.A(_02768_),
    .B(_10660_),
    .X(_10661_));
 sky130_fd_sc_hd__nand3_1 _31230_ (.A(net857),
    .B(net1039),
    .C(_10661_),
    .Y(_10662_));
 sky130_fd_sc_hd__nand3_1 _31231_ (.A(net852),
    .B(\inst$top.soc.cpu.divider.remainder[25] ),
    .C(net1039),
    .Y(_10663_));
 sky130_fd_sc_hd__nor4_1 _31232_ (.A(\inst$top.soc.cpu.divider.remainder[22] ),
    .B(\inst$top.soc.cpu.divider.remainder[23] ),
    .C(\inst$top.soc.cpu.divider.remainder[24] ),
    .D(\inst$top.soc.cpu.divider.remainder[25] ),
    .Y(_10664_));
 sky130_fd_sc_hd__inv_1 _31233_ (.A(_10664_),
    .Y(_10665_));
 sky130_fd_sc_hd__o21ai_0 _31234_ (.A1(_10665_),
    .A2(_10594_),
    .B1(\inst$top.soc.cpu.divider.remainder[26] ),
    .Y(_10666_));
 sky130_fd_sc_hd__nor2_1 _31235_ (.A(_10665_),
    .B(_10594_),
    .Y(_10667_));
 sky130_fd_sc_hd__inv_1 _31236_ (.A(\inst$top.soc.cpu.divider.remainder[26] ),
    .Y(_10668_));
 sky130_fd_sc_hd__nand2_1 _31237_ (.A(_10667_),
    .B(_10668_),
    .Y(_10669_));
 sky130_fd_sc_hd__nand3_1 _31238_ (.A(_10666_),
    .B(_10669_),
    .C(net1664),
    .Y(_10670_));
 sky130_fd_sc_hd__nand3_1 _31239_ (.A(_10662_),
    .B(_10663_),
    .C(_10670_),
    .Y(_10671_));
 sky130_fd_sc_hd__nand2_1 _31240_ (.A(_10671_),
    .B(net2929),
    .Y(_10672_));
 sky130_fd_sc_hd__nand2_1 _31241_ (.A(net606),
    .B(net1253),
    .Y(_10673_));
 sky130_fd_sc_hd__nand3_1 _31242_ (.A(_10672_),
    .B(_10673_),
    .C(net726),
    .Y(_10674_));
 sky130_fd_sc_hd__a21oi_1 _31243_ (.A1(net750),
    .A2(_10668_),
    .B1(net2977),
    .Y(_10675_));
 sky130_fd_sc_hd__nand2_1 _31244_ (.A(_10674_),
    .B(_10675_),
    .Y(_10676_));
 sky130_fd_sc_hd__inv_2 _31245_ (.A(_10676_),
    .Y(_03762_));
 sky130_fd_sc_hd__nand2_1 _31246_ (.A(net836),
    .B(\inst$top.soc.cpu.divider.remainder[26] ),
    .Y(_10677_));
 sky130_fd_sc_hd__inv_1 _31247_ (.A(_10524_),
    .Y(_10678_));
 sky130_fd_sc_hd__nand2_1 _31248_ (.A(_10489_),
    .B(_10678_),
    .Y(_10679_));
 sky130_fd_sc_hd__nor3_1 _31249_ (.A(_10446_),
    .B(_10447_),
    .C(_10679_),
    .Y(_10680_));
 sky130_fd_sc_hd__inv_1 _31250_ (.A(_10606_),
    .Y(_10681_));
 sky130_fd_sc_hd__nand2_1 _31251_ (.A(_02768_),
    .B(_02771_),
    .Y(_10682_));
 sky130_fd_sc_hd__nor2_1 _31252_ (.A(_10642_),
    .B(_10682_),
    .Y(_10683_));
 sky130_fd_sc_hd__inv_1 _31253_ (.A(_10683_),
    .Y(_10684_));
 sky130_fd_sc_hd__nor2_1 _31254_ (.A(_10681_),
    .B(_10684_),
    .Y(_10685_));
 sky130_fd_sc_hd__nand3_1 _31255_ (.A(_10365_),
    .B(_10680_),
    .C(_10685_),
    .Y(_10686_));
 sky130_fd_sc_hd__nand3_1 _31256_ (.A(_10453_),
    .B(_10489_),
    .C(_10678_),
    .Y(_10687_));
 sky130_fd_sc_hd__o21a_1 _31257_ (.A1(_10524_),
    .A2(_10490_),
    .B1(_10525_),
    .X(_10688_));
 sky130_fd_sc_hd__nand2_1 _31258_ (.A(_10687_),
    .B(_10688_),
    .Y(_10689_));
 sky130_fd_sc_hd__a21oi_1 _31259_ (.A1(_02768_),
    .A2(_02770_),
    .B1(_02767_),
    .Y(_10690_));
 sky130_fd_sc_hd__o21ai_0 _31260_ (.A1(_10682_),
    .A2(_10643_),
    .B1(_10690_),
    .Y(_10691_));
 sky130_fd_sc_hd__a221oi_1 _31261_ (.A1(_10608_),
    .A2(_10683_),
    .B1(_10689_),
    .B2(_10685_),
    .C1(_10691_),
    .Y(_10692_));
 sky130_fd_sc_hd__nand2_1 _31262_ (.A(_10686_),
    .B(_10692_),
    .Y(_10693_));
 sky130_fd_sc_hd__xor2_1 _31263_ (.A(_02765_),
    .B(_10693_),
    .X(_10694_));
 sky130_fd_sc_hd__nand3_1 _31264_ (.A(net857),
    .B(net1040),
    .C(_10694_),
    .Y(_10695_));
 sky130_fd_sc_hd__nor4_1 _31265_ (.A(\inst$top.soc.cpu.divider.remainder[23] ),
    .B(\inst$top.soc.cpu.divider.remainder[24] ),
    .C(\inst$top.soc.cpu.divider.remainder[25] ),
    .D(\inst$top.soc.cpu.divider.remainder[26] ),
    .Y(_10696_));
 sky130_fd_sc_hd__inv_1 _31266_ (.A(_10696_),
    .Y(_10697_));
 sky130_fd_sc_hd__o21ai_0 _31267_ (.A1(_10697_),
    .A2(_10615_),
    .B1(\inst$top.soc.cpu.divider.remainder[27] ),
    .Y(_10698_));
 sky130_fd_sc_hd__inv_1 _31268_ (.A(\inst$top.soc.cpu.divider.remainder[27] ),
    .Y(_10699_));
 sky130_fd_sc_hd__nand4_1 _31269_ (.A(_10532_),
    .B(_10699_),
    .C(_10614_),
    .D(_10696_),
    .Y(_10700_));
 sky130_fd_sc_hd__nand3_1 _31270_ (.A(_10698_),
    .B(_10700_),
    .C(net1664),
    .Y(_10701_));
 sky130_fd_sc_hd__nand3_1 _31271_ (.A(_10677_),
    .B(_10695_),
    .C(_10701_),
    .Y(_10702_));
 sky130_fd_sc_hd__nand2_1 _31272_ (.A(_10702_),
    .B(net2928),
    .Y(_10703_));
 sky130_fd_sc_hd__nand2_1 _31273_ (.A(net608),
    .B(net1453),
    .Y(_10704_));
 sky130_fd_sc_hd__nand3_1 _31274_ (.A(_10703_),
    .B(net725),
    .C(_10704_),
    .Y(_10705_));
 sky130_fd_sc_hd__a21oi_1 _31275_ (.A1(net751),
    .A2(_10699_),
    .B1(net2976),
    .Y(_10706_));
 sky130_fd_sc_hd__nand2_1 _31276_ (.A(_10705_),
    .B(_10706_),
    .Y(_10707_));
 sky130_fd_sc_hd__inv_2 _31277_ (.A(_10707_),
    .Y(_03763_));
 sky130_fd_sc_hd__nand4_1 _31278_ (.A(_10664_),
    .B(_10668_),
    .C(_10699_),
    .D(_10593_),
    .Y(_10708_));
 sky130_fd_sc_hd__nor3_1 _31279_ (.A(\inst$top.soc.cpu.divider.remainder[28] ),
    .B(_10708_),
    .C(_10555_),
    .Y(_10709_));
 sky130_fd_sc_hd__o21ai_0 _31280_ (.A1(_10708_),
    .A2(_10555_),
    .B1(\inst$top.soc.cpu.divider.remainder[28] ),
    .Y(_10710_));
 sky130_fd_sc_hd__nand2_1 _31281_ (.A(_10710_),
    .B(net1664),
    .Y(_10711_));
 sky130_fd_sc_hd__xor2_1 _31282_ (.A(_02762_),
    .B(_09983_),
    .X(_10712_));
 sky130_fd_sc_hd__nand3_1 _31283_ (.A(net857),
    .B(net1039),
    .C(_10712_),
    .Y(_10713_));
 sky130_fd_sc_hd__nand2_1 _31284_ (.A(net835),
    .B(\inst$top.soc.cpu.divider.remainder[27] ),
    .Y(_10714_));
 sky130_fd_sc_hd__o211ai_1 _31285_ (.A1(_10709_),
    .A2(_10711_),
    .B1(_10713_),
    .C1(_10714_),
    .Y(_10715_));
 sky130_fd_sc_hd__nand2_1 _31286_ (.A(_10715_),
    .B(net2928),
    .Y(_10716_));
 sky130_fd_sc_hd__o21ai_1 _31287_ (.A1(net1460),
    .A2(net749),
    .B1(net610),
    .Y(_10717_));
 sky130_fd_sc_hd__o21ai_0 _31288_ (.A1(\inst$top.soc.cpu.divider.remainder[28] ),
    .A2(net725),
    .B1(net2116),
    .Y(_10718_));
 sky130_fd_sc_hd__a21oi_4 _31289_ (.A1(_10716_),
    .A2(_10717_),
    .B1(_10718_),
    .Y(_03764_));
 sky130_fd_sc_hd__a21oi_1 _31290_ (.A1(net607),
    .A2(net1468),
    .B1(net749),
    .Y(_10719_));
 sky130_fd_sc_hd__nor4_1 _31291_ (.A(_10447_),
    .B(_10488_),
    .C(_10524_),
    .D(_10572_),
    .Y(_10720_));
 sky130_fd_sc_hd__nor2_1 _31292_ (.A(_10605_),
    .B(_10642_),
    .Y(_10721_));
 sky130_fd_sc_hd__nand2_1 _31293_ (.A(_02762_),
    .B(_02765_),
    .Y(_10722_));
 sky130_fd_sc_hd__nor2_1 _31294_ (.A(_10682_),
    .B(_10722_),
    .Y(_10723_));
 sky130_fd_sc_hd__nand4_1 _31295_ (.A(_10406_),
    .B(_10720_),
    .C(_10721_),
    .D(_10723_),
    .Y(_10724_));
 sky130_fd_sc_hd__o21ai_0 _31296_ (.A1(_10642_),
    .A2(_10607_),
    .B1(_10643_),
    .Y(_10725_));
 sky130_fd_sc_hd__a21oi_1 _31297_ (.A1(_02762_),
    .A2(_02764_),
    .B1(_02761_),
    .Y(_10726_));
 sky130_fd_sc_hd__o21ai_0 _31298_ (.A1(_10722_),
    .A2(_10690_),
    .B1(_10726_),
    .Y(_10727_));
 sky130_fd_sc_hd__nand2_1 _31299_ (.A(_10721_),
    .B(_10723_),
    .Y(_10728_));
 sky130_fd_sc_hd__o21ai_0 _31300_ (.A1(_10488_),
    .A2(_10452_),
    .B1(_10490_),
    .Y(_10729_));
 sky130_fd_sc_hd__o21ai_0 _31301_ (.A1(_10572_),
    .A2(_10525_),
    .B1(_10574_),
    .Y(_10730_));
 sky130_fd_sc_hd__a31oi_1 _31302_ (.A1(_10729_),
    .A2(_10678_),
    .A3(_10573_),
    .B1(_10730_),
    .Y(_10731_));
 sky130_fd_sc_hd__nor2_1 _31303_ (.A(_10728_),
    .B(_10731_),
    .Y(_10732_));
 sky130_fd_sc_hd__a211oi_1 _31304_ (.A1(_10725_),
    .A2(_10723_),
    .B1(_10727_),
    .C1(_10732_),
    .Y(_10733_));
 sky130_fd_sc_hd__nand2_1 _31305_ (.A(_10724_),
    .B(_10733_),
    .Y(_10734_));
 sky130_fd_sc_hd__xor2_1 _31306_ (.A(_02759_),
    .B(_10734_),
    .X(_10735_));
 sky130_fd_sc_hd__nand3_1 _31307_ (.A(_10735_),
    .B(net1039),
    .C(net857),
    .Y(_10736_));
 sky130_fd_sc_hd__nand2_1 _31308_ (.A(net835),
    .B(\inst$top.soc.cpu.divider.remainder[28] ),
    .Y(_10737_));
 sky130_fd_sc_hd__nor2_1 _31309_ (.A(\inst$top.soc.cpu.divider.remainder[27] ),
    .B(\inst$top.soc.cpu.divider.remainder[28] ),
    .Y(_10738_));
 sky130_fd_sc_hd__nand4_1 _31310_ (.A(_10532_),
    .B(_10614_),
    .C(_10696_),
    .D(_10738_),
    .Y(_10739_));
 sky130_fd_sc_hd__xor2_1 _31311_ (.A(\inst$top.soc.cpu.divider.remainder[29] ),
    .B(_10739_),
    .X(_10740_));
 sky130_fd_sc_hd__nand2_1 _31312_ (.A(_10740_),
    .B(net1666),
    .Y(_10741_));
 sky130_fd_sc_hd__nand3_1 _31313_ (.A(_10736_),
    .B(_10737_),
    .C(_10741_),
    .Y(_10742_));
 sky130_fd_sc_hd__nand2_1 _31314_ (.A(_10742_),
    .B(net2929),
    .Y(_10743_));
 sky130_fd_sc_hd__nand2_1 _31315_ (.A(_10719_),
    .B(_10743_),
    .Y(_10744_));
 sky130_fd_sc_hd__inv_1 _31316_ (.A(\inst$top.soc.cpu.divider.remainder[29] ),
    .Y(_10745_));
 sky130_fd_sc_hd__a21oi_1 _31317_ (.A1(net750),
    .A2(_10745_),
    .B1(net2977),
    .Y(_10746_));
 sky130_fd_sc_hd__nand2_1 _31318_ (.A(_10744_),
    .B(_10746_),
    .Y(_10747_));
 sky130_fd_sc_hd__inv_2 _31319_ (.A(_10747_),
    .Y(_03765_));
 sky130_fd_sc_hd__a21oi_1 _31320_ (.A1(net607),
    .A2(net1153),
    .B1(net749),
    .Y(_10748_));
 sky130_fd_sc_hd__xor2_1 _31321_ (.A(\inst$top.soc.cpu.divider.remainder[2] ),
    .B(_02855_),
    .X(_10749_));
 sky130_fd_sc_hd__nor2_1 _31322_ (.A(_10749_),
    .B(net1245),
    .Y(_10750_));
 sky130_fd_sc_hd__xor2_1 _31323_ (.A(_02543_),
    .B(_02840_),
    .X(_10751_));
 sky130_fd_sc_hd__nand3_1 _31324_ (.A(net857),
    .B(net1039),
    .C(_10751_),
    .Y(_10752_));
 sky130_fd_sc_hd__nand3_1 _31325_ (.A(net852),
    .B(\inst$top.soc.cpu.divider.remainder[1] ),
    .C(net1039),
    .Y(_10753_));
 sky130_fd_sc_hd__nand2_1 _31326_ (.A(_10752_),
    .B(_10753_),
    .Y(_10754_));
 sky130_fd_sc_hd__o21ai_0 _31327_ (.A1(_10750_),
    .A2(_10754_),
    .B1(net2928),
    .Y(_10755_));
 sky130_fd_sc_hd__nand2_1 _31328_ (.A(_10748_),
    .B(_10755_),
    .Y(_10756_));
 sky130_fd_sc_hd__a21oi_1 _31329_ (.A1(net751),
    .A2(_10328_),
    .B1(net2976),
    .Y(_10757_));
 sky130_fd_sc_hd__nand2_1 _31330_ (.A(_10756_),
    .B(_10757_),
    .Y(_10758_));
 sky130_fd_sc_hd__inv_2 _31331_ (.A(_10758_),
    .Y(_03766_));
 sky130_fd_sc_hd__nand2_1 _31332_ (.A(net835),
    .B(\inst$top.soc.cpu.divider.remainder[29] ),
    .Y(_10759_));
 sky130_fd_sc_hd__nor2_1 _31333_ (.A(_09986_),
    .B(_09977_),
    .Y(_10760_));
 sky130_fd_sc_hd__o21ai_0 _31334_ (.A1(_09986_),
    .A2(_09981_),
    .B1(_09988_),
    .Y(_10761_));
 sky130_fd_sc_hd__a21oi_1 _31335_ (.A1(_10660_),
    .A2(_10760_),
    .B1(_10761_),
    .Y(_10762_));
 sky130_fd_sc_hd__xor2_1 _31336_ (.A(_09985_),
    .B(_10762_),
    .X(_10763_));
 sky130_fd_sc_hd__nand3_1 _31337_ (.A(net857),
    .B(net1039),
    .C(_10763_),
    .Y(_10764_));
 sky130_fd_sc_hd__nand4_1 _31338_ (.A(_10667_),
    .B(_10668_),
    .C(_10745_),
    .D(_10738_),
    .Y(_10765_));
 sky130_fd_sc_hd__xor2_1 _31339_ (.A(\inst$top.soc.cpu.divider.remainder[30] ),
    .B(_10765_),
    .X(_10766_));
 sky130_fd_sc_hd__nand2_1 _31340_ (.A(_10766_),
    .B(net1664),
    .Y(_10767_));
 sky130_fd_sc_hd__nand3_1 _31341_ (.A(_10759_),
    .B(_10764_),
    .C(_10767_),
    .Y(_10768_));
 sky130_fd_sc_hd__nand2_1 _31342_ (.A(_10768_),
    .B(net2929),
    .Y(_10769_));
 sky130_fd_sc_hd__nand2_1 _31343_ (.A(net607),
    .B(net1475),
    .Y(_10770_));
 sky130_fd_sc_hd__nand3_1 _31344_ (.A(_10769_),
    .B(net726),
    .C(_10770_),
    .Y(_10771_));
 sky130_fd_sc_hd__inv_1 _31345_ (.A(\inst$top.soc.cpu.divider.remainder[30] ),
    .Y(_10772_));
 sky130_fd_sc_hd__a21oi_1 _31346_ (.A1(net750),
    .A2(_10772_),
    .B1(net2977),
    .Y(_10773_));
 sky130_fd_sc_hd__nand2_1 _31347_ (.A(_10771_),
    .B(_10773_),
    .Y(_10774_));
 sky130_fd_sc_hd__inv_2 _31348_ (.A(_10774_),
    .Y(_03767_));
 sky130_fd_sc_hd__nand2_1 _31349_ (.A(net836),
    .B(\inst$top.soc.cpu.divider.remainder[30] ),
    .Y(_10775_));
 sky130_fd_sc_hd__inv_1 _31350_ (.A(_02759_),
    .Y(_10776_));
 sky130_fd_sc_hd__nor3_1 _31351_ (.A(_09985_),
    .B(_10776_),
    .C(_10722_),
    .Y(_10777_));
 sky130_fd_sc_hd__nand2_1 _31352_ (.A(_10693_),
    .B(_10777_),
    .Y(_10778_));
 sky130_fd_sc_hd__o21bai_1 _31353_ (.A1(_10776_),
    .A2(_10726_),
    .B1_N(_02758_),
    .Y(_10779_));
 sky130_fd_sc_hd__a21oi_1 _31354_ (.A1(_10779_),
    .A2(_02756_),
    .B1(_02755_),
    .Y(_10780_));
 sky130_fd_sc_hd__nand2_1 _31355_ (.A(_10778_),
    .B(_10780_),
    .Y(_10781_));
 sky130_fd_sc_hd__xor2_1 _31356_ (.A(_02753_),
    .B(_10781_),
    .X(_10782_));
 sky130_fd_sc_hd__nand3_1 _31357_ (.A(net857),
    .B(_10782_),
    .C(net1039),
    .Y(_10783_));
 sky130_fd_sc_hd__nand3_1 _31358_ (.A(_10738_),
    .B(_10745_),
    .C(_10772_),
    .Y(_10784_));
 sky130_fd_sc_hd__nor3_1 _31359_ (.A(_10697_),
    .B(_10784_),
    .C(_10615_),
    .Y(_10785_));
 sky130_fd_sc_hd__xor2_1 _31360_ (.A(_09930_),
    .B(_10785_),
    .X(_10786_));
 sky130_fd_sc_hd__nand2_1 _31361_ (.A(_10786_),
    .B(net1664),
    .Y(_10787_));
 sky130_fd_sc_hd__nand3_1 _31362_ (.A(_10775_),
    .B(_10783_),
    .C(_10787_),
    .Y(_10788_));
 sky130_fd_sc_hd__nand2_1 _31363_ (.A(_10788_),
    .B(net2929),
    .Y(_10789_));
 sky130_fd_sc_hd__nand2_1 _31364_ (.A(net606),
    .B(net1482),
    .Y(_10790_));
 sky130_fd_sc_hd__nand3_1 _31365_ (.A(_10789_),
    .B(net726),
    .C(_10790_),
    .Y(_10791_));
 sky130_fd_sc_hd__a21oi_1 _31366_ (.A1(net749),
    .A2(_09930_),
    .B1(net2977),
    .Y(_10792_));
 sky130_fd_sc_hd__nand2_1 _31367_ (.A(_10791_),
    .B(_10792_),
    .Y(_10793_));
 sky130_fd_sc_hd__inv_2 _31368_ (.A(_10793_),
    .Y(_03768_));
 sky130_fd_sc_hd__nand2_1 _31369_ (.A(net606),
    .B(net1361),
    .Y(_10794_));
 sky130_fd_sc_hd__nand2_1 _31370_ (.A(_10356_),
    .B(_02837_),
    .Y(_10795_));
 sky130_fd_sc_hd__nand3_1 _31371_ (.A(_10354_),
    .B(_10352_),
    .C(_10355_),
    .Y(_10796_));
 sky130_fd_sc_hd__nand4_1 _31372_ (.A(net856),
    .B(net1039),
    .C(_10795_),
    .D(_10796_),
    .Y(_10797_));
 sky130_fd_sc_hd__nand2_1 _31373_ (.A(net836),
    .B(\inst$top.soc.cpu.divider.remainder[2] ),
    .Y(_10798_));
 sky130_fd_sc_hd__xor2_1 _31374_ (.A(_10329_),
    .B(_10368_),
    .X(_10799_));
 sky130_fd_sc_hd__a21oi_1 _31375_ (.A1(net1102),
    .A2(_10799_),
    .B1(net751),
    .Y(_10800_));
 sky130_fd_sc_hd__nand4_1 _31376_ (.A(_10794_),
    .B(_10797_),
    .C(_10798_),
    .D(_10800_),
    .Y(_10801_));
 sky130_fd_sc_hd__a21oi_1 _31377_ (.A1(net751),
    .A2(_10329_),
    .B1(net2975),
    .Y(_10802_));
 sky130_fd_sc_hd__nand2_1 _31378_ (.A(_10801_),
    .B(_10802_),
    .Y(_10803_));
 sky130_fd_sc_hd__inv_2 _31379_ (.A(_10803_),
    .Y(_03769_));
 sky130_fd_sc_hd__a21oi_1 _31380_ (.A1(net608),
    .A2(net1356),
    .B1(net751),
    .Y(_10804_));
 sky130_fd_sc_hd__nand3_1 _31381_ (.A(_02543_),
    .B(_02837_),
    .C(_02840_),
    .Y(_10805_));
 sky130_fd_sc_hd__nand2_1 _31382_ (.A(_09935_),
    .B(_10805_),
    .Y(_10806_));
 sky130_fd_sc_hd__nand2_1 _31383_ (.A(_10806_),
    .B(_02834_),
    .Y(_10807_));
 sky130_fd_sc_hd__nand3_1 _31384_ (.A(_09935_),
    .B(_10351_),
    .C(_10805_),
    .Y(_10808_));
 sky130_fd_sc_hd__nand4_1 _31385_ (.A(net856),
    .B(net1038),
    .C(_10807_),
    .D(_10808_),
    .Y(_10809_));
 sky130_fd_sc_hd__nand2_1 _31386_ (.A(net836),
    .B(\inst$top.soc.cpu.divider.remainder[3] ),
    .Y(_10810_));
 sky130_fd_sc_hd__nand3_1 _31387_ (.A(_10809_),
    .B(_10810_),
    .C(net1245),
    .Y(_10811_));
 sky130_fd_sc_hd__nand3_1 _31388_ (.A(_10328_),
    .B(_10329_),
    .C(_02855_),
    .Y(_10812_));
 sky130_fd_sc_hd__xor2_1 _31389_ (.A(_10369_),
    .B(_10812_),
    .X(_10813_));
 sky130_fd_sc_hd__a21oi_1 _31390_ (.A1(_10813_),
    .A2(net1664),
    .B1(net2025),
    .Y(_10814_));
 sky130_fd_sc_hd__nand2_1 _31391_ (.A(_10811_),
    .B(_10814_),
    .Y(_10815_));
 sky130_fd_sc_hd__nand2_1 _31392_ (.A(_10804_),
    .B(_10815_),
    .Y(_10816_));
 sky130_fd_sc_hd__a21oi_1 _31394_ (.A1(net751),
    .A2(_10369_),
    .B1(net2976),
    .Y(_10818_));
 sky130_fd_sc_hd__nand2_1 _31395_ (.A(_10816_),
    .B(_10818_),
    .Y(_10819_));
 sky130_fd_sc_hd__inv_2 _31396_ (.A(_10819_),
    .Y(_03770_));
 sky130_fd_sc_hd__inv_1 _31397_ (.A(_02836_),
    .Y(_10820_));
 sky130_fd_sc_hd__a21oi_1 _31398_ (.A1(_10795_),
    .A2(_10820_),
    .B1(_10351_),
    .Y(_10821_));
 sky130_fd_sc_hd__nor2_1 _31399_ (.A(_02833_),
    .B(_10821_),
    .Y(_10822_));
 sky130_fd_sc_hd__xor2_1 _31400_ (.A(_02831_),
    .B(_10822_),
    .X(_10823_));
 sky130_fd_sc_hd__nand3b_1 _31401_ (.A_N(_10823_),
    .B(net856),
    .C(net1038),
    .Y(_10824_));
 sky130_fd_sc_hd__nand3_1 _31402_ (.A(net852),
    .B(\inst$top.soc.cpu.divider.remainder[4] ),
    .C(net1038),
    .Y(_10825_));
 sky130_fd_sc_hd__xor2_1 _31403_ (.A(\inst$top.soc.cpu.divider.remainder[5] ),
    .B(_10370_),
    .X(_10826_));
 sky130_fd_sc_hd__nand2_1 _31404_ (.A(_10826_),
    .B(net1664),
    .Y(_10827_));
 sky130_fd_sc_hd__nand3_1 _31405_ (.A(_10824_),
    .B(_10825_),
    .C(_10827_),
    .Y(_10828_));
 sky130_fd_sc_hd__nand2_1 _31406_ (.A(_10828_),
    .B(net2925),
    .Y(_10829_));
 sky130_fd_sc_hd__nand2_1 _31407_ (.A(net605),
    .B(net1351),
    .Y(_10830_));
 sky130_fd_sc_hd__nand3_1 _31408_ (.A(_10829_),
    .B(_10830_),
    .C(net725),
    .Y(_10831_));
 sky130_fd_sc_hd__inv_1 _31409_ (.A(\inst$top.soc.cpu.divider.remainder[5] ),
    .Y(_10832_));
 sky130_fd_sc_hd__a21oi_1 _31410_ (.A1(net751),
    .A2(_10832_),
    .B1(net2974),
    .Y(_10833_));
 sky130_fd_sc_hd__nand2_1 _31411_ (.A(_10831_),
    .B(_10833_),
    .Y(_10834_));
 sky130_fd_sc_hd__inv_2 _31412_ (.A(_10834_),
    .Y(_03771_));
 sky130_fd_sc_hd__xnor2_1 _31413_ (.A(_02828_),
    .B(_09938_),
    .Y(_10835_));
 sky130_fd_sc_hd__nand3_1 _31414_ (.A(net855),
    .B(net1034),
    .C(_10835_),
    .Y(_10836_));
 sky130_fd_sc_hd__nand3_1 _31415_ (.A(net852),
    .B(\inst$top.soc.cpu.divider.remainder[5] ),
    .C(net1034),
    .Y(_10837_));
 sky130_fd_sc_hd__xor2_1 _31416_ (.A(\inst$top.soc.cpu.divider.remainder[6] ),
    .B(_10330_),
    .X(_10838_));
 sky130_fd_sc_hd__nand2_1 _31417_ (.A(_10838_),
    .B(net1665),
    .Y(_10839_));
 sky130_fd_sc_hd__nand3_1 _31418_ (.A(_10836_),
    .B(_10837_),
    .C(_10839_),
    .Y(_10840_));
 sky130_fd_sc_hd__nand2_1 _31419_ (.A(_10840_),
    .B(net2925),
    .Y(_10841_));
 sky130_fd_sc_hd__nand2_1 _31420_ (.A(net605),
    .B(net1350),
    .Y(_10842_));
 sky130_fd_sc_hd__nand3_1 _31421_ (.A(_10841_),
    .B(_10842_),
    .C(net724),
    .Y(_10843_));
 sky130_fd_sc_hd__a21oi_1 _31422_ (.A1(net745),
    .A2(_10322_),
    .B1(net2974),
    .Y(_10844_));
 sky130_fd_sc_hd__nand2_1 _31423_ (.A(_10843_),
    .B(_10844_),
    .Y(_10845_));
 sky130_fd_sc_hd__inv_2 _31424_ (.A(_10845_),
    .Y(_03772_));
 sky130_fd_sc_hd__a21oi_1 _31425_ (.A1(net605),
    .A2(net1346),
    .B1(net745),
    .Y(_10846_));
 sky130_fd_sc_hd__nand2_1 _31426_ (.A(_10358_),
    .B(_02825_),
    .Y(_10847_));
 sky130_fd_sc_hd__nand3_1 _31427_ (.A(_10350_),
    .B(_10444_),
    .C(_10357_),
    .Y(_10848_));
 sky130_fd_sc_hd__nand4_1 _31428_ (.A(net854),
    .B(net1032),
    .C(_10847_),
    .D(_10848_),
    .Y(_10849_));
 sky130_fd_sc_hd__nand2_1 _31429_ (.A(net835),
    .B(\inst$top.soc.cpu.divider.remainder[6] ),
    .Y(_10850_));
 sky130_fd_sc_hd__xor2_1 _31430_ (.A(_10323_),
    .B(_10371_),
    .X(_10851_));
 sky130_fd_sc_hd__nand2_1 _31431_ (.A(_10851_),
    .B(net1665),
    .Y(_10852_));
 sky130_fd_sc_hd__nand3_1 _31432_ (.A(_10849_),
    .B(_10850_),
    .C(_10852_),
    .Y(_10853_));
 sky130_fd_sc_hd__nand2_1 _31433_ (.A(_10853_),
    .B(net2927),
    .Y(_10854_));
 sky130_fd_sc_hd__nand2_1 _31434_ (.A(_10846_),
    .B(_10854_),
    .Y(_10855_));
 sky130_fd_sc_hd__a21oi_1 _31435_ (.A1(net744),
    .A2(_10323_),
    .B1(net2978),
    .Y(_10856_));
 sky130_fd_sc_hd__nand2_1 _31436_ (.A(_10855_),
    .B(_10856_),
    .Y(_10857_));
 sky130_fd_sc_hd__inv_2 _31437_ (.A(_10857_),
    .Y(_03773_));
 sky130_fd_sc_hd__xor2_1 _31438_ (.A(_02822_),
    .B(_09940_),
    .X(_10858_));
 sky130_fd_sc_hd__nand3_1 _31439_ (.A(net854),
    .B(net1032),
    .C(_10858_),
    .Y(_10859_));
 sky130_fd_sc_hd__nand3_1 _31440_ (.A(net852),
    .B(\inst$top.soc.cpu.divider.remainder[7] ),
    .C(net1032),
    .Y(_10860_));
 sky130_fd_sc_hd__xor2_1 _31441_ (.A(_10324_),
    .B(_10391_),
    .X(_10861_));
 sky130_fd_sc_hd__nand2_1 _31442_ (.A(_10861_),
    .B(net1665),
    .Y(_10862_));
 sky130_fd_sc_hd__nand3_1 _31443_ (.A(_10859_),
    .B(_10860_),
    .C(_10862_),
    .Y(_10863_));
 sky130_fd_sc_hd__nand2_1 _31444_ (.A(_10863_),
    .B(net2927),
    .Y(_10864_));
 sky130_fd_sc_hd__nand2_1 _31445_ (.A(net606),
    .B(net1341),
    .Y(_10865_));
 sky130_fd_sc_hd__nand3_1 _31446_ (.A(_10864_),
    .B(_10865_),
    .C(net723),
    .Y(_10866_));
 sky130_fd_sc_hd__a21oi_1 _31447_ (.A1(net746),
    .A2(_10324_),
    .B1(net2967),
    .Y(_10867_));
 sky130_fd_sc_hd__nand2_1 _31448_ (.A(_10866_),
    .B(_10867_),
    .Y(_10868_));
 sky130_fd_sc_hd__inv_2 _31449_ (.A(_10868_),
    .Y(_03774_));
 sky130_fd_sc_hd__xor2_1 _31450_ (.A(_02819_),
    .B(_10360_),
    .X(_10869_));
 sky130_fd_sc_hd__nand3_1 _31451_ (.A(net854),
    .B(net1032),
    .C(_10869_),
    .Y(_10870_));
 sky130_fd_sc_hd__nand3_1 _31452_ (.A(net852),
    .B(\inst$top.soc.cpu.divider.remainder[8] ),
    .C(net1032),
    .Y(_10871_));
 sky130_fd_sc_hd__nand2_1 _31453_ (.A(_10371_),
    .B(_10372_),
    .Y(_10872_));
 sky130_fd_sc_hd__a21oi_1 _31454_ (.A1(_10872_),
    .A2(\inst$top.soc.cpu.divider.remainder[9] ),
    .B1(net1245),
    .Y(_10873_));
 sky130_fd_sc_hd__o21ai_0 _31455_ (.A1(\inst$top.soc.cpu.divider.remainder[9] ),
    .A2(_10872_),
    .B1(_10873_),
    .Y(_10874_));
 sky130_fd_sc_hd__nand3_1 _31456_ (.A(_10870_),
    .B(_10871_),
    .C(_10874_),
    .Y(_10875_));
 sky130_fd_sc_hd__nand2_1 _31457_ (.A(_10875_),
    .B(net2927),
    .Y(_10876_));
 sky130_fd_sc_hd__nand2_1 _31458_ (.A(net605),
    .B(net1337),
    .Y(_10877_));
 sky130_fd_sc_hd__nand3_1 _31459_ (.A(_10876_),
    .B(_10877_),
    .C(net723),
    .Y(_10878_));
 sky130_fd_sc_hd__a21oi_1 _31460_ (.A1(net744),
    .A2(_10325_),
    .B1(net2967),
    .Y(_10879_));
 sky130_fd_sc_hd__nand2_1 _31461_ (.A(_10878_),
    .B(_10879_),
    .Y(_10880_));
 sky130_fd_sc_hd__inv_2 _31462_ (.A(_10880_),
    .Y(_03775_));
 sky130_fd_sc_hd__nand2_1 _31463_ (.A(net611),
    .B(net1104),
    .Y(_10881_));
 sky130_fd_sc_hd__nand2_1 _31464_ (.A(_10881_),
    .B(\inst$top.soc.cpu.divider.timer[0] ),
    .Y(_10882_));
 sky130_fd_sc_hd__a21oi_1 _31465_ (.A1(net1104),
    .A2(_02857_),
    .B1(net2967),
    .Y(_10883_));
 sky130_fd_sc_hd__nand2_1 _31466_ (.A(_10882_),
    .B(_10883_),
    .Y(_10884_));
 sky130_fd_sc_hd__inv_2 _31467_ (.A(_10884_),
    .Y(_03776_));
 sky130_fd_sc_hd__nand3_1 _31468_ (.A(net611),
    .B(\inst$top.soc.cpu.divider.timer[1] ),
    .C(net1104),
    .Y(_10885_));
 sky130_fd_sc_hd__or2_2 _31469_ (.A(_02860_),
    .B(net1104),
    .X(_10886_));
 sky130_fd_sc_hd__a21oi_4 _31470_ (.A1(_10885_),
    .A2(_10886_),
    .B1(net2967),
    .Y(_03777_));
 sky130_fd_sc_hd__xnor2_1 _31471_ (.A(\inst$top.soc.cpu.divider.timer[2] ),
    .B(_02859_),
    .Y(_10887_));
 sky130_fd_sc_hd__nor2_1 _31472_ (.A(net2026),
    .B(_10887_),
    .Y(_10888_));
 sky130_fd_sc_hd__nand2_1 _31473_ (.A(_10881_),
    .B(_10888_),
    .Y(_10889_));
 sky130_fd_sc_hd__nand3_2 _31474_ (.A(net611),
    .B(\inst$top.soc.cpu.divider.timer[2] ),
    .C(net1104),
    .Y(_10890_));
 sky130_fd_sc_hd__a21oi_4 _31475_ (.A1(_10889_),
    .A2(_10890_),
    .B1(net2967),
    .Y(_03778_));
 sky130_fd_sc_hd__nor2_1 _31476_ (.A(\inst$top.soc.cpu.divider.timer[2] ),
    .B(\inst$top.soc.cpu.divider.timer[1] ),
    .Y(_10891_));
 sky130_fd_sc_hd__nand2_1 _31477_ (.A(_10891_),
    .B(_02857_),
    .Y(_10892_));
 sky130_fd_sc_hd__xor2_1 _31478_ (.A(\inst$top.soc.cpu.divider.timer[3] ),
    .B(_10892_),
    .X(_10893_));
 sky130_fd_sc_hd__nor2_1 _31479_ (.A(net2026),
    .B(_10893_),
    .Y(_10894_));
 sky130_fd_sc_hd__nand2_1 _31480_ (.A(_10881_),
    .B(_10894_),
    .Y(_10895_));
 sky130_fd_sc_hd__nand3_2 _31481_ (.A(net611),
    .B(\inst$top.soc.cpu.divider.timer[3] ),
    .C(net1104),
    .Y(_10896_));
 sky130_fd_sc_hd__a21oi_4 _31482_ (.A1(_10895_),
    .A2(_10896_),
    .B1(net2967),
    .Y(_03779_));
 sky130_fd_sc_hd__xor2_1 _31483_ (.A(\inst$top.soc.cpu.divider.timer[4] ),
    .B(_09905_),
    .X(_10897_));
 sky130_fd_sc_hd__nor2_1 _31484_ (.A(net2026),
    .B(_10897_),
    .Y(_10898_));
 sky130_fd_sc_hd__nand2_1 _31485_ (.A(_10881_),
    .B(_10898_),
    .Y(_10899_));
 sky130_fd_sc_hd__nand3_2 _31486_ (.A(net611),
    .B(\inst$top.soc.cpu.divider.timer[4] ),
    .C(net1104),
    .Y(_10900_));
 sky130_fd_sc_hd__a21oi_4 _31487_ (.A1(_10899_),
    .A2(_10900_),
    .B1(net2967),
    .Y(_03780_));
 sky130_fd_sc_hd__nor2_1 _31488_ (.A(\inst$top.soc.cpu.divider.timer[3] ),
    .B(\inst$top.soc.cpu.divider.timer[4] ),
    .Y(_10901_));
 sky130_fd_sc_hd__nand3_1 _31489_ (.A(_10891_),
    .B(_10901_),
    .C(_02857_),
    .Y(_10902_));
 sky130_fd_sc_hd__or2_2 _31490_ (.A(\inst$top.soc.cpu.divider.timer[5] ),
    .B(_10902_),
    .X(_10903_));
 sky130_fd_sc_hd__nand2_1 _31491_ (.A(_10902_),
    .B(\inst$top.soc.cpu.divider.timer[5] ),
    .Y(_10904_));
 sky130_fd_sc_hd__nand3_1 _31492_ (.A(_10903_),
    .B(net2927),
    .C(_10904_),
    .Y(_10905_));
 sky130_fd_sc_hd__nand2_1 _31493_ (.A(_10881_),
    .B(_10905_),
    .Y(_10906_));
 sky130_fd_sc_hd__nand3_1 _31496_ (.A(net611),
    .B(\inst$top.soc.cpu.divider.timer[5] ),
    .C(net1104),
    .Y(_10909_));
 sky130_fd_sc_hd__nand3_2 _31497_ (.A(_10906_),
    .B(net2118),
    .C(_10909_),
    .Y(_03781_));
 sky130_fd_sc_hd__nand2_1 _31498_ (.A(\inst$top.soc.cpu.d.sink__payload$16.csr_rdy ),
    .B(\inst$top.soc.cpu.csrf.bank_300_w_select ),
    .Y(_10910_));
 sky130_fd_sc_hd__nor2_1 _31499_ (.A(_10910_),
    .B(_20368_),
    .Y(_10911_));
 sky130_fd_sc_hd__nand2_1 _31500_ (.A(net1807),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause_w_select ),
    .Y(_10912_));
 sky130_fd_sc_hd__nand2_1 _31501_ (.A(\inst$top.soc.cpu.exception.w_trap ),
    .B(\inst$top.soc.cpu.m.source__valid ),
    .Y(_10913_));
 sky130_fd_sc_hd__nand2_1 _31502_ (.A(_10912_),
    .B(_10913_),
    .Y(_10914_));
 sky130_fd_sc_hd__inv_1 _31503_ (.A(_10914_),
    .Y(_10915_));
 sky130_fd_sc_hd__nand2_1 _31505_ (.A(net1096),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[0] ),
    .Y(_10917_));
 sky130_fd_sc_hd__inv_1 _31506_ (.A(_10912_),
    .Y(_10918_));
 sky130_fd_sc_hd__nand2_1 _31508_ (.A(net1241),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[0] ),
    .Y(_10920_));
 sky130_fd_sc_hd__inv_2 _31509_ (.A(_10913_),
    .Y(_10921_));
 sky130_fd_sc_hd__nand2_1 _31512_ (.A(net1873),
    .B(\inst$top.soc.cpu.exception.w_data$48[0] ),
    .Y(_10924_));
 sky130_fd_sc_hd__a31oi_1 _31514_ (.A1(_10917_),
    .A2(_10920_),
    .A3(_10924_),
    .B1(net2960),
    .Y(_03782_));
 sky130_fd_sc_hd__nand2_1 _31516_ (.A(net1097),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[10] ),
    .Y(_10927_));
 sky130_fd_sc_hd__nand2_1 _31518_ (.A(net1242),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[10] ),
    .Y(_10929_));
 sky130_fd_sc_hd__a21oi_1 _31520_ (.A1(_10927_),
    .A2(_10929_),
    .B1(net2968),
    .Y(_03783_));
 sky130_fd_sc_hd__nand2_1 _31521_ (.A(net1099),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[11] ),
    .Y(_10931_));
 sky130_fd_sc_hd__nand2_1 _31522_ (.A(net1244),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[11] ),
    .Y(_10932_));
 sky130_fd_sc_hd__a21oi_1 _31523_ (.A1(_10931_),
    .A2(_10932_),
    .B1(net2961),
    .Y(_03784_));
 sky130_fd_sc_hd__nand2_1 _31524_ (.A(net1098),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[12] ),
    .Y(_10933_));
 sky130_fd_sc_hd__nand2_1 _31525_ (.A(net1243),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[12] ),
    .Y(_10934_));
 sky130_fd_sc_hd__a21oi_1 _31526_ (.A1(_10933_),
    .A2(_10934_),
    .B1(net2939),
    .Y(_03785_));
 sky130_fd_sc_hd__nand2_1 _31527_ (.A(net1097),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[13] ),
    .Y(_10935_));
 sky130_fd_sc_hd__nand2_1 _31528_ (.A(net1242),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[13] ),
    .Y(_10936_));
 sky130_fd_sc_hd__a21oi_1 _31529_ (.A1(_10935_),
    .A2(_10936_),
    .B1(net2968),
    .Y(_03786_));
 sky130_fd_sc_hd__nand2_1 _31530_ (.A(net1097),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[14] ),
    .Y(_10937_));
 sky130_fd_sc_hd__nand2_1 _31531_ (.A(net1242),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[14] ),
    .Y(_10938_));
 sky130_fd_sc_hd__a21oi_1 _31532_ (.A1(_10937_),
    .A2(_10938_),
    .B1(net2952),
    .Y(_03787_));
 sky130_fd_sc_hd__nand2_1 _31533_ (.A(net1097),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[15] ),
    .Y(_10939_));
 sky130_fd_sc_hd__nand2_1 _31534_ (.A(net1242),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[15] ),
    .Y(_10940_));
 sky130_fd_sc_hd__a21oi_1 _31535_ (.A1(_10939_),
    .A2(_10940_),
    .B1(net2952),
    .Y(_03788_));
 sky130_fd_sc_hd__nand2_1 _31536_ (.A(net1096),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[16] ),
    .Y(_10941_));
 sky130_fd_sc_hd__nand2_1 _31537_ (.A(net1241),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[16] ),
    .Y(_10942_));
 sky130_fd_sc_hd__a21oi_1 _31538_ (.A1(_10941_),
    .A2(_10942_),
    .B1(net2958),
    .Y(_03789_));
 sky130_fd_sc_hd__nand2_1 _31539_ (.A(net1098),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[17] ),
    .Y(_10943_));
 sky130_fd_sc_hd__nand2_1 _31540_ (.A(net1243),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[17] ),
    .Y(_10944_));
 sky130_fd_sc_hd__a21oi_1 _31541_ (.A1(_10943_),
    .A2(_10944_),
    .B1(net2964),
    .Y(_03790_));
 sky130_fd_sc_hd__nand2_1 _31542_ (.A(net1098),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[18] ),
    .Y(_10945_));
 sky130_fd_sc_hd__nand2_1 _31543_ (.A(net1243),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[18] ),
    .Y(_10946_));
 sky130_fd_sc_hd__a21oi_1 _31544_ (.A1(_10945_),
    .A2(_10946_),
    .B1(net2964),
    .Y(_03791_));
 sky130_fd_sc_hd__nand2_1 _31545_ (.A(net1098),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[19] ),
    .Y(_10947_));
 sky130_fd_sc_hd__nand2_1 _31546_ (.A(net1243),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[19] ),
    .Y(_10948_));
 sky130_fd_sc_hd__a21oi_1 _31547_ (.A1(_10947_),
    .A2(_10948_),
    .B1(net2965),
    .Y(_03792_));
 sky130_fd_sc_hd__nand2_1 _31548_ (.A(net1096),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[1] ),
    .Y(_10949_));
 sky130_fd_sc_hd__nand2_1 _31549_ (.A(net1241),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[1] ),
    .Y(_10950_));
 sky130_fd_sc_hd__nand2_1 _31550_ (.A(net1873),
    .B(\inst$top.soc.cpu.exception.w_data$48[1] ),
    .Y(_10951_));
 sky130_fd_sc_hd__a31oi_1 _31551_ (.A1(_10949_),
    .A2(_10950_),
    .A3(_10951_),
    .B1(net2958),
    .Y(_03793_));
 sky130_fd_sc_hd__nand2_1 _31553_ (.A(net1099),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[20] ),
    .Y(_10953_));
 sky130_fd_sc_hd__nand2_1 _31555_ (.A(net1244),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[20] ),
    .Y(_10955_));
 sky130_fd_sc_hd__a21oi_1 _31557_ (.A1(_10953_),
    .A2(_10955_),
    .B1(net2965),
    .Y(_03794_));
 sky130_fd_sc_hd__nand2_1 _31558_ (.A(net1098),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[21] ),
    .Y(_10957_));
 sky130_fd_sc_hd__nand2_1 _31559_ (.A(net1243),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[21] ),
    .Y(_10958_));
 sky130_fd_sc_hd__a21oi_1 _31560_ (.A1(_10957_),
    .A2(_10958_),
    .B1(net2961),
    .Y(_03795_));
 sky130_fd_sc_hd__nand2_1 _31561_ (.A(net1098),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[22] ),
    .Y(_10959_));
 sky130_fd_sc_hd__nand2_1 _31562_ (.A(net1243),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[22] ),
    .Y(_10960_));
 sky130_fd_sc_hd__a21oi_1 _31563_ (.A1(_10959_),
    .A2(_10960_),
    .B1(net2971),
    .Y(_03796_));
 sky130_fd_sc_hd__nand2_1 _31564_ (.A(net1098),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[23] ),
    .Y(_10961_));
 sky130_fd_sc_hd__nand2_1 _31565_ (.A(net1243),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[23] ),
    .Y(_10962_));
 sky130_fd_sc_hd__a21oi_1 _31566_ (.A1(_10961_),
    .A2(_10962_),
    .B1(net2971),
    .Y(_03797_));
 sky130_fd_sc_hd__nand2_1 _31567_ (.A(net1099),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[24] ),
    .Y(_10963_));
 sky130_fd_sc_hd__nand2_1 _31568_ (.A(net1244),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[24] ),
    .Y(_10964_));
 sky130_fd_sc_hd__a21oi_1 _31569_ (.A1(_10963_),
    .A2(_10964_),
    .B1(net2969),
    .Y(_03798_));
 sky130_fd_sc_hd__nand2_1 _31570_ (.A(net1096),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[25] ),
    .Y(_10965_));
 sky130_fd_sc_hd__nand2_1 _31571_ (.A(net1241),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[25] ),
    .Y(_10966_));
 sky130_fd_sc_hd__a21oi_1 _31572_ (.A1(_10965_),
    .A2(_10966_),
    .B1(net2960),
    .Y(_03799_));
 sky130_fd_sc_hd__nand2_1 _31573_ (.A(net1097),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[26] ),
    .Y(_10967_));
 sky130_fd_sc_hd__nand2_1 _31574_ (.A(net1242),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[26] ),
    .Y(_10968_));
 sky130_fd_sc_hd__a21oi_1 _31575_ (.A1(_10967_),
    .A2(_10968_),
    .B1(net2971),
    .Y(_03800_));
 sky130_fd_sc_hd__nand2_1 _31576_ (.A(net1097),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[27] ),
    .Y(_10969_));
 sky130_fd_sc_hd__nand2_1 _31577_ (.A(net1242),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[27] ),
    .Y(_10970_));
 sky130_fd_sc_hd__a21oi_1 _31578_ (.A1(_10969_),
    .A2(_10970_),
    .B1(net2971),
    .Y(_03801_));
 sky130_fd_sc_hd__nand2_1 _31579_ (.A(net1097),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[28] ),
    .Y(_10971_));
 sky130_fd_sc_hd__nand2_1 _31580_ (.A(net1242),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[28] ),
    .Y(_10972_));
 sky130_fd_sc_hd__a21oi_1 _31581_ (.A1(_10971_),
    .A2(_10972_),
    .B1(net2969),
    .Y(_03802_));
 sky130_fd_sc_hd__nand2_1 _31582_ (.A(net1097),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[29] ),
    .Y(_10973_));
 sky130_fd_sc_hd__nand2_1 _31583_ (.A(net1242),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[29] ),
    .Y(_10974_));
 sky130_fd_sc_hd__a21oi_1 _31584_ (.A1(_10973_),
    .A2(_10974_),
    .B1(net2968),
    .Y(_03803_));
 sky130_fd_sc_hd__nand2_1 _31585_ (.A(net1096),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[2] ),
    .Y(_10975_));
 sky130_fd_sc_hd__nand2_1 _31586_ (.A(net1241),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[2] ),
    .Y(_10976_));
 sky130_fd_sc_hd__nand2_1 _31587_ (.A(net1874),
    .B(\inst$top.soc.cpu.exception.w_data$48[2] ),
    .Y(_10977_));
 sky130_fd_sc_hd__a31oi_1 _31590_ (.A1(_10975_),
    .A2(_10976_),
    .A3(_10977_),
    .B1(net2936),
    .Y(_03804_));
 sky130_fd_sc_hd__nand2_1 _31591_ (.A(net1097),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[30] ),
    .Y(_10980_));
 sky130_fd_sc_hd__nand2_1 _31592_ (.A(net1242),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[30] ),
    .Y(_10981_));
 sky130_fd_sc_hd__a21oi_1 _31595_ (.A1(_10980_),
    .A2(_10981_),
    .B1(net2962),
    .Y(_03805_));
 sky130_fd_sc_hd__nand2_1 _31596_ (.A(net1096),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[31] ),
    .Y(_10984_));
 sky130_fd_sc_hd__nand2_1 _31597_ (.A(net1241),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[31] ),
    .Y(_10985_));
 sky130_fd_sc_hd__nand2_1 _31598_ (.A(net1872),
    .B(\inst$top.soc.cpu.exception.w_data$48[31] ),
    .Y(_10986_));
 sky130_fd_sc_hd__a31oi_1 _31599_ (.A1(_10984_),
    .A2(_10985_),
    .A3(_10986_),
    .B1(net2937),
    .Y(_03806_));
 sky130_fd_sc_hd__nand2_1 _31600_ (.A(net1096),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[3] ),
    .Y(_10987_));
 sky130_fd_sc_hd__nand2_1 _31601_ (.A(net1241),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[3] ),
    .Y(_10988_));
 sky130_fd_sc_hd__nand2_1 _31602_ (.A(net1873),
    .B(\inst$top.soc.cpu.exception.w_data$48[3] ),
    .Y(_10989_));
 sky130_fd_sc_hd__a31oi_1 _31603_ (.A1(_10987_),
    .A2(_10988_),
    .A3(_10989_),
    .B1(net2958),
    .Y(_03807_));
 sky130_fd_sc_hd__nand2_1 _31604_ (.A(net1096),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[4] ),
    .Y(_10990_));
 sky130_fd_sc_hd__nand2_1 _31605_ (.A(net1241),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[4] ),
    .Y(_10991_));
 sky130_fd_sc_hd__nand2_1 _31606_ (.A(net1872),
    .B(\inst$top.soc.cpu.exception.w_data$48[4] ),
    .Y(_10992_));
 sky130_fd_sc_hd__a31oi_1 _31607_ (.A1(_10990_),
    .A2(_10991_),
    .A3(_10992_),
    .B1(net2936),
    .Y(_03808_));
 sky130_fd_sc_hd__nand2_1 _31608_ (.A(net1098),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[5] ),
    .Y(_10993_));
 sky130_fd_sc_hd__nand2_1 _31609_ (.A(net1243),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[5] ),
    .Y(_10994_));
 sky130_fd_sc_hd__a21oi_1 _31610_ (.A1(_10993_),
    .A2(_10994_),
    .B1(net2939),
    .Y(_03809_));
 sky130_fd_sc_hd__nand2_1 _31611_ (.A(net1096),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[6] ),
    .Y(_10995_));
 sky130_fd_sc_hd__nand2_1 _31612_ (.A(net1241),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[6] ),
    .Y(_10996_));
 sky130_fd_sc_hd__a21oi_1 _31613_ (.A1(_10995_),
    .A2(_10996_),
    .B1(net2939),
    .Y(_03810_));
 sky130_fd_sc_hd__nand2_1 _31614_ (.A(net1096),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[7] ),
    .Y(_10997_));
 sky130_fd_sc_hd__nand2_1 _31615_ (.A(net1241),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[7] ),
    .Y(_10998_));
 sky130_fd_sc_hd__a21oi_1 _31616_ (.A1(_10997_),
    .A2(_10998_),
    .B1(net2937),
    .Y(_03811_));
 sky130_fd_sc_hd__nand2_1 _31617_ (.A(net1097),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[8] ),
    .Y(_10999_));
 sky130_fd_sc_hd__nand2_1 _31618_ (.A(net1242),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[8] ),
    .Y(_11000_));
 sky130_fd_sc_hd__a21oi_1 _31619_ (.A1(_10999_),
    .A2(_11000_),
    .B1(net2942),
    .Y(_03812_));
 sky130_fd_sc_hd__nand2_1 _31620_ (.A(net1098),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[9] ),
    .Y(_11001_));
 sky130_fd_sc_hd__nand2_1 _31621_ (.A(net1243),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[9] ),
    .Y(_11002_));
 sky130_fd_sc_hd__a21oi_1 _31622_ (.A1(_11001_),
    .A2(_11002_),
    .B1(net2941),
    .Y(_03813_));
 sky130_fd_sc_hd__nor2_1 _31625_ (.A(net2912),
    .B(net1883),
    .Y(_11005_));
 sky130_fd_sc_hd__o21ai_0 _31628_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause_m_select ),
    .A2(net2216),
    .B1(net2031),
    .Y(_11008_));
 sky130_fd_sc_hd__nor2_1 _31629_ (.A(_11005_),
    .B(_11008_),
    .Y(_03814_));
 sky130_fd_sc_hd__nor2_1 _31630_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause_m_select ),
    .B(net1883),
    .Y(_11009_));
 sky130_fd_sc_hd__o21ai_0 _31632_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause_w_select ),
    .A2(net2220),
    .B1(net2031),
    .Y(_11011_));
 sky130_fd_sc_hd__nor2_1 _31633_ (.A(_11009_),
    .B(_11011_),
    .Y(_03815_));
 sky130_fd_sc_hd__nor2_1 _31634_ (.A(net2912),
    .B(net672),
    .Y(_11012_));
 sky130_fd_sc_hd__nand2_1 _31635_ (.A(_06037_),
    .B(\inst$top.soc.cpu.sink__payload$6[40] ),
    .Y(_11013_));
 sky130_fd_sc_hd__o21ai_4 _31636_ (.A1(_20261_),
    .A2(_06041_),
    .B1(_11013_),
    .Y(_11014_));
 sky130_fd_sc_hd__inv_1 _31637_ (.A(_11014_),
    .Y(_11015_));
 sky130_fd_sc_hd__a22oi_1 _31638_ (.A1(\inst$top.soc.cpu.sink__payload$6[39] ),
    .A2(_09363_),
    .B1(_09360_),
    .B2(net2687),
    .Y(_11016_));
 sky130_fd_sc_hd__inv_1 _31639_ (.A(net1031),
    .Y(_11017_));
 sky130_fd_sc_hd__nor2_1 _31640_ (.A(_06044_),
    .B(net884),
    .Y(_11018_));
 sky130_fd_sc_hd__inv_1 _31641_ (.A(_11018_),
    .Y(_11019_));
 sky130_fd_sc_hd__inv_1 _31642_ (.A(\inst$top.soc.cpu.csrf.d_addr[6] ),
    .Y(_11020_));
 sky130_fd_sc_hd__or2_2 _31643_ (.A(\inst$top.soc.cpu.csrf.d_addr[5] ),
    .B(\inst$top.soc.cpu.csrf.d_addr[4] ),
    .X(_11021_));
 sky130_fd_sc_hd__nor2_1 _31644_ (.A(_11020_),
    .B(_11021_),
    .Y(_11022_));
 sky130_fd_sc_hd__inv_1 _31645_ (.A(_11022_),
    .Y(_11023_));
 sky130_fd_sc_hd__nor4_1 _31646_ (.A(_11015_),
    .B(_11017_),
    .C(_11019_),
    .D(_11023_),
    .Y(_11024_));
 sky130_fd_sc_hd__o21ai_1 _31649_ (.A1(_11024_),
    .A2(net633),
    .B1(net2033),
    .Y(_11027_));
 sky130_fd_sc_hd__nor2_4 _31650_ (.A(_11012_),
    .B(_11027_),
    .Y(_03816_));
 sky130_fd_sc_hd__nand2_1 _31651_ (.A(net1807),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc_w_select ),
    .Y(_11028_));
 sky130_fd_sc_hd__nand2_1 _31652_ (.A(_11028_),
    .B(_10913_),
    .Y(_11029_));
 sky130_fd_sc_hd__inv_1 _31653_ (.A(_11029_),
    .Y(_11030_));
 sky130_fd_sc_hd__nand2_1 _31655_ (.A(net1092),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[0] ),
    .Y(_11032_));
 sky130_fd_sc_hd__inv_1 _31656_ (.A(_11028_),
    .Y(_11033_));
 sky130_fd_sc_hd__nand2_1 _31658_ (.A(net1237),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[2] ),
    .Y(_11035_));
 sky130_fd_sc_hd__nand2_1 _31659_ (.A(net1872),
    .B(\inst$top.soc.cpu.sink__payload$24[2] ),
    .Y(_11036_));
 sky130_fd_sc_hd__a31oi_1 _31660_ (.A1(_11032_),
    .A2(_11035_),
    .A3(_11036_),
    .B1(net2936),
    .Y(_03817_));
 sky130_fd_sc_hd__nand2_1 _31661_ (.A(net1094),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[10] ),
    .Y(_11037_));
 sky130_fd_sc_hd__nand2_1 _31662_ (.A(net1239),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[12] ),
    .Y(_11038_));
 sky130_fd_sc_hd__nand2_1 _31663_ (.A(net1876),
    .B(\inst$top.soc.cpu.sink__payload$24[12] ),
    .Y(_11039_));
 sky130_fd_sc_hd__a31oi_1 _31664_ (.A1(_11037_),
    .A2(_11038_),
    .A3(_11039_),
    .B1(net2941),
    .Y(_03818_));
 sky130_fd_sc_hd__nand2_1 _31665_ (.A(net1093),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[11] ),
    .Y(_11040_));
 sky130_fd_sc_hd__nand2_1 _31666_ (.A(net1238),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[13] ),
    .Y(_11041_));
 sky130_fd_sc_hd__nand2_1 _31667_ (.A(net1879),
    .B(\inst$top.soc.cpu.sink__payload$24[13] ),
    .Y(_11042_));
 sky130_fd_sc_hd__a31oi_1 _31668_ (.A1(_11040_),
    .A2(_11041_),
    .A3(_11042_),
    .B1(net2968),
    .Y(_03819_));
 sky130_fd_sc_hd__nand2_1 _31669_ (.A(net1093),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[12] ),
    .Y(_11043_));
 sky130_fd_sc_hd__nand2_1 _31670_ (.A(net1238),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[14] ),
    .Y(_11044_));
 sky130_fd_sc_hd__nand2_1 _31671_ (.A(net1879),
    .B(\inst$top.soc.cpu.sink__payload$24[14] ),
    .Y(_11045_));
 sky130_fd_sc_hd__a31oi_1 _31672_ (.A1(_11043_),
    .A2(_11044_),
    .A3(_11045_),
    .B1(net2952),
    .Y(_03820_));
 sky130_fd_sc_hd__nand2_1 _31673_ (.A(net1093),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[13] ),
    .Y(_11046_));
 sky130_fd_sc_hd__nand2_1 _31674_ (.A(net1238),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[15] ),
    .Y(_11047_));
 sky130_fd_sc_hd__nand2_1 _31676_ (.A(net1879),
    .B(\inst$top.soc.cpu.sink__payload$24[15] ),
    .Y(_11049_));
 sky130_fd_sc_hd__a31oi_1 _31677_ (.A1(_11046_),
    .A2(_11047_),
    .A3(_11049_),
    .B1(net2952),
    .Y(_03821_));
 sky130_fd_sc_hd__nand2_1 _31678_ (.A(net1092),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[14] ),
    .Y(_11050_));
 sky130_fd_sc_hd__nand2_1 _31679_ (.A(net1237),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[16] ),
    .Y(_11051_));
 sky130_fd_sc_hd__nand2_1 _31680_ (.A(net1875),
    .B(\inst$top.soc.cpu.sink__payload$24[16] ),
    .Y(_11052_));
 sky130_fd_sc_hd__a31oi_1 _31681_ (.A1(_11050_),
    .A2(_11051_),
    .A3(_11052_),
    .B1(net2961),
    .Y(_03822_));
 sky130_fd_sc_hd__nand2_1 _31682_ (.A(net1094),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[15] ),
    .Y(_11053_));
 sky130_fd_sc_hd__nand2_1 _31683_ (.A(net1239),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[17] ),
    .Y(_11054_));
 sky130_fd_sc_hd__nand2_1 _31684_ (.A(net1876),
    .B(\inst$top.soc.cpu.sink__payload$24[17] ),
    .Y(_11055_));
 sky130_fd_sc_hd__a31oi_1 _31686_ (.A1(_11053_),
    .A2(_11054_),
    .A3(_11055_),
    .B1(net2962),
    .Y(_03823_));
 sky130_fd_sc_hd__nand2_1 _31687_ (.A(net1092),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[16] ),
    .Y(_11057_));
 sky130_fd_sc_hd__nand2_1 _31688_ (.A(net1237),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[18] ),
    .Y(_11058_));
 sky130_fd_sc_hd__nand2_1 _31689_ (.A(net1875),
    .B(\inst$top.soc.cpu.sink__payload$24[18] ),
    .Y(_11059_));
 sky130_fd_sc_hd__a31oi_1 _31690_ (.A1(_11057_),
    .A2(_11058_),
    .A3(_11059_),
    .B1(net2963),
    .Y(_03824_));
 sky130_fd_sc_hd__nand2_1 _31691_ (.A(net1092),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[17] ),
    .Y(_11060_));
 sky130_fd_sc_hd__nand2_1 _31692_ (.A(net1237),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[19] ),
    .Y(_11061_));
 sky130_fd_sc_hd__nand2_1 _31693_ (.A(net1876),
    .B(\inst$top.soc.cpu.sink__payload$24[19] ),
    .Y(_11062_));
 sky130_fd_sc_hd__a31oi_1 _31694_ (.A1(_11060_),
    .A2(_11061_),
    .A3(_11062_),
    .B1(net2963),
    .Y(_03825_));
 sky130_fd_sc_hd__nand2_1 _31695_ (.A(net1092),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[18] ),
    .Y(_11063_));
 sky130_fd_sc_hd__nand2_1 _31696_ (.A(net1237),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[20] ),
    .Y(_11064_));
 sky130_fd_sc_hd__nand2_1 _31697_ (.A(net1875),
    .B(\inst$top.soc.cpu.sink__payload$24[20] ),
    .Y(_11065_));
 sky130_fd_sc_hd__a31oi_1 _31698_ (.A1(_11063_),
    .A2(_11064_),
    .A3(_11065_),
    .B1(net2961),
    .Y(_03826_));
 sky130_fd_sc_hd__nand2_1 _31700_ (.A(net1095),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[19] ),
    .Y(_11067_));
 sky130_fd_sc_hd__nand2_1 _31702_ (.A(net1240),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[21] ),
    .Y(_11069_));
 sky130_fd_sc_hd__nand2_1 _31703_ (.A(net1874),
    .B(\inst$top.soc.cpu.sink__payload$24[21] ),
    .Y(_11070_));
 sky130_fd_sc_hd__a31oi_1 _31704_ (.A1(_11067_),
    .A2(_11069_),
    .A3(_11070_),
    .B1(net2961),
    .Y(_03827_));
 sky130_fd_sc_hd__nand2_1 _31705_ (.A(net1092),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[1] ),
    .Y(_11071_));
 sky130_fd_sc_hd__nand2_1 _31706_ (.A(net1237),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[3] ),
    .Y(_11072_));
 sky130_fd_sc_hd__nand2_1 _31707_ (.A(net1873),
    .B(\inst$top.soc.cpu.sink__payload$24[3] ),
    .Y(_11073_));
 sky130_fd_sc_hd__a31oi_1 _31708_ (.A1(_11071_),
    .A2(_11072_),
    .A3(_11073_),
    .B1(net2958),
    .Y(_03828_));
 sky130_fd_sc_hd__nand2_1 _31709_ (.A(net1094),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[20] ),
    .Y(_11074_));
 sky130_fd_sc_hd__nand2_1 _31710_ (.A(net1239),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[22] ),
    .Y(_11075_));
 sky130_fd_sc_hd__nand2_1 _31711_ (.A(net1877),
    .B(\inst$top.soc.cpu.sink__payload$24[22] ),
    .Y(_11076_));
 sky130_fd_sc_hd__a31oi_1 _31712_ (.A1(_11074_),
    .A2(_11075_),
    .A3(_11076_),
    .B1(net2969),
    .Y(_03829_));
 sky130_fd_sc_hd__nand2_1 _31713_ (.A(net1094),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[21] ),
    .Y(_11077_));
 sky130_fd_sc_hd__nand2_1 _31714_ (.A(net1239),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[23] ),
    .Y(_11078_));
 sky130_fd_sc_hd__nand2_1 _31715_ (.A(net1877),
    .B(\inst$top.soc.cpu.sink__payload$24[23] ),
    .Y(_11079_));
 sky130_fd_sc_hd__a31oi_1 _31716_ (.A1(_11077_),
    .A2(_11078_),
    .A3(_11079_),
    .B1(net2971),
    .Y(_03830_));
 sky130_fd_sc_hd__nand2_1 _31717_ (.A(net1093),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[22] ),
    .Y(_11080_));
 sky130_fd_sc_hd__nand2_1 _31718_ (.A(net1238),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[24] ),
    .Y(_11081_));
 sky130_fd_sc_hd__nand2_1 _31720_ (.A(net1877),
    .B(\inst$top.soc.cpu.sink__payload$24[24] ),
    .Y(_11083_));
 sky130_fd_sc_hd__a31oi_1 _31721_ (.A1(_11080_),
    .A2(_11081_),
    .A3(_11083_),
    .B1(net2970),
    .Y(_03831_));
 sky130_fd_sc_hd__nand2_1 _31722_ (.A(net1092),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[23] ),
    .Y(_11084_));
 sky130_fd_sc_hd__nand2_1 _31723_ (.A(net1237),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[25] ),
    .Y(_11085_));
 sky130_fd_sc_hd__nand2_1 _31724_ (.A(net1873),
    .B(\inst$top.soc.cpu.sink__payload$24[25] ),
    .Y(_11086_));
 sky130_fd_sc_hd__a31oi_1 _31725_ (.A1(_11084_),
    .A2(_11085_),
    .A3(_11086_),
    .B1(net2957),
    .Y(_03832_));
 sky130_fd_sc_hd__nand2_1 _31726_ (.A(net1093),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[24] ),
    .Y(_11087_));
 sky130_fd_sc_hd__nand2_1 _31727_ (.A(net1238),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[26] ),
    .Y(_11088_));
 sky130_fd_sc_hd__nand2_1 _31728_ (.A(net1877),
    .B(\inst$top.soc.cpu.sink__payload$24[26] ),
    .Y(_11089_));
 sky130_fd_sc_hd__a31oi_1 _31730_ (.A1(_11087_),
    .A2(_11088_),
    .A3(_11089_),
    .B1(net2973),
    .Y(_03833_));
 sky130_fd_sc_hd__nand2_1 _31731_ (.A(net1093),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[25] ),
    .Y(_11091_));
 sky130_fd_sc_hd__nand2_1 _31732_ (.A(net1238),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[27] ),
    .Y(_11092_));
 sky130_fd_sc_hd__nand2_1 _31733_ (.A(net1877),
    .B(\inst$top.soc.cpu.sink__payload$24[27] ),
    .Y(_11093_));
 sky130_fd_sc_hd__a31oi_1 _31734_ (.A1(_11091_),
    .A2(_11092_),
    .A3(_11093_),
    .B1(net2970),
    .Y(_03834_));
 sky130_fd_sc_hd__nand2_1 _31735_ (.A(net1093),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[26] ),
    .Y(_11094_));
 sky130_fd_sc_hd__nand2_1 _31736_ (.A(net1238),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[28] ),
    .Y(_11095_));
 sky130_fd_sc_hd__nand2_1 _31737_ (.A(net1877),
    .B(\inst$top.soc.cpu.sink__payload$24[28] ),
    .Y(_11096_));
 sky130_fd_sc_hd__a31oi_1 _31738_ (.A1(_11094_),
    .A2(_11095_),
    .A3(_11096_),
    .B1(net2970),
    .Y(_03835_));
 sky130_fd_sc_hd__nand2_1 _31739_ (.A(net1093),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[27] ),
    .Y(_11097_));
 sky130_fd_sc_hd__nand2_1 _31740_ (.A(net1238),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[29] ),
    .Y(_11098_));
 sky130_fd_sc_hd__nand2_1 _31741_ (.A(net1877),
    .B(\inst$top.soc.cpu.sink__payload$24[29] ),
    .Y(_11099_));
 sky130_fd_sc_hd__a31oi_1 _31742_ (.A1(_11097_),
    .A2(_11098_),
    .A3(_11099_),
    .B1(net2970),
    .Y(_03836_));
 sky130_fd_sc_hd__nand2_1 _31744_ (.A(net1093),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[28] ),
    .Y(_11101_));
 sky130_fd_sc_hd__nand2_1 _31746_ (.A(net1238),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[30] ),
    .Y(_11103_));
 sky130_fd_sc_hd__nand2_1 _31747_ (.A(net1879),
    .B(\inst$top.soc.cpu.sink__payload$24[30] ),
    .Y(_11104_));
 sky130_fd_sc_hd__a31oi_1 _31748_ (.A1(_11101_),
    .A2(_11103_),
    .A3(_11104_),
    .B1(net2970),
    .Y(_03837_));
 sky130_fd_sc_hd__nand2_1 _31749_ (.A(net1092),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[29] ),
    .Y(_11105_));
 sky130_fd_sc_hd__nand2_1 _31750_ (.A(net1237),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[31] ),
    .Y(_11106_));
 sky130_fd_sc_hd__nand2_1 _31751_ (.A(net1872),
    .B(\inst$top.soc.cpu.sink__payload$24[31] ),
    .Y(_11107_));
 sky130_fd_sc_hd__a31oi_1 _31752_ (.A1(_11105_),
    .A2(_11106_),
    .A3(_11107_),
    .B1(net2937),
    .Y(_03838_));
 sky130_fd_sc_hd__nand2_1 _31753_ (.A(net1092),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[2] ),
    .Y(_11108_));
 sky130_fd_sc_hd__nand2_1 _31754_ (.A(net1237),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[4] ),
    .Y(_11109_));
 sky130_fd_sc_hd__nand2_1 _31755_ (.A(net1872),
    .B(\inst$top.soc.cpu.sink__payload$24[4] ),
    .Y(_11110_));
 sky130_fd_sc_hd__a31oi_1 _31756_ (.A1(_11108_),
    .A2(_11109_),
    .A3(_11110_),
    .B1(net2937),
    .Y(_03839_));
 sky130_fd_sc_hd__nand2_1 _31757_ (.A(net1095),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[3] ),
    .Y(_11111_));
 sky130_fd_sc_hd__nand2_1 _31758_ (.A(net1240),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[5] ),
    .Y(_11112_));
 sky130_fd_sc_hd__nand2_1 _31759_ (.A(net1874),
    .B(\inst$top.soc.cpu.sink__payload$24[5] ),
    .Y(_11113_));
 sky130_fd_sc_hd__a31oi_1 _31760_ (.A1(_11111_),
    .A2(_11112_),
    .A3(_11113_),
    .B1(net2939),
    .Y(_03840_));
 sky130_fd_sc_hd__nand2_1 _31761_ (.A(net1095),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[4] ),
    .Y(_11114_));
 sky130_fd_sc_hd__nand2_1 _31762_ (.A(net1240),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[6] ),
    .Y(_11115_));
 sky130_fd_sc_hd__nand2_1 _31764_ (.A(net1874),
    .B(\inst$top.soc.cpu.sink__payload$24[6] ),
    .Y(_11117_));
 sky130_fd_sc_hd__a31oi_1 _31765_ (.A1(_11114_),
    .A2(_11115_),
    .A3(_11117_),
    .B1(net2940),
    .Y(_03841_));
 sky130_fd_sc_hd__nand2_1 _31766_ (.A(net1092),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[5] ),
    .Y(_11118_));
 sky130_fd_sc_hd__nand2_1 _31767_ (.A(net1237),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[7] ),
    .Y(_11119_));
 sky130_fd_sc_hd__nand2_1 _31768_ (.A(net1872),
    .B(\inst$top.soc.cpu.sink__payload$24[7] ),
    .Y(_11120_));
 sky130_fd_sc_hd__a31oi_1 _31769_ (.A1(_11118_),
    .A2(_11119_),
    .A3(_11120_),
    .B1(net2937),
    .Y(_03842_));
 sky130_fd_sc_hd__nand2_1 _31770_ (.A(net1094),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[6] ),
    .Y(_11121_));
 sky130_fd_sc_hd__nand2_1 _31771_ (.A(net1239),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[8] ),
    .Y(_11122_));
 sky130_fd_sc_hd__nand2_1 _31772_ (.A(net1876),
    .B(\inst$top.soc.cpu.sink__payload$24[8] ),
    .Y(_11123_));
 sky130_fd_sc_hd__a31oi_1 _31774_ (.A1(_11121_),
    .A2(_11122_),
    .A3(_11123_),
    .B1(net2941),
    .Y(_03843_));
 sky130_fd_sc_hd__nand2_1 _31775_ (.A(net1094),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[7] ),
    .Y(_11125_));
 sky130_fd_sc_hd__nand2_1 _31776_ (.A(net1239),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[9] ),
    .Y(_11126_));
 sky130_fd_sc_hd__nand2_1 _31777_ (.A(net1876),
    .B(\inst$top.soc.cpu.sink__payload$24[9] ),
    .Y(_11127_));
 sky130_fd_sc_hd__a31oi_1 _31778_ (.A1(_11125_),
    .A2(_11126_),
    .A3(_11127_),
    .B1(net2941),
    .Y(_03844_));
 sky130_fd_sc_hd__nand2_1 _31779_ (.A(net1093),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[8] ),
    .Y(_11128_));
 sky130_fd_sc_hd__nand2_1 _31780_ (.A(net1238),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[10] ),
    .Y(_11129_));
 sky130_fd_sc_hd__nand2_1 _31781_ (.A(net1879),
    .B(\inst$top.soc.cpu.sink__payload$24[10] ),
    .Y(_11130_));
 sky130_fd_sc_hd__a31oi_1 _31782_ (.A1(_11128_),
    .A2(_11129_),
    .A3(_11130_),
    .B1(net2953),
    .Y(_03845_));
 sky130_fd_sc_hd__nand2_1 _31783_ (.A(net1095),
    .B(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[9] ),
    .Y(_11131_));
 sky130_fd_sc_hd__nand2_1 _31784_ (.A(net1240),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[11] ),
    .Y(_11132_));
 sky130_fd_sc_hd__nand2_1 _31785_ (.A(net1874),
    .B(\inst$top.soc.cpu.sink__payload$24[11] ),
    .Y(_11133_));
 sky130_fd_sc_hd__a31oi_1 _31786_ (.A1(_11131_),
    .A2(_11132_),
    .A3(_11133_),
    .B1(net2961),
    .Y(_03846_));
 sky130_fd_sc_hd__nor2_1 _31788_ (.A(net2908),
    .B(net1883),
    .Y(_11135_));
 sky130_fd_sc_hd__o21ai_0 _31790_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mepc_m_select ),
    .A2(net2220),
    .B1(net2083),
    .Y(_11137_));
 sky130_fd_sc_hd__nor2_1 _31791_ (.A(_11135_),
    .B(_11137_),
    .Y(_03847_));
 sky130_fd_sc_hd__nor2_1 _31792_ (.A(\inst$top.soc.cpu.exception.csr_bank.mepc_m_select ),
    .B(net1883),
    .Y(_11138_));
 sky130_fd_sc_hd__o21ai_0 _31793_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mepc_w_select ),
    .A2(net2220),
    .B1(net2083),
    .Y(_11139_));
 sky130_fd_sc_hd__nor2_1 _31794_ (.A(_11138_),
    .B(_11139_),
    .Y(_03848_));
 sky130_fd_sc_hd__nor2_1 _31795_ (.A(net2908),
    .B(net672),
    .Y(_11140_));
 sky130_fd_sc_hd__nor2_1 _31796_ (.A(net1031),
    .B(_11014_),
    .Y(_11141_));
 sky130_fd_sc_hd__nand2_1 _31797_ (.A(_11018_),
    .B(_11141_),
    .Y(_11142_));
 sky130_fd_sc_hd__nor2_1 _31798_ (.A(_11142_),
    .B(_11023_),
    .Y(_11143_));
 sky130_fd_sc_hd__o21ai_1 _31799_ (.A1(_11143_),
    .A2(net633),
    .B1(net2033),
    .Y(_11144_));
 sky130_fd_sc_hd__nor2_4 _31800_ (.A(_11140_),
    .B(_11144_),
    .Y(_03849_));
 sky130_fd_sc_hd__nand2_1 _31801_ (.A(net1807),
    .B(\inst$top.soc.cpu.exception.csr_bank.mie_w_select ),
    .Y(_11145_));
 sky130_fd_sc_hd__nand2_1 _31803_ (.A(net1663),
    .B(\inst$top.soc.cpu.exception.csr_bank.mie.meie.x_data ),
    .Y(_11147_));
 sky130_fd_sc_hd__nand3_1 _31806_ (.A(net1808),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[11] ),
    .C(\inst$top.soc.cpu.exception.csr_bank.mie_w_select ),
    .Y(_11150_));
 sky130_fd_sc_hd__a21oi_1 _31807_ (.A1(_11147_),
    .A2(_11150_),
    .B1(net2957),
    .Y(_03850_));
 sky130_fd_sc_hd__nand2_1 _31808_ (.A(net1663),
    .B(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[0] ),
    .Y(_11151_));
 sky130_fd_sc_hd__nand3_1 _31810_ (.A(net1809),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[16] ),
    .C(\inst$top.soc.cpu.exception.csr_bank.mie_w_select ),
    .Y(_11153_));
 sky130_fd_sc_hd__a21oi_1 _31811_ (.A1(_11151_),
    .A2(_11153_),
    .B1(net2957),
    .Y(_03851_));
 sky130_fd_sc_hd__o21ai_0 _31813_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[26] ),
    .A2(net1661),
    .B1(net2099),
    .Y(_11155_));
 sky130_fd_sc_hd__a21oi_1 _31814_ (.A1(_05815_),
    .A2(net1661),
    .B1(_11155_),
    .Y(_03852_));
 sky130_fd_sc_hd__o21ai_0 _31816_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[27] ),
    .A2(net1660),
    .B1(net2095),
    .Y(_11157_));
 sky130_fd_sc_hd__a21oi_1 _31817_ (.A1(_05828_),
    .A2(net1660),
    .B1(_11157_),
    .Y(_03853_));
 sky130_fd_sc_hd__o21ai_0 _31818_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[28] ),
    .A2(net1660),
    .B1(net2095),
    .Y(_11158_));
 sky130_fd_sc_hd__a21oi_1 _31819_ (.A1(_05841_),
    .A2(net1660),
    .B1(_11158_),
    .Y(_03854_));
 sky130_fd_sc_hd__o21ai_0 _31820_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[29] ),
    .A2(net1660),
    .B1(net2095),
    .Y(_11159_));
 sky130_fd_sc_hd__a21oi_1 _31821_ (.A1(_05854_),
    .A2(net1660),
    .B1(_11159_),
    .Y(_03855_));
 sky130_fd_sc_hd__o21ai_0 _31823_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[30] ),
    .A2(net1660),
    .B1(net2095),
    .Y(_11161_));
 sky130_fd_sc_hd__a21oi_1 _31824_ (.A1(_05863_),
    .A2(net1660),
    .B1(_11161_),
    .Y(_03856_));
 sky130_fd_sc_hd__nand2_1 _31825_ (.A(net1663),
    .B(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[15] ),
    .Y(_11162_));
 sky130_fd_sc_hd__nand3_1 _31826_ (.A(net1809),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[31] ),
    .C(\inst$top.soc.cpu.exception.csr_bank.mie_w_select ),
    .Y(_11163_));
 sky130_fd_sc_hd__a21oi_1 _31827_ (.A1(_11162_),
    .A2(_11163_),
    .B1(net2957),
    .Y(_03857_));
 sky130_fd_sc_hd__o21ai_0 _31828_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[17] ),
    .A2(net1662),
    .B1(net2098),
    .Y(_11164_));
 sky130_fd_sc_hd__a21oi_1 _31829_ (.A1(_05631_),
    .A2(net1662),
    .B1(_11164_),
    .Y(_03858_));
 sky130_fd_sc_hd__o21ai_0 _31830_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[18] ),
    .A2(net1662),
    .B1(net2098),
    .Y(_11165_));
 sky130_fd_sc_hd__a21oi_1 _31831_ (.A1(_05652_),
    .A2(net1662),
    .B1(_11165_),
    .Y(_03859_));
 sky130_fd_sc_hd__o21ai_0 _31832_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[19] ),
    .A2(net1662),
    .B1(net2098),
    .Y(_11166_));
 sky130_fd_sc_hd__a21oi_1 _31833_ (.A1(_05674_),
    .A2(net1662),
    .B1(_11166_),
    .Y(_03860_));
 sky130_fd_sc_hd__o21ai_0 _31834_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[20] ),
    .A2(net1663),
    .B1(net2090),
    .Y(_11167_));
 sky130_fd_sc_hd__a21oi_1 _31835_ (.A1(_05699_),
    .A2(net1663),
    .B1(_11167_),
    .Y(_03861_));
 sky130_fd_sc_hd__o21ai_0 _31836_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[21] ),
    .A2(net1662),
    .B1(net2094),
    .Y(_11168_));
 sky130_fd_sc_hd__a21oi_1 _31837_ (.A1(_05720_),
    .A2(net1662),
    .B1(_11168_),
    .Y(_03862_));
 sky130_fd_sc_hd__o21ai_0 _31838_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[22] ),
    .A2(net1661),
    .B1(net2099),
    .Y(_11169_));
 sky130_fd_sc_hd__a21oi_1 _31839_ (.A1(_05738_),
    .A2(net1661),
    .B1(_11169_),
    .Y(_03863_));
 sky130_fd_sc_hd__o21ai_0 _31840_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[23] ),
    .A2(net1661),
    .B1(net2099),
    .Y(_11170_));
 sky130_fd_sc_hd__a21oi_1 _31841_ (.A1(_05759_),
    .A2(net1661),
    .B1(_11170_),
    .Y(_03864_));
 sky130_fd_sc_hd__o21ai_0 _31842_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[24] ),
    .A2(net1660),
    .B1(net2096),
    .Y(_11171_));
 sky130_fd_sc_hd__a21oi_1 _31843_ (.A1(_05776_),
    .A2(net1660),
    .B1(_11171_),
    .Y(_03865_));
 sky130_fd_sc_hd__o21ai_0 _31844_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[25] ),
    .A2(net1663),
    .B1(net2092),
    .Y(_11172_));
 sky130_fd_sc_hd__a21oi_1 _31845_ (.A1(_05796_),
    .A2(net1663),
    .B1(_11172_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand2_1 _31846_ (.A(net1663),
    .B(\inst$top.soc.cpu.exception.csr_bank.mie.msie.x_data ),
    .Y(_11173_));
 sky130_fd_sc_hd__nand3_1 _31847_ (.A(net1808),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[3] ),
    .C(\inst$top.soc.cpu.exception.csr_bank.mie_w_select ),
    .Y(_11174_));
 sky130_fd_sc_hd__a21oi_1 _31848_ (.A1(_11173_),
    .A2(_11174_),
    .B1(net2957),
    .Y(_03867_));
 sky130_fd_sc_hd__nand2_1 _31849_ (.A(net1663),
    .B(\inst$top.soc.cpu.exception.csr_bank.mie.mtie.x_data ),
    .Y(_11175_));
 sky130_fd_sc_hd__nand3_1 _31850_ (.A(net1808),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[7] ),
    .C(\inst$top.soc.cpu.exception.csr_bank.mie_w_select ),
    .Y(_11176_));
 sky130_fd_sc_hd__a21oi_1 _31852_ (.A1(_11175_),
    .A2(_11176_),
    .B1(net2957),
    .Y(_03868_));
 sky130_fd_sc_hd__o21ai_0 _31854_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mie_m_select ),
    .A2(net2222),
    .B1(net2085),
    .Y(_11179_));
 sky130_fd_sc_hd__a21oi_1 _31855_ (.A1(net2195),
    .A2(net2221),
    .B1(_11179_),
    .Y(_03869_));
 sky130_fd_sc_hd__nor2_1 _31856_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie_m_select ),
    .B(net1884),
    .Y(_11180_));
 sky130_fd_sc_hd__o21ai_0 _31857_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mie_w_select ),
    .A2(net2221),
    .B1(net2085),
    .Y(_11181_));
 sky130_fd_sc_hd__nor2_1 _31858_ (.A(_11180_),
    .B(_11181_),
    .Y(_03870_));
 sky130_fd_sc_hd__nor2_1 _31859_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie_x_select ),
    .B(net671),
    .Y(_11182_));
 sky130_fd_sc_hd__inv_1 _31861_ (.A(_06044_),
    .Y(_11184_));
 sky130_fd_sc_hd__nor4_1 _31862_ (.A(_11017_),
    .B(_11014_),
    .C(net884),
    .D(_11184_),
    .Y(_11185_));
 sky130_fd_sc_hd__nor2_1 _31863_ (.A(\inst$top.soc.cpu.csrf.d_addr[6] ),
    .B(_11021_),
    .Y(_11186_));
 sky130_fd_sc_hd__nand2_1 _31864_ (.A(_11185_),
    .B(_11186_),
    .Y(_11187_));
 sky130_fd_sc_hd__nand2_1 _31865_ (.A(net671),
    .B(_11187_),
    .Y(_11188_));
 sky130_fd_sc_hd__nand2_1 _31867_ (.A(_11188_),
    .B(net2031),
    .Y(_11190_));
 sky130_fd_sc_hd__nor2_4 _31868_ (.A(_11182_),
    .B(_11190_),
    .Y(_03871_));
 sky130_fd_sc_hd__nand3_1 _31871_ (.A(net1808),
    .B(net2906),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[11] ),
    .Y(_11193_));
 sky130_fd_sc_hd__clkinv_1 _31872_ (.A(\inst$top.soc.cpu.m.source__valid ),
    .Y(_11194_));
 sky130_fd_sc_hd__nand2_1 _31874_ (.A(net2021),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.meip.x_data ),
    .Y(_11196_));
 sky130_fd_sc_hd__a21oi_1 _31875_ (.A1(_11193_),
    .A2(_11196_),
    .B1(net2958),
    .Y(_03872_));
 sky130_fd_sc_hd__nand3_1 _31876_ (.A(net1809),
    .B(net2906),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[16] ),
    .Y(_11197_));
 sky130_fd_sc_hd__nand2_1 _31877_ (.A(net2021),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[0] ),
    .Y(_11198_));
 sky130_fd_sc_hd__a21oi_1 _31878_ (.A1(_11197_),
    .A2(_11198_),
    .B1(net2959),
    .Y(_03873_));
 sky130_fd_sc_hd__nand3_1 _31879_ (.A(net1812),
    .B(net2907),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[26] ),
    .Y(_11199_));
 sky130_fd_sc_hd__nand2_1 _31880_ (.A(net2022),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[10] ),
    .Y(_11200_));
 sky130_fd_sc_hd__a21oi_1 _31881_ (.A1(_11199_),
    .A2(_11200_),
    .B1(net2964),
    .Y(_03874_));
 sky130_fd_sc_hd__nand3_1 _31882_ (.A(net1812),
    .B(net2907),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[27] ),
    .Y(_11201_));
 sky130_fd_sc_hd__nand2_1 _31883_ (.A(net2022),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[11] ),
    .Y(_11202_));
 sky130_fd_sc_hd__a21oi_1 _31884_ (.A1(_11201_),
    .A2(_11202_),
    .B1(net2962),
    .Y(_03875_));
 sky130_fd_sc_hd__nand3_1 _31885_ (.A(net1812),
    .B(net2907),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[28] ),
    .Y(_11203_));
 sky130_fd_sc_hd__nand2_1 _31886_ (.A(net2022),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[12] ),
    .Y(_11204_));
 sky130_fd_sc_hd__a21oi_1 _31887_ (.A1(_11203_),
    .A2(_11204_),
    .B1(net2962),
    .Y(_03876_));
 sky130_fd_sc_hd__nand3_1 _31888_ (.A(net1814),
    .B(net2907),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[29] ),
    .Y(_11205_));
 sky130_fd_sc_hd__nand2_1 _31889_ (.A(net2022),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[13] ),
    .Y(_11206_));
 sky130_fd_sc_hd__a21oi_1 _31890_ (.A1(_11205_),
    .A2(_11206_),
    .B1(net2962),
    .Y(_03877_));
 sky130_fd_sc_hd__nand3_1 _31891_ (.A(net1811),
    .B(net2907),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[30] ),
    .Y(_11207_));
 sky130_fd_sc_hd__nand2_1 _31892_ (.A(net2022),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[14] ),
    .Y(_11208_));
 sky130_fd_sc_hd__a21oi_1 _31893_ (.A1(_11207_),
    .A2(_11208_),
    .B1(net2962),
    .Y(_03878_));
 sky130_fd_sc_hd__nand3_1 _31894_ (.A(net1809),
    .B(net2906),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[31] ),
    .Y(_11209_));
 sky130_fd_sc_hd__nand2_1 _31895_ (.A(net2021),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[15] ),
    .Y(_11210_));
 sky130_fd_sc_hd__a21oi_1 _31896_ (.A1(_11209_),
    .A2(_11210_),
    .B1(net2959),
    .Y(_03879_));
 sky130_fd_sc_hd__nand3_1 _31897_ (.A(net1813),
    .B(net2907),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[17] ),
    .Y(_11211_));
 sky130_fd_sc_hd__nand2_1 _31898_ (.A(net2022),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[1] ),
    .Y(_11212_));
 sky130_fd_sc_hd__a21oi_1 _31899_ (.A1(_11211_),
    .A2(_11212_),
    .B1(net2964),
    .Y(_03880_));
 sky130_fd_sc_hd__nand3_1 _31900_ (.A(net1810),
    .B(net2906),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[18] ),
    .Y(_11213_));
 sky130_fd_sc_hd__nand2_1 _31901_ (.A(net2021),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[2] ),
    .Y(_11214_));
 sky130_fd_sc_hd__a21oi_1 _31903_ (.A1(_11213_),
    .A2(_11214_),
    .B1(net2965),
    .Y(_03881_));
 sky130_fd_sc_hd__nand3_1 _31905_ (.A(net1813),
    .B(net2906),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[19] ),
    .Y(_11217_));
 sky130_fd_sc_hd__nand2_1 _31906_ (.A(net2021),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[3] ),
    .Y(_11218_));
 sky130_fd_sc_hd__a21oi_1 _31907_ (.A1(_11217_),
    .A2(_11218_),
    .B1(net2965),
    .Y(_03882_));
 sky130_fd_sc_hd__nand3_1 _31908_ (.A(net1810),
    .B(net2906),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[20] ),
    .Y(_11219_));
 sky130_fd_sc_hd__nand2_1 _31909_ (.A(net2021),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[4] ),
    .Y(_11220_));
 sky130_fd_sc_hd__a21oi_1 _31910_ (.A1(_11219_),
    .A2(_11220_),
    .B1(net2960),
    .Y(_03883_));
 sky130_fd_sc_hd__nand3_1 _31911_ (.A(net1813),
    .B(net2907),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[21] ),
    .Y(_11221_));
 sky130_fd_sc_hd__nand2_1 _31912_ (.A(net2021),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[5] ),
    .Y(_11222_));
 sky130_fd_sc_hd__a21oi_1 _31913_ (.A1(_11221_),
    .A2(_11222_),
    .B1(net2963),
    .Y(_03884_));
 sky130_fd_sc_hd__nand3_1 _31914_ (.A(net1812),
    .B(net2907),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[22] ),
    .Y(_11223_));
 sky130_fd_sc_hd__nand2_1 _31915_ (.A(net2022),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[6] ),
    .Y(_11224_));
 sky130_fd_sc_hd__a21oi_1 _31916_ (.A1(_11223_),
    .A2(_11224_),
    .B1(net2964),
    .Y(_03885_));
 sky130_fd_sc_hd__nand3_1 _31917_ (.A(net1812),
    .B(net2907),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[23] ),
    .Y(_11225_));
 sky130_fd_sc_hd__nand2_1 _31918_ (.A(net2022),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[7] ),
    .Y(_11226_));
 sky130_fd_sc_hd__a21oi_1 _31919_ (.A1(_11225_),
    .A2(_11226_),
    .B1(net2964),
    .Y(_03886_));
 sky130_fd_sc_hd__nand3_1 _31920_ (.A(net1813),
    .B(net2907),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[24] ),
    .Y(_11227_));
 sky130_fd_sc_hd__nand2_1 _31921_ (.A(net2022),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[8] ),
    .Y(_11228_));
 sky130_fd_sc_hd__a21oi_1 _31922_ (.A1(_11227_),
    .A2(_11228_),
    .B1(net2963),
    .Y(_03887_));
 sky130_fd_sc_hd__nand3_1 _31923_ (.A(net1809),
    .B(net2906),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[25] ),
    .Y(_11229_));
 sky130_fd_sc_hd__nand2_1 _31924_ (.A(net2021),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[9] ),
    .Y(_11230_));
 sky130_fd_sc_hd__a21oi_1 _31925_ (.A1(_11229_),
    .A2(_11230_),
    .B1(net2960),
    .Y(_03888_));
 sky130_fd_sc_hd__nand3_1 _31926_ (.A(net1807),
    .B(net2906),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[3] ),
    .Y(_11231_));
 sky130_fd_sc_hd__nand2_1 _31927_ (.A(net2021),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.msip.x_data ),
    .Y(_11232_));
 sky130_fd_sc_hd__a21oi_1 _31928_ (.A1(_11231_),
    .A2(_11232_),
    .B1(net2958),
    .Y(_03889_));
 sky130_fd_sc_hd__nand3_1 _31929_ (.A(net1807),
    .B(net2906),
    .C(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[7] ),
    .Y(_11233_));
 sky130_fd_sc_hd__nand2_1 _31930_ (.A(net2021),
    .B(\inst$top.soc.cpu.exception.csr_bank.mip.mtip.x_data ),
    .Y(_11234_));
 sky130_fd_sc_hd__a21oi_1 _31931_ (.A1(_11233_),
    .A2(_11234_),
    .B1(net2959),
    .Y(_03890_));
 sky130_fd_sc_hd__o21ai_0 _31932_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mip_m_select ),
    .A2(net2253),
    .B1(net2090),
    .Y(_11235_));
 sky130_fd_sc_hd__a21oi_1 _31933_ (.A1(_20509_),
    .A2(net2253),
    .B1(_11235_),
    .Y(_03891_));
 sky130_fd_sc_hd__nor2_1 _31934_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip_m_select ),
    .B(net1893),
    .Y(_11236_));
 sky130_fd_sc_hd__o21ai_0 _31935_ (.A1(net2906),
    .A2(net2253),
    .B1(net2090),
    .Y(_11237_));
 sky130_fd_sc_hd__nor2_1 _31936_ (.A(_11236_),
    .B(_11237_),
    .Y(_03892_));
 sky130_fd_sc_hd__nor2_1 _31937_ (.A(net2905),
    .B(net671),
    .Y(_11238_));
 sky130_fd_sc_hd__nand2_1 _31938_ (.A(_11185_),
    .B(_11022_),
    .Y(_11239_));
 sky130_fd_sc_hd__nand2_1 _31939_ (.A(net671),
    .B(_11239_),
    .Y(_11240_));
 sky130_fd_sc_hd__nand2_1 _31941_ (.A(_11240_),
    .B(net2033),
    .Y(_11242_));
 sky130_fd_sc_hd__nor2_4 _31942_ (.A(_11238_),
    .B(_11242_),
    .Y(_03893_));
 sky130_fd_sc_hd__nand2_1 _31943_ (.A(net1809),
    .B(\inst$top.soc.cpu.exception.csr_bank.misa_w_select ),
    .Y(_11243_));
 sky130_fd_sc_hd__o21ai_0 _31946_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[0] ),
    .A2(net1654),
    .B1(net2090),
    .Y(_11246_));
 sky130_fd_sc_hd__a21oi_1 _31947_ (.A1(_20385_),
    .A2(net1654),
    .B1(_11246_),
    .Y(_03894_));
 sky130_fd_sc_hd__o21ai_0 _31948_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[10] ),
    .A2(net1656),
    .B1(net2068),
    .Y(_11247_));
 sky130_fd_sc_hd__a21oi_1 _31949_ (.A1(_20713_),
    .A2(net1656),
    .B1(_11247_),
    .Y(_03895_));
 sky130_fd_sc_hd__o21ai_0 _31951_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[11] ),
    .A2(net1653),
    .B1(net2084),
    .Y(_11249_));
 sky130_fd_sc_hd__a21oi_1 _31952_ (.A1(_20740_),
    .A2(net1653),
    .B1(_11249_),
    .Y(_03896_));
 sky130_fd_sc_hd__inv_1 _31953_ (.A(net1656),
    .Y(_11250_));
 sky130_fd_sc_hd__nand2_1 _31954_ (.A(_11250_),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[12] ),
    .Y(_11251_));
 sky130_fd_sc_hd__nand2_1 _31955_ (.A(net1656),
    .B(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[12] ),
    .Y(_11252_));
 sky130_fd_sc_hd__nand3_1 _31956_ (.A(_11251_),
    .B(net2044),
    .C(_11252_),
    .Y(_03897_));
 sky130_fd_sc_hd__nand2_1 _31957_ (.A(_11250_),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[13] ),
    .Y(_11253_));
 sky130_fd_sc_hd__nand2_1 _31958_ (.A(net1657),
    .B(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[13] ),
    .Y(_11254_));
 sky130_fd_sc_hd__a21oi_1 _31960_ (.A1(_11253_),
    .A2(_11254_),
    .B1(net2968),
    .Y(_03898_));
 sky130_fd_sc_hd__nand2_1 _31961_ (.A(_11250_),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[14] ),
    .Y(_11256_));
 sky130_fd_sc_hd__nand2_1 _31962_ (.A(net1656),
    .B(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[14] ),
    .Y(_11257_));
 sky130_fd_sc_hd__a21oi_1 _31963_ (.A1(_11256_),
    .A2(_11257_),
    .B1(net2953),
    .Y(_03899_));
 sky130_fd_sc_hd__o21ai_0 _31964_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[15] ),
    .A2(net1656),
    .B1(net2068),
    .Y(_11258_));
 sky130_fd_sc_hd__a21oi_1 _31965_ (.A1(_20816_),
    .A2(net1656),
    .B1(_11258_),
    .Y(_03900_));
 sky130_fd_sc_hd__o21ai_0 _31966_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[16] ),
    .A2(net1655),
    .B1(net2085),
    .Y(_11259_));
 sky130_fd_sc_hd__a21oi_1 _31967_ (.A1(_05611_),
    .A2(net1654),
    .B1(_11259_),
    .Y(_03901_));
 sky130_fd_sc_hd__o21ai_0 _31968_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[17] ),
    .A2(net1658),
    .B1(net2099),
    .Y(_11260_));
 sky130_fd_sc_hd__a21oi_1 _31969_ (.A1(_05629_),
    .A2(net1658),
    .B1(_11260_),
    .Y(_03902_));
 sky130_fd_sc_hd__o21ai_0 _31970_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[18] ),
    .A2(net1658),
    .B1(net2098),
    .Y(_11261_));
 sky130_fd_sc_hd__a21oi_1 _31971_ (.A1(_05651_),
    .A2(net1658),
    .B1(_11261_),
    .Y(_03903_));
 sky130_fd_sc_hd__o21ai_0 _31973_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[19] ),
    .A2(net1658),
    .B1(net2098),
    .Y(_11263_));
 sky130_fd_sc_hd__a21oi_1 _31974_ (.A1(_05679_),
    .A2(net1658),
    .B1(_11263_),
    .Y(_03904_));
 sky130_fd_sc_hd__o21ai_0 _31976_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[1] ),
    .A2(net1654),
    .B1(net2087),
    .Y(_11265_));
 sky130_fd_sc_hd__a21oi_1 _31977_ (.A1(_20436_),
    .A2(net1655),
    .B1(_11265_),
    .Y(_03905_));
 sky130_fd_sc_hd__o21ai_0 _31978_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[20] ),
    .A2(net1654),
    .B1(net2091),
    .Y(_11266_));
 sky130_fd_sc_hd__a21oi_1 _31979_ (.A1(_05698_),
    .A2(net1655),
    .B1(_11266_),
    .Y(_03906_));
 sky130_fd_sc_hd__o21ai_0 _31980_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[21] ),
    .A2(net1657),
    .B1(net2093),
    .Y(_11267_));
 sky130_fd_sc_hd__a21oi_1 _31981_ (.A1(_05719_),
    .A2(net1658),
    .B1(_11267_),
    .Y(_03907_));
 sky130_fd_sc_hd__o21ai_0 _31982_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[22] ),
    .A2(net1658),
    .B1(net2099),
    .Y(_11268_));
 sky130_fd_sc_hd__a21oi_1 _31983_ (.A1(_05737_),
    .A2(net1659),
    .B1(_11268_),
    .Y(_03908_));
 sky130_fd_sc_hd__o21ai_0 _31985_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[23] ),
    .A2(net1659),
    .B1(net2099),
    .Y(_11270_));
 sky130_fd_sc_hd__a21oi_1 _31986_ (.A1(_05758_),
    .A2(net1658),
    .B1(_11270_),
    .Y(_03909_));
 sky130_fd_sc_hd__o21ai_0 _31987_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[24] ),
    .A2(net1659),
    .B1(net2095),
    .Y(_11271_));
 sky130_fd_sc_hd__a21oi_1 _31988_ (.A1(_05775_),
    .A2(net1658),
    .B1(_11271_),
    .Y(_03910_));
 sky130_fd_sc_hd__o21ai_0 _31989_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[25] ),
    .A2(net1655),
    .B1(net2092),
    .Y(_11272_));
 sky130_fd_sc_hd__a21oi_1 _31990_ (.A1(_05795_),
    .A2(net1655),
    .B1(_11272_),
    .Y(_03911_));
 sky130_fd_sc_hd__o21ai_0 _31991_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[2] ),
    .A2(net1654),
    .B1(net2034),
    .Y(_11273_));
 sky130_fd_sc_hd__a21oi_1 _31992_ (.A1(_20471_),
    .A2(net1654),
    .B1(_11273_),
    .Y(_03912_));
 sky130_fd_sc_hd__o21ai_0 _31993_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[3] ),
    .A2(net1653),
    .B1(net2084),
    .Y(_11274_));
 sky130_fd_sc_hd__a21oi_1 _31994_ (.A1(_20517_),
    .A2(net1653),
    .B1(_11274_),
    .Y(_03913_));
 sky130_fd_sc_hd__o21ai_0 _31995_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[4] ),
    .A2(net1653),
    .B1(net2032),
    .Y(_11275_));
 sky130_fd_sc_hd__a21oi_1 _31996_ (.A1(_20547_),
    .A2(net1653),
    .B1(_11275_),
    .Y(_03914_));
 sky130_fd_sc_hd__o21ai_0 _31998_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[5] ),
    .A2(net1657),
    .B1(net2042),
    .Y(_11277_));
 sky130_fd_sc_hd__a21oi_1 _31999_ (.A1(_20574_),
    .A2(net1657),
    .B1(_11277_),
    .Y(_03915_));
 sky130_fd_sc_hd__o21ai_0 _32000_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[6] ),
    .A2(net1654),
    .B1(net2042),
    .Y(_11278_));
 sky130_fd_sc_hd__a21oi_1 _32001_ (.A1(_20602_),
    .A2(net1654),
    .B1(_11278_),
    .Y(_03916_));
 sky130_fd_sc_hd__o21ai_0 _32002_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[7] ),
    .A2(net1653),
    .B1(net2083),
    .Y(_11279_));
 sky130_fd_sc_hd__a21oi_1 _32003_ (.A1(_20634_),
    .A2(net1653),
    .B1(_11279_),
    .Y(_03917_));
 sky130_fd_sc_hd__nand2_1 _32004_ (.A(_11250_),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[8] ),
    .Y(_11280_));
 sky130_fd_sc_hd__nand2_1 _32007_ (.A(net1656),
    .B(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[8] ),
    .Y(_11283_));
 sky130_fd_sc_hd__nand3_1 _32008_ (.A(_11280_),
    .B(net2045),
    .C(_11283_),
    .Y(_03918_));
 sky130_fd_sc_hd__o21ai_0 _32009_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[9] ),
    .A2(net1656),
    .B1(net2045),
    .Y(_11284_));
 sky130_fd_sc_hd__a21oi_1 _32010_ (.A1(_20692_),
    .A2(net1656),
    .B1(_11284_),
    .Y(_03919_));
 sky130_fd_sc_hd__nand2_1 _32011_ (.A(_11250_),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[30] ),
    .Y(_11285_));
 sky130_fd_sc_hd__nand2_1 _32012_ (.A(net1657),
    .B(\inst$top.soc.cpu.exception.csr_bank.misa.mxl.x_data[0] ),
    .Y(_11286_));
 sky130_fd_sc_hd__nand3_1 _32013_ (.A(_11285_),
    .B(net2097),
    .C(_11286_),
    .Y(_03920_));
 sky130_fd_sc_hd__o21ai_0 _32014_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[31] ),
    .A2(net1653),
    .B1(net2032),
    .Y(_11287_));
 sky130_fd_sc_hd__a21oi_1 _32015_ (.A1(_05879_),
    .A2(net1653),
    .B1(_11287_),
    .Y(_03921_));
 sky130_fd_sc_hd__o21ai_0 _32016_ (.A1(\inst$top.soc.cpu.exception.csr_bank.misa_m_select ),
    .A2(net2252),
    .B1(net2092),
    .Y(_11288_));
 sky130_fd_sc_hd__a21oi_1 _32017_ (.A1(net2211),
    .A2(net2252),
    .B1(_11288_),
    .Y(_03922_));
 sky130_fd_sc_hd__nor2_1 _32018_ (.A(\inst$top.soc.cpu.exception.csr_bank.misa_m_select ),
    .B(net1893),
    .Y(_11289_));
 sky130_fd_sc_hd__o21ai_0 _32019_ (.A1(\inst$top.soc.cpu.exception.csr_bank.misa_w_select ),
    .A2(net2252),
    .B1(net2092),
    .Y(_11290_));
 sky130_fd_sc_hd__nor2_1 _32020_ (.A(_11289_),
    .B(_11290_),
    .Y(_03923_));
 sky130_fd_sc_hd__inv_1 _32021_ (.A(_11186_),
    .Y(_11291_));
 sky130_fd_sc_hd__nor2_1 _32022_ (.A(_11142_),
    .B(_11291_),
    .Y(_11292_));
 sky130_fd_sc_hd__nand2_1 _32023_ (.A(net633),
    .B(net2211),
    .Y(_11293_));
 sky130_fd_sc_hd__o21ai_1 _32024_ (.A1(_11292_),
    .A2(net633),
    .B1(_11293_),
    .Y(_11294_));
 sky130_fd_sc_hd__nor2_4 _32025_ (.A(net2936),
    .B(_11294_),
    .Y(_03924_));
 sky130_fd_sc_hd__nand2_1 _32026_ (.A(net1809),
    .B(net2901),
    .Y(_11295_));
 sky130_fd_sc_hd__o21ai_0 _32028_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[0] ),
    .A2(net1649),
    .B1(net2090),
    .Y(_11297_));
 sky130_fd_sc_hd__a21oi_1 _32029_ (.A1(_20391_),
    .A2(net1650),
    .B1(_11297_),
    .Y(_03925_));
 sky130_fd_sc_hd__nand2_1 _32030_ (.A(net1651),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[10] ),
    .Y(_11298_));
 sky130_fd_sc_hd__nand3_1 _32032_ (.A(net1811),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[10] ),
    .C(net2902),
    .Y(_11300_));
 sky130_fd_sc_hd__a21oi_1 _32033_ (.A1(_11298_),
    .A2(_11300_),
    .B1(net2953),
    .Y(_03926_));
 sky130_fd_sc_hd__nand2_1 _32034_ (.A(net1649),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[11] ),
    .Y(_11301_));
 sky130_fd_sc_hd__nand3_1 _32035_ (.A(net1808),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[11] ),
    .C(net2901),
    .Y(_11302_));
 sky130_fd_sc_hd__a21oi_1 _32036_ (.A1(_11301_),
    .A2(_11302_),
    .B1(net2958),
    .Y(_03927_));
 sky130_fd_sc_hd__nand2_1 _32037_ (.A(net1651),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[12] ),
    .Y(_11303_));
 sky130_fd_sc_hd__nand3_1 _32038_ (.A(net1811),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[12] ),
    .C(net2903),
    .Y(_11304_));
 sky130_fd_sc_hd__a21oi_1 _32039_ (.A1(_11303_),
    .A2(_11304_),
    .B1(net2961),
    .Y(_03928_));
 sky130_fd_sc_hd__nand2_1 _32040_ (.A(net1651),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[13] ),
    .Y(_11305_));
 sky130_fd_sc_hd__nand3_1 _32041_ (.A(net1811),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[13] ),
    .C(net2902),
    .Y(_11306_));
 sky130_fd_sc_hd__a21oi_1 _32042_ (.A1(_11305_),
    .A2(_11306_),
    .B1(net2968),
    .Y(_03929_));
 sky130_fd_sc_hd__nand2_1 _32043_ (.A(net1651),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[14] ),
    .Y(_11307_));
 sky130_fd_sc_hd__nand3_1 _32044_ (.A(net1811),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[14] ),
    .C(net2902),
    .Y(_11308_));
 sky130_fd_sc_hd__a21oi_1 _32045_ (.A1(_11307_),
    .A2(_11308_),
    .B1(net2953),
    .Y(_03930_));
 sky130_fd_sc_hd__nand2_1 _32046_ (.A(net1651),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[15] ),
    .Y(_11309_));
 sky130_fd_sc_hd__nand3_1 _32047_ (.A(net1811),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[15] ),
    .C(net2902),
    .Y(_11310_));
 sky130_fd_sc_hd__a21oi_1 _32048_ (.A1(_11309_),
    .A2(_11310_),
    .B1(net2952),
    .Y(_03931_));
 sky130_fd_sc_hd__nand2_1 _32049_ (.A(net1650),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[16] ),
    .Y(_11311_));
 sky130_fd_sc_hd__nand3_1 _32051_ (.A(net1809),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[16] ),
    .C(net2901),
    .Y(_11313_));
 sky130_fd_sc_hd__a21oi_1 _32052_ (.A1(_11311_),
    .A2(_11313_),
    .B1(net2960),
    .Y(_03932_));
 sky130_fd_sc_hd__nand2_1 _32053_ (.A(net1652),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[17] ),
    .Y(_11314_));
 sky130_fd_sc_hd__nand3_1 _32054_ (.A(net1813),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[17] ),
    .C(net2903),
    .Y(_11315_));
 sky130_fd_sc_hd__a21oi_1 _32055_ (.A1(_11314_),
    .A2(_11315_),
    .B1(net2964),
    .Y(_03933_));
 sky130_fd_sc_hd__nand2_1 _32057_ (.A(net1652),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[18] ),
    .Y(_11317_));
 sky130_fd_sc_hd__nand3_1 _32058_ (.A(net1813),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[18] ),
    .C(net2903),
    .Y(_11318_));
 sky130_fd_sc_hd__a21oi_1 _32060_ (.A1(_11317_),
    .A2(_11318_),
    .B1(net2965),
    .Y(_03934_));
 sky130_fd_sc_hd__nand2_1 _32061_ (.A(net1652),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[19] ),
    .Y(_11320_));
 sky130_fd_sc_hd__nand3_1 _32062_ (.A(net1813),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[19] ),
    .C(net2903),
    .Y(_11321_));
 sky130_fd_sc_hd__a21oi_1 _32063_ (.A1(_11320_),
    .A2(_11321_),
    .B1(net2965),
    .Y(_03935_));
 sky130_fd_sc_hd__o21ai_0 _32064_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[1] ),
    .A2(net1649),
    .B1(net2087),
    .Y(_11322_));
 sky130_fd_sc_hd__a21oi_1 _32065_ (.A1(_20433_),
    .A2(net1650),
    .B1(_11322_),
    .Y(_03936_));
 sky130_fd_sc_hd__nand2_1 _32066_ (.A(net1650),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[20] ),
    .Y(_11323_));
 sky130_fd_sc_hd__nand3_1 _32068_ (.A(net1810),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[20] ),
    .C(net2901),
    .Y(_11325_));
 sky130_fd_sc_hd__a21oi_1 _32069_ (.A1(_11323_),
    .A2(_11325_),
    .B1(net2960),
    .Y(_03937_));
 sky130_fd_sc_hd__nand2_1 _32070_ (.A(net1649),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[21] ),
    .Y(_11326_));
 sky130_fd_sc_hd__nand3_1 _32071_ (.A(net1811),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[21] ),
    .C(net2903),
    .Y(_11327_));
 sky130_fd_sc_hd__a21oi_1 _32072_ (.A1(_11326_),
    .A2(_11327_),
    .B1(net2961),
    .Y(_03938_));
 sky130_fd_sc_hd__nand2_1 _32073_ (.A(net1652),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[22] ),
    .Y(_11328_));
 sky130_fd_sc_hd__nand3_1 _32074_ (.A(net1812),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[22] ),
    .C(net2903),
    .Y(_11329_));
 sky130_fd_sc_hd__a21oi_1 _32075_ (.A1(_11328_),
    .A2(_11329_),
    .B1(net2964),
    .Y(_03939_));
 sky130_fd_sc_hd__nand2_1 _32076_ (.A(net1652),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[23] ),
    .Y(_11330_));
 sky130_fd_sc_hd__nand3_1 _32077_ (.A(net1812),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[23] ),
    .C(net2903),
    .Y(_11331_));
 sky130_fd_sc_hd__a21oi_1 _32078_ (.A1(_11330_),
    .A2(_11331_),
    .B1(net2971),
    .Y(_03940_));
 sky130_fd_sc_hd__nand2_1 _32079_ (.A(net1652),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[24] ),
    .Y(_11332_));
 sky130_fd_sc_hd__nand3_1 _32080_ (.A(net1812),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[24] ),
    .C(net2904),
    .Y(_11333_));
 sky130_fd_sc_hd__a21oi_1 _32081_ (.A1(_11332_),
    .A2(_11333_),
    .B1(net2969),
    .Y(_03941_));
 sky130_fd_sc_hd__nand2_1 _32082_ (.A(net1650),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[25] ),
    .Y(_11334_));
 sky130_fd_sc_hd__nand3_1 _32083_ (.A(net1809),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[25] ),
    .C(net2901),
    .Y(_11335_));
 sky130_fd_sc_hd__a21oi_1 _32084_ (.A1(_11334_),
    .A2(_11335_),
    .B1(net2960),
    .Y(_03942_));
 sky130_fd_sc_hd__nand2_1 _32085_ (.A(net1652),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[26] ),
    .Y(_11336_));
 sky130_fd_sc_hd__nand3_1 _32087_ (.A(net1813),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[26] ),
    .C(net2902),
    .Y(_11338_));
 sky130_fd_sc_hd__a21oi_1 _32088_ (.A1(_11336_),
    .A2(_11338_),
    .B1(net2971),
    .Y(_03943_));
 sky130_fd_sc_hd__nand2_1 _32089_ (.A(net1652),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[27] ),
    .Y(_11339_));
 sky130_fd_sc_hd__nand3_1 _32090_ (.A(net1812),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[27] ),
    .C(net2902),
    .Y(_11340_));
 sky130_fd_sc_hd__a21oi_1 _32091_ (.A1(_11339_),
    .A2(_11340_),
    .B1(net2969),
    .Y(_03944_));
 sky130_fd_sc_hd__nand2_1 _32093_ (.A(net1652),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[28] ),
    .Y(_11342_));
 sky130_fd_sc_hd__nand3_1 _32094_ (.A(net1812),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[28] ),
    .C(net2902),
    .Y(_11343_));
 sky130_fd_sc_hd__a21oi_1 _32096_ (.A1(_11342_),
    .A2(_11343_),
    .B1(net2969),
    .Y(_03945_));
 sky130_fd_sc_hd__nand2_1 _32097_ (.A(net1651),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[29] ),
    .Y(_11345_));
 sky130_fd_sc_hd__nand3_1 _32098_ (.A(net1814),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[29] ),
    .C(net2902),
    .Y(_11346_));
 sky130_fd_sc_hd__a21oi_1 _32099_ (.A1(_11345_),
    .A2(_11346_),
    .B1(net2968),
    .Y(_03946_));
 sky130_fd_sc_hd__nand2_1 _32100_ (.A(net1649),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[2] ),
    .Y(_11347_));
 sky130_fd_sc_hd__nand3_1 _32102_ (.A(net1808),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[2] ),
    .C(net2904),
    .Y(_11349_));
 sky130_fd_sc_hd__a21oi_1 _32103_ (.A1(_11347_),
    .A2(_11349_),
    .B1(net2936),
    .Y(_03947_));
 sky130_fd_sc_hd__nand2_1 _32104_ (.A(net1651),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[30] ),
    .Y(_11350_));
 sky130_fd_sc_hd__nand3_1 _32105_ (.A(net1814),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[30] ),
    .C(net2902),
    .Y(_11351_));
 sky130_fd_sc_hd__a21oi_1 _32106_ (.A1(_11350_),
    .A2(_11351_),
    .B1(net2962),
    .Y(_03948_));
 sky130_fd_sc_hd__nand2_1 _32107_ (.A(net1649),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[31] ),
    .Y(_11352_));
 sky130_fd_sc_hd__nand3_1 _32108_ (.A(net1807),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[31] ),
    .C(net2901),
    .Y(_11353_));
 sky130_fd_sc_hd__a21oi_1 _32109_ (.A1(_11352_),
    .A2(_11353_),
    .B1(net2937),
    .Y(_03949_));
 sky130_fd_sc_hd__nand2_1 _32110_ (.A(net1649),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[3] ),
    .Y(_11354_));
 sky130_fd_sc_hd__nand3_1 _32111_ (.A(net1808),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[3] ),
    .C(net2901),
    .Y(_11355_));
 sky130_fd_sc_hd__a21oi_1 _32112_ (.A1(_11354_),
    .A2(_11355_),
    .B1(net2958),
    .Y(_03950_));
 sky130_fd_sc_hd__nand2_1 _32113_ (.A(net1649),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[4] ),
    .Y(_11356_));
 sky130_fd_sc_hd__nand3_1 _32114_ (.A(net1807),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[4] ),
    .C(net2901),
    .Y(_11357_));
 sky130_fd_sc_hd__a21oi_1 _32115_ (.A1(_11356_),
    .A2(_11357_),
    .B1(net2936),
    .Y(_03951_));
 sky130_fd_sc_hd__nand2_1 _32116_ (.A(net1651),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[5] ),
    .Y(_11358_));
 sky130_fd_sc_hd__nand3_1 _32117_ (.A(net1811),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[5] ),
    .C(net2903),
    .Y(_11359_));
 sky130_fd_sc_hd__a21oi_1 _32118_ (.A1(_11358_),
    .A2(_11359_),
    .B1(net2940),
    .Y(_03952_));
 sky130_fd_sc_hd__nand2_1 _32119_ (.A(net1649),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[6] ),
    .Y(_11360_));
 sky130_fd_sc_hd__nand3_1 _32120_ (.A(net1808),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[6] ),
    .C(net2904),
    .Y(_11361_));
 sky130_fd_sc_hd__a21oi_1 _32121_ (.A1(_11360_),
    .A2(_11361_),
    .B1(net2940),
    .Y(_03953_));
 sky130_fd_sc_hd__nand2_1 _32122_ (.A(net1649),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[7] ),
    .Y(_11362_));
 sky130_fd_sc_hd__nand3_1 _32123_ (.A(net1807),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[7] ),
    .C(net2901),
    .Y(_11363_));
 sky130_fd_sc_hd__a21oi_1 _32124_ (.A1(_11362_),
    .A2(_11363_),
    .B1(net2937),
    .Y(_03954_));
 sky130_fd_sc_hd__nand2_1 _32125_ (.A(net1651),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[8] ),
    .Y(_11364_));
 sky130_fd_sc_hd__nand3_1 _32126_ (.A(net1811),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[8] ),
    .C(net2902),
    .Y(_11365_));
 sky130_fd_sc_hd__a21oi_1 _32128_ (.A1(_11364_),
    .A2(_11365_),
    .B1(net2942),
    .Y(_03955_));
 sky130_fd_sc_hd__nand2_1 _32129_ (.A(net1651),
    .B(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[9] ),
    .Y(_11367_));
 sky130_fd_sc_hd__nand3_1 _32130_ (.A(net1811),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[9] ),
    .C(net2903),
    .Y(_11368_));
 sky130_fd_sc_hd__a21oi_1 _32131_ (.A1(_11367_),
    .A2(_11368_),
    .B1(net2942),
    .Y(_03956_));
 sky130_fd_sc_hd__o21ai_0 _32132_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mscratch_m_select ),
    .A2(net2251),
    .B1(net2085),
    .Y(_11369_));
 sky130_fd_sc_hd__a21oi_1 _32133_ (.A1(_20390_),
    .A2(net2251),
    .B1(_11369_),
    .Y(_03957_));
 sky130_fd_sc_hd__inv_1 _32134_ (.A(\inst$top.soc.cpu.exception.csr_bank.mscratch_m_select ),
    .Y(_11370_));
 sky130_fd_sc_hd__o21ai_0 _32135_ (.A1(net2901),
    .A2(net2251),
    .B1(net2085),
    .Y(_11371_));
 sky130_fd_sc_hd__a21oi_1 _32136_ (.A1(_11370_),
    .A2(net2251),
    .B1(_11371_),
    .Y(_03958_));
 sky130_fd_sc_hd__nor2_1 _32137_ (.A(net2897),
    .B(net671),
    .Y(_11372_));
 sky130_fd_sc_hd__nor2_1 _32138_ (.A(_11017_),
    .B(_11014_),
    .Y(_11373_));
 sky130_fd_sc_hd__nand2_1 _32139_ (.A(_11018_),
    .B(_11373_),
    .Y(_11374_));
 sky130_fd_sc_hd__nor2_1 _32140_ (.A(_11374_),
    .B(_11023_),
    .Y(_11375_));
 sky130_fd_sc_hd__o21ai_1 _32141_ (.A1(_11375_),
    .A2(net633),
    .B1(net2033),
    .Y(_11376_));
 sky130_fd_sc_hd__nor2_4 _32142_ (.A(_11372_),
    .B(_11376_),
    .Y(_03959_));
 sky130_fd_sc_hd__nand2_1 _32143_ (.A(net1807),
    .B(\inst$top.soc.cpu.exception.csr_bank.mstatus_w_select ),
    .Y(_11377_));
 sky130_fd_sc_hd__nand3_1 _32144_ (.A(\inst$top.soc.cpu.m.source__valid ),
    .B(\inst$top.soc.cpu.exception.w_mret ),
    .C(\inst$top.soc.cpu.exception.w_mstatus.mpie ),
    .Y(_11378_));
 sky130_fd_sc_hd__nand2_1 _32145_ (.A(\inst$top.soc.cpu.m.source__valid ),
    .B(\inst$top.soc.cpu.exception.w_mret ),
    .Y(_11379_));
 sky130_fd_sc_hd__nand3_1 _32146_ (.A(_10913_),
    .B(_11379_),
    .C(\inst$top.soc.cpu.exception.csr_bank.mstatus.mie.x_data ),
    .Y(_11380_));
 sky130_fd_sc_hd__o21ai_0 _32147_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[3] ),
    .A2(_11377_),
    .B1(net2084),
    .Y(_11381_));
 sky130_fd_sc_hd__a31oi_1 _32148_ (.A1(_11377_),
    .A2(_11378_),
    .A3(_11380_),
    .B1(_11381_),
    .Y(_03960_));
 sky130_fd_sc_hd__nand2_1 _32149_ (.A(_10913_),
    .B(_20636_),
    .Y(_11382_));
 sky130_fd_sc_hd__o21ai_0 _32150_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mstatus.mpie.w_data ),
    .A2(_10913_),
    .B1(_11382_),
    .Y(_11383_));
 sky130_fd_sc_hd__o21ai_0 _32152_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[7] ),
    .A2(_11377_),
    .B1(net2083),
    .Y(_11385_));
 sky130_fd_sc_hd__a21oi_1 _32153_ (.A1(_11377_),
    .A2(_11383_),
    .B1(_11385_),
    .Y(_03961_));
 sky130_fd_sc_hd__inv_1 _32154_ (.A(_11377_),
    .Y(_11386_));
 sky130_fd_sc_hd__nand2_1 _32155_ (.A(_11386_),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[11] ),
    .Y(_11387_));
 sky130_fd_sc_hd__nand2_1 _32156_ (.A(_11377_),
    .B(\inst$top.soc.cpu.exception.csr_bank.mstatus.mpp.x_data[0] ),
    .Y(_11388_));
 sky130_fd_sc_hd__nand3_1 _32157_ (.A(_11387_),
    .B(net2088),
    .C(_11388_),
    .Y(_03962_));
 sky130_fd_sc_hd__nand2_1 _32158_ (.A(_11386_),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[12] ),
    .Y(_11389_));
 sky130_fd_sc_hd__nand2_1 _32159_ (.A(_11377_),
    .B(\inst$top.soc.cpu.exception.csr_bank.mstatus.mpp.x_data[1] ),
    .Y(_11390_));
 sky130_fd_sc_hd__nand3_1 _32160_ (.A(_11389_),
    .B(net2088),
    .C(_11390_),
    .Y(_03963_));
 sky130_fd_sc_hd__o21ai_0 _32161_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mstatus_m_select ),
    .A2(net2221),
    .B1(net2083),
    .Y(_11391_));
 sky130_fd_sc_hd__a21oi_1 _32162_ (.A1(_20635_),
    .A2(net2221),
    .B1(_11391_),
    .Y(_03964_));
 sky130_fd_sc_hd__nor2_1 _32163_ (.A(\inst$top.soc.cpu.exception.csr_bank.mstatus_m_select ),
    .B(net1884),
    .Y(_11392_));
 sky130_fd_sc_hd__o21ai_0 _32164_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mstatus_w_select ),
    .A2(net2221),
    .B1(net2083),
    .Y(_11393_));
 sky130_fd_sc_hd__nor2_1 _32165_ (.A(_11392_),
    .B(_11393_),
    .Y(_03965_));
 sky130_fd_sc_hd__nor2_1 _32166_ (.A(_11374_),
    .B(_11291_),
    .Y(_11394_));
 sky130_fd_sc_hd__nand2_1 _32167_ (.A(net633),
    .B(_20635_),
    .Y(_11395_));
 sky130_fd_sc_hd__o21ai_1 _32168_ (.A1(_11394_),
    .A2(net633),
    .B1(_11395_),
    .Y(_11396_));
 sky130_fd_sc_hd__nor2_4 _32169_ (.A(net2958),
    .B(_11396_),
    .Y(_03966_));
 sky130_fd_sc_hd__nand2_1 _32170_ (.A(net1807),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval_w_select ),
    .Y(_11397_));
 sky130_fd_sc_hd__nand2_1 _32171_ (.A(_11397_),
    .B(_10913_),
    .Y(_11398_));
 sky130_fd_sc_hd__inv_1 _32172_ (.A(_11398_),
    .Y(_11399_));
 sky130_fd_sc_hd__nand2_1 _32174_ (.A(net1088),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[0] ),
    .Y(_11401_));
 sky130_fd_sc_hd__inv_1 _32175_ (.A(_11397_),
    .Y(_11402_));
 sky130_fd_sc_hd__nand2_1 _32177_ (.A(net1233),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[0] ),
    .Y(_11404_));
 sky130_fd_sc_hd__nand2_1 _32178_ (.A(net1873),
    .B(\inst$top.soc.cpu.exception.w_data$51[0] ),
    .Y(_11405_));
 sky130_fd_sc_hd__a31oi_1 _32179_ (.A1(_11401_),
    .A2(_11404_),
    .A3(_11405_),
    .B1(net2959),
    .Y(_03967_));
 sky130_fd_sc_hd__nand2_1 _32180_ (.A(net1089),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[10] ),
    .Y(_11406_));
 sky130_fd_sc_hd__nand2_1 _32181_ (.A(net1234),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[10] ),
    .Y(_11407_));
 sky130_fd_sc_hd__nand2_1 _32182_ (.A(net1879),
    .B(\inst$top.soc.cpu.exception.w_data$51[10] ),
    .Y(_11408_));
 sky130_fd_sc_hd__a31oi_1 _32183_ (.A1(_11406_),
    .A2(_11407_),
    .A3(_11408_),
    .B1(net2968),
    .Y(_03968_));
 sky130_fd_sc_hd__nand2_1 _32184_ (.A(net1088),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[11] ),
    .Y(_11409_));
 sky130_fd_sc_hd__nand2_1 _32185_ (.A(net1233),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[11] ),
    .Y(_11410_));
 sky130_fd_sc_hd__nand2_1 _32186_ (.A(net1874),
    .B(\inst$top.soc.cpu.exception.w_data$51[11] ),
    .Y(_11411_));
 sky130_fd_sc_hd__a31oi_1 _32187_ (.A1(_11409_),
    .A2(_11410_),
    .A3(_11411_),
    .B1(net2961),
    .Y(_03969_));
 sky130_fd_sc_hd__nand2_1 _32188_ (.A(net1090),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[12] ),
    .Y(_11412_));
 sky130_fd_sc_hd__nand2_1 _32189_ (.A(net1235),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[12] ),
    .Y(_11413_));
 sky130_fd_sc_hd__nand2_1 _32190_ (.A(net1876),
    .B(\inst$top.soc.cpu.exception.w_data$51[12] ),
    .Y(_11414_));
 sky130_fd_sc_hd__a31oi_1 _32191_ (.A1(_11412_),
    .A2(_11413_),
    .A3(_11414_),
    .B1(net2962),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2_1 _32192_ (.A(net1089),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[13] ),
    .Y(_11415_));
 sky130_fd_sc_hd__nand2_1 _32193_ (.A(net1234),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[13] ),
    .Y(_11416_));
 sky130_fd_sc_hd__nand2_1 _32195_ (.A(net1879),
    .B(\inst$top.soc.cpu.exception.w_data$51[13] ),
    .Y(_11418_));
 sky130_fd_sc_hd__a31oi_1 _32196_ (.A1(_11415_),
    .A2(_11416_),
    .A3(_11418_),
    .B1(net2968),
    .Y(_03971_));
 sky130_fd_sc_hd__nand2_1 _32197_ (.A(net1089),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[14] ),
    .Y(_11419_));
 sky130_fd_sc_hd__nand2_1 _32198_ (.A(net1234),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[14] ),
    .Y(_11420_));
 sky130_fd_sc_hd__nand2_1 _32199_ (.A(net1879),
    .B(\inst$top.soc.cpu.exception.w_data$51[14] ),
    .Y(_11421_));
 sky130_fd_sc_hd__a31oi_1 _32200_ (.A1(_11419_),
    .A2(_11420_),
    .A3(_11421_),
    .B1(net2952),
    .Y(_03972_));
 sky130_fd_sc_hd__nand2_1 _32201_ (.A(net1089),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[15] ),
    .Y(_11422_));
 sky130_fd_sc_hd__nand2_1 _32202_ (.A(net1234),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[15] ),
    .Y(_11423_));
 sky130_fd_sc_hd__nand2_1 _32203_ (.A(net1879),
    .B(\inst$top.soc.cpu.exception.w_data$51[15] ),
    .Y(_11424_));
 sky130_fd_sc_hd__a31oi_1 _32205_ (.A1(_11422_),
    .A2(_11423_),
    .A3(_11424_),
    .B1(net2953),
    .Y(_03973_));
 sky130_fd_sc_hd__nand2_1 _32206_ (.A(net1090),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[16] ),
    .Y(_11426_));
 sky130_fd_sc_hd__nand2_1 _32207_ (.A(net1235),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[16] ),
    .Y(_11427_));
 sky130_fd_sc_hd__nand2_1 _32208_ (.A(net1880),
    .B(\inst$top.soc.cpu.exception.w_data$51[16] ),
    .Y(_11428_));
 sky130_fd_sc_hd__a31oi_1 _32209_ (.A1(_11426_),
    .A2(_11427_),
    .A3(_11428_),
    .B1(net2962),
    .Y(_03974_));
 sky130_fd_sc_hd__nand2_1 _32210_ (.A(net1090),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[17] ),
    .Y(_11429_));
 sky130_fd_sc_hd__nand2_1 _32211_ (.A(net1235),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[17] ),
    .Y(_11430_));
 sky130_fd_sc_hd__nand2_1 _32212_ (.A(net1880),
    .B(\inst$top.soc.cpu.exception.w_data$51[17] ),
    .Y(_11431_));
 sky130_fd_sc_hd__a31oi_1 _32213_ (.A1(_11429_),
    .A2(_11430_),
    .A3(_11431_),
    .B1(net2964),
    .Y(_03975_));
 sky130_fd_sc_hd__nand2_1 _32214_ (.A(net1090),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[18] ),
    .Y(_11432_));
 sky130_fd_sc_hd__nand2_1 _32215_ (.A(net1235),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[18] ),
    .Y(_11433_));
 sky130_fd_sc_hd__nand2_1 _32216_ (.A(net1876),
    .B(\inst$top.soc.cpu.exception.w_data$51[18] ),
    .Y(_11434_));
 sky130_fd_sc_hd__a31oi_1 _32217_ (.A1(_11432_),
    .A2(_11433_),
    .A3(_11434_),
    .B1(net2963),
    .Y(_03976_));
 sky130_fd_sc_hd__nand2_1 _32219_ (.A(net1090),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[19] ),
    .Y(_11436_));
 sky130_fd_sc_hd__nand2_1 _32221_ (.A(net1235),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[19] ),
    .Y(_11438_));
 sky130_fd_sc_hd__nand2_1 _32222_ (.A(net1876),
    .B(\inst$top.soc.cpu.exception.w_data$51[19] ),
    .Y(_11439_));
 sky130_fd_sc_hd__a31oi_1 _32223_ (.A1(_11436_),
    .A2(_11438_),
    .A3(_11439_),
    .B1(net2963),
    .Y(_03977_));
 sky130_fd_sc_hd__nand2_1 _32224_ (.A(net1088),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[1] ),
    .Y(_11440_));
 sky130_fd_sc_hd__nand2_1 _32225_ (.A(net1233),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[1] ),
    .Y(_11441_));
 sky130_fd_sc_hd__nand2_1 _32226_ (.A(net1875),
    .B(\inst$top.soc.cpu.exception.w_data$51[1] ),
    .Y(_11442_));
 sky130_fd_sc_hd__a31oi_1 _32227_ (.A1(_11440_),
    .A2(_11441_),
    .A3(_11442_),
    .B1(net2959),
    .Y(_03978_));
 sky130_fd_sc_hd__nand2_1 _32228_ (.A(net1088),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[20] ),
    .Y(_11443_));
 sky130_fd_sc_hd__nand2_1 _32229_ (.A(net1233),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[20] ),
    .Y(_11444_));
 sky130_fd_sc_hd__nand2_1 _32230_ (.A(net1875),
    .B(\inst$top.soc.cpu.exception.w_data$51[20] ),
    .Y(_11445_));
 sky130_fd_sc_hd__a31oi_1 _32231_ (.A1(_11443_),
    .A2(_11444_),
    .A3(_11445_),
    .B1(net2965),
    .Y(_03979_));
 sky130_fd_sc_hd__nand2_1 _32232_ (.A(net1090),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[21] ),
    .Y(_11446_));
 sky130_fd_sc_hd__nand2_1 _32233_ (.A(net1235),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[21] ),
    .Y(_11447_));
 sky130_fd_sc_hd__nand2_1 _32234_ (.A(net1874),
    .B(\inst$top.soc.cpu.exception.w_data$51[21] ),
    .Y(_11448_));
 sky130_fd_sc_hd__a31oi_1 _32235_ (.A1(_11446_),
    .A2(_11447_),
    .A3(_11448_),
    .B1(net2961),
    .Y(_03980_));
 sky130_fd_sc_hd__nand2_1 _32236_ (.A(net1091),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[22] ),
    .Y(_11449_));
 sky130_fd_sc_hd__nand2_1 _32237_ (.A(net1236),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[22] ),
    .Y(_11450_));
 sky130_fd_sc_hd__nand2_1 _32239_ (.A(net1878),
    .B(\inst$top.soc.cpu.exception.w_data$51[22] ),
    .Y(_11452_));
 sky130_fd_sc_hd__a31oi_1 _32240_ (.A1(_11449_),
    .A2(_11450_),
    .A3(_11452_),
    .B1(net2971),
    .Y(_03981_));
 sky130_fd_sc_hd__nand2_1 _32241_ (.A(net1089),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[23] ),
    .Y(_11453_));
 sky130_fd_sc_hd__nand2_1 _32242_ (.A(net1234),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[23] ),
    .Y(_11454_));
 sky130_fd_sc_hd__nand2_1 _32243_ (.A(net1878),
    .B(\inst$top.soc.cpu.exception.w_data$51[23] ),
    .Y(_11455_));
 sky130_fd_sc_hd__a31oi_1 _32244_ (.A1(_11453_),
    .A2(_11454_),
    .A3(_11455_),
    .B1(net2971),
    .Y(_03982_));
 sky130_fd_sc_hd__nand2_1 _32245_ (.A(net1089),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[24] ),
    .Y(_11456_));
 sky130_fd_sc_hd__nand2_1 _32246_ (.A(net1234),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[24] ),
    .Y(_11457_));
 sky130_fd_sc_hd__nand2_1 _32247_ (.A(net1877),
    .B(\inst$top.soc.cpu.exception.w_data$51[24] ),
    .Y(_11458_));
 sky130_fd_sc_hd__a31oi_1 _32249_ (.A1(_11456_),
    .A2(_11457_),
    .A3(_11458_),
    .B1(net2969),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_1 _32250_ (.A(net1088),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[25] ),
    .Y(_11460_));
 sky130_fd_sc_hd__nand2_1 _32251_ (.A(net1233),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[25] ),
    .Y(_11461_));
 sky130_fd_sc_hd__nand2_1 _32252_ (.A(net1873),
    .B(\inst$top.soc.cpu.exception.w_data$51[25] ),
    .Y(_11462_));
 sky130_fd_sc_hd__a31oi_1 _32253_ (.A1(_11460_),
    .A2(_11461_),
    .A3(_11462_),
    .B1(net2966),
    .Y(_03984_));
 sky130_fd_sc_hd__nand2_1 _32254_ (.A(net1089),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[26] ),
    .Y(_11463_));
 sky130_fd_sc_hd__nand2_1 _32255_ (.A(net1234),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[26] ),
    .Y(_11464_));
 sky130_fd_sc_hd__nand2_1 _32256_ (.A(net1878),
    .B(\inst$top.soc.cpu.exception.w_data$51[26] ),
    .Y(_11465_));
 sky130_fd_sc_hd__a31oi_1 _32257_ (.A1(_11463_),
    .A2(_11464_),
    .A3(_11465_),
    .B1(net2973),
    .Y(_03985_));
 sky130_fd_sc_hd__nand2_1 _32258_ (.A(net1089),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[27] ),
    .Y(_11466_));
 sky130_fd_sc_hd__nand2_1 _32259_ (.A(net1234),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[27] ),
    .Y(_11467_));
 sky130_fd_sc_hd__nand2_1 _32260_ (.A(net1877),
    .B(\inst$top.soc.cpu.exception.w_data$51[27] ),
    .Y(_11468_));
 sky130_fd_sc_hd__a31oi_1 _32261_ (.A1(_11466_),
    .A2(_11467_),
    .A3(_11468_),
    .B1(net2970),
    .Y(_03986_));
 sky130_fd_sc_hd__nand2_1 _32263_ (.A(net1090),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[28] ),
    .Y(_11470_));
 sky130_fd_sc_hd__nand2_1 _32265_ (.A(net1235),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[28] ),
    .Y(_11472_));
 sky130_fd_sc_hd__nand2_1 _32266_ (.A(net1877),
    .B(\inst$top.soc.cpu.exception.w_data$51[28] ),
    .Y(_11473_));
 sky130_fd_sc_hd__a31oi_1 _32267_ (.A1(_11470_),
    .A2(_11472_),
    .A3(_11473_),
    .B1(net2969),
    .Y(_03987_));
 sky130_fd_sc_hd__nand2_1 _32268_ (.A(net1091),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[29] ),
    .Y(_11474_));
 sky130_fd_sc_hd__nand2_1 _32269_ (.A(net1236),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[29] ),
    .Y(_11475_));
 sky130_fd_sc_hd__nand2_1 _32270_ (.A(net1878),
    .B(\inst$top.soc.cpu.exception.w_data$51[29] ),
    .Y(_11476_));
 sky130_fd_sc_hd__a31oi_1 _32271_ (.A1(_11474_),
    .A2(_11475_),
    .A3(_11476_),
    .B1(net2968),
    .Y(_03988_));
 sky130_fd_sc_hd__nand2_1 _32272_ (.A(net1091),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[2] ),
    .Y(_11477_));
 sky130_fd_sc_hd__nand2_1 _32273_ (.A(net1236),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[2] ),
    .Y(_11478_));
 sky130_fd_sc_hd__nand2_1 _32274_ (.A(net1874),
    .B(\inst$top.soc.cpu.exception.w_data$51[2] ),
    .Y(_11479_));
 sky130_fd_sc_hd__a31oi_1 _32275_ (.A1(_11477_),
    .A2(_11478_),
    .A3(_11479_),
    .B1(net2936),
    .Y(_03989_));
 sky130_fd_sc_hd__nand2_1 _32276_ (.A(net1089),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[30] ),
    .Y(_11480_));
 sky130_fd_sc_hd__nand2_1 _32277_ (.A(net1234),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[30] ),
    .Y(_11481_));
 sky130_fd_sc_hd__nand2_1 _32278_ (.A(net1879),
    .B(\inst$top.soc.cpu.exception.w_data$51[30] ),
    .Y(_11482_));
 sky130_fd_sc_hd__a31oi_1 _32279_ (.A1(_11480_),
    .A2(_11481_),
    .A3(_11482_),
    .B1(net2962),
    .Y(_03990_));
 sky130_fd_sc_hd__nand2_1 _32280_ (.A(net1088),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[31] ),
    .Y(_11483_));
 sky130_fd_sc_hd__nand2_1 _32281_ (.A(net1233),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[31] ),
    .Y(_11484_));
 sky130_fd_sc_hd__nand2_1 _32282_ (.A(net1872),
    .B(\inst$top.soc.cpu.exception.w_data$51[31] ),
    .Y(_11485_));
 sky130_fd_sc_hd__a31oi_1 _32283_ (.A1(_11483_),
    .A2(_11484_),
    .A3(_11485_),
    .B1(net2937),
    .Y(_03991_));
 sky130_fd_sc_hd__nand2_1 _32284_ (.A(net1088),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[3] ),
    .Y(_11486_));
 sky130_fd_sc_hd__nand2_1 _32285_ (.A(net1233),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[3] ),
    .Y(_11487_));
 sky130_fd_sc_hd__nand2_1 _32286_ (.A(net1872),
    .B(\inst$top.soc.cpu.exception.w_data$51[3] ),
    .Y(_11488_));
 sky130_fd_sc_hd__a31oi_1 _32287_ (.A1(_11486_),
    .A2(_11487_),
    .A3(_11488_),
    .B1(net2958),
    .Y(_03992_));
 sky130_fd_sc_hd__nand2_1 _32288_ (.A(net1088),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[4] ),
    .Y(_11489_));
 sky130_fd_sc_hd__nand2_1 _32289_ (.A(net1233),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[4] ),
    .Y(_11490_));
 sky130_fd_sc_hd__nand2_1 _32290_ (.A(net1872),
    .B(\inst$top.soc.cpu.exception.w_data$51[4] ),
    .Y(_11491_));
 sky130_fd_sc_hd__a31oi_1 _32292_ (.A1(_11489_),
    .A2(_11490_),
    .A3(_11491_),
    .B1(net2937),
    .Y(_03993_));
 sky130_fd_sc_hd__nand2_1 _32293_ (.A(net1090),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[5] ),
    .Y(_11493_));
 sky130_fd_sc_hd__nand2_1 _32294_ (.A(net1235),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[5] ),
    .Y(_11494_));
 sky130_fd_sc_hd__nand2_1 _32295_ (.A(net1874),
    .B(\inst$top.soc.cpu.exception.w_data$51[5] ),
    .Y(_11495_));
 sky130_fd_sc_hd__a31oi_1 _32296_ (.A1(_11493_),
    .A2(_11494_),
    .A3(_11495_),
    .B1(net2940),
    .Y(_03994_));
 sky130_fd_sc_hd__nand2_1 _32297_ (.A(net1088),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[6] ),
    .Y(_11496_));
 sky130_fd_sc_hd__nand2_1 _32298_ (.A(net1233),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[6] ),
    .Y(_11497_));
 sky130_fd_sc_hd__nand2_1 _32299_ (.A(net1874),
    .B(\inst$top.soc.cpu.exception.w_data$51[6] ),
    .Y(_11498_));
 sky130_fd_sc_hd__a31oi_1 _32300_ (.A1(_11496_),
    .A2(_11497_),
    .A3(_11498_),
    .B1(net2940),
    .Y(_03995_));
 sky130_fd_sc_hd__nand2_1 _32301_ (.A(net1088),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[7] ),
    .Y(_11499_));
 sky130_fd_sc_hd__nand2_1 _32302_ (.A(net1233),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[7] ),
    .Y(_11500_));
 sky130_fd_sc_hd__nand2_1 _32303_ (.A(net1872),
    .B(\inst$top.soc.cpu.exception.w_data$51[7] ),
    .Y(_11501_));
 sky130_fd_sc_hd__a31oi_1 _32304_ (.A1(_11499_),
    .A2(_11500_),
    .A3(_11501_),
    .B1(net2957),
    .Y(_03996_));
 sky130_fd_sc_hd__nand2_1 _32305_ (.A(net1089),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[8] ),
    .Y(_11502_));
 sky130_fd_sc_hd__nand2_1 _32306_ (.A(net1234),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[8] ),
    .Y(_11503_));
 sky130_fd_sc_hd__nand2_1 _32307_ (.A(net1876),
    .B(\inst$top.soc.cpu.exception.w_data$51[8] ),
    .Y(_11504_));
 sky130_fd_sc_hd__a31oi_1 _32308_ (.A1(_11502_),
    .A2(_11503_),
    .A3(_11504_),
    .B1(net2953),
    .Y(_03997_));
 sky130_fd_sc_hd__nand2_1 _32309_ (.A(net1090),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[9] ),
    .Y(_11505_));
 sky130_fd_sc_hd__nand2_1 _32310_ (.A(net1235),
    .B(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[9] ),
    .Y(_11506_));
 sky130_fd_sc_hd__nand2_1 _32311_ (.A(net1876),
    .B(\inst$top.soc.cpu.exception.w_data$51[9] ),
    .Y(_11507_));
 sky130_fd_sc_hd__a31oi_1 _32312_ (.A1(_11505_),
    .A2(_11506_),
    .A3(_11507_),
    .B1(net2942),
    .Y(_03998_));
 sky130_fd_sc_hd__nor2_1 _32313_ (.A(net2893),
    .B(net1883),
    .Y(_11508_));
 sky130_fd_sc_hd__o21ai_0 _32315_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mtval_m_select ),
    .A2(net2220),
    .B1(net2083),
    .Y(_11510_));
 sky130_fd_sc_hd__nor2_1 _32316_ (.A(_11508_),
    .B(_11510_),
    .Y(_03999_));
 sky130_fd_sc_hd__nor2_1 _32317_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtval_m_select ),
    .B(net1883),
    .Y(_11511_));
 sky130_fd_sc_hd__o21ai_0 _32318_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mtval_w_select ),
    .A2(net2220),
    .B1(net2083),
    .Y(_11512_));
 sky130_fd_sc_hd__nor2_1 _32319_ (.A(_11511_),
    .B(_11512_),
    .Y(_04000_));
 sky130_fd_sc_hd__nand2_1 _32320_ (.A(net633),
    .B(net2893),
    .Y(_11513_));
 sky130_fd_sc_hd__nor4_1 _32321_ (.A(_11015_),
    .B(net1031),
    .C(_11019_),
    .D(_11023_),
    .Y(_11514_));
 sky130_fd_sc_hd__nand3_1 _32322_ (.A(net663),
    .B(net753),
    .C(_11514_),
    .Y(_11515_));
 sky130_fd_sc_hd__a21oi_4 _32323_ (.A1(_11513_),
    .A2(_11515_),
    .B1(net2936),
    .Y(_04001_));
 sky130_fd_sc_hd__nand2_1 _32324_ (.A(net1809),
    .B(\inst$top.soc.cpu.exception.csr_bank.mtvec_w_select ),
    .Y(_11516_));
 sky130_fd_sc_hd__o21ai_0 _32327_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[2] ),
    .A2(net1641),
    .B1(net2034),
    .Y(_11519_));
 sky130_fd_sc_hd__a21oi_1 _32328_ (.A1(_20472_),
    .A2(net1641),
    .B1(_11519_),
    .Y(_04002_));
 sky130_fd_sc_hd__o21ai_0 _32329_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[12] ),
    .A2(net1644),
    .B1(net2043),
    .Y(_11520_));
 sky130_fd_sc_hd__a21oi_1 _32330_ (.A1(_20760_),
    .A2(net1644),
    .B1(_11520_),
    .Y(_04003_));
 sky130_fd_sc_hd__o21ai_0 _32331_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[13] ),
    .A2(net1643),
    .B1(net2104),
    .Y(_11521_));
 sky130_fd_sc_hd__a21oi_1 _32332_ (.A1(_20778_),
    .A2(net1643),
    .B1(_11521_),
    .Y(_04004_));
 sky130_fd_sc_hd__o21ai_0 _32333_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[14] ),
    .A2(net1643),
    .B1(net2069),
    .Y(_11522_));
 sky130_fd_sc_hd__a21oi_1 _32334_ (.A1(_20796_),
    .A2(net1643),
    .B1(_11522_),
    .Y(_04005_));
 sky130_fd_sc_hd__o21ai_0 _32335_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[15] ),
    .A2(net1643),
    .B1(net2068),
    .Y(_11523_));
 sky130_fd_sc_hd__a21oi_1 _32336_ (.A1(_20817_),
    .A2(net1643),
    .B1(_11523_),
    .Y(_04006_));
 sky130_fd_sc_hd__o21ai_0 _32337_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[16] ),
    .A2(net1645),
    .B1(net2097),
    .Y(_11524_));
 sky130_fd_sc_hd__a21oi_1 _32338_ (.A1(_05605_),
    .A2(net1645),
    .B1(_11524_),
    .Y(_04007_));
 sky130_fd_sc_hd__inv_1 _32339_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[15] ),
    .Y(_11525_));
 sky130_fd_sc_hd__o21ai_0 _32340_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[17] ),
    .A2(net1647),
    .B1(net2099),
    .Y(_11526_));
 sky130_fd_sc_hd__a21oi_1 _32341_ (.A1(_11525_),
    .A2(net1647),
    .B1(_11526_),
    .Y(_04008_));
 sky130_fd_sc_hd__inv_1 _32342_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[16] ),
    .Y(_11527_));
 sky130_fd_sc_hd__o21ai_0 _32343_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[18] ),
    .A2(net1647),
    .B1(net2098),
    .Y(_11528_));
 sky130_fd_sc_hd__a21oi_1 _32344_ (.A1(_11527_),
    .A2(net1647),
    .B1(_11528_),
    .Y(_04009_));
 sky130_fd_sc_hd__inv_1 _32345_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[17] ),
    .Y(_11529_));
 sky130_fd_sc_hd__o21ai_0 _32348_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[19] ),
    .A2(net1647),
    .B1(net2098),
    .Y(_11532_));
 sky130_fd_sc_hd__a21oi_1 _32349_ (.A1(_11529_),
    .A2(net1647),
    .B1(_11532_),
    .Y(_04010_));
 sky130_fd_sc_hd__o21ai_0 _32350_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[20] ),
    .A2(net1648),
    .B1(net2098),
    .Y(_11533_));
 sky130_fd_sc_hd__a21oi_1 _32351_ (.A1(_05695_),
    .A2(net1642),
    .B1(_11533_),
    .Y(_04011_));
 sky130_fd_sc_hd__inv_1 _32352_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[19] ),
    .Y(_11534_));
 sky130_fd_sc_hd__o21ai_0 _32354_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[21] ),
    .A2(net1644),
    .B1(net2093),
    .Y(_11536_));
 sky130_fd_sc_hd__a21oi_1 _32355_ (.A1(_11534_),
    .A2(net1644),
    .B1(_11536_),
    .Y(_04012_));
 sky130_fd_sc_hd__o21ai_0 _32356_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[3] ),
    .A2(net1641),
    .B1(net2088),
    .Y(_11537_));
 sky130_fd_sc_hd__a21oi_1 _32357_ (.A1(_20512_),
    .A2(net1642),
    .B1(_11537_),
    .Y(_04013_));
 sky130_fd_sc_hd__o21ai_0 _32358_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[22] ),
    .A2(net1645),
    .B1(net2110),
    .Y(_11538_));
 sky130_fd_sc_hd__a21oi_1 _32359_ (.A1(_05734_),
    .A2(net1646),
    .B1(_11538_),
    .Y(_04014_));
 sky130_fd_sc_hd__inv_1 _32360_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[21] ),
    .Y(_11539_));
 sky130_fd_sc_hd__o21ai_0 _32361_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[23] ),
    .A2(net1645),
    .B1(net2110),
    .Y(_11540_));
 sky130_fd_sc_hd__a21oi_1 _32362_ (.A1(_11539_),
    .A2(net1646),
    .B1(_11540_),
    .Y(_04015_));
 sky130_fd_sc_hd__inv_1 _32363_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[22] ),
    .Y(_11541_));
 sky130_fd_sc_hd__o21ai_0 _32364_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[24] ),
    .A2(net1645),
    .B1(net2105),
    .Y(_11542_));
 sky130_fd_sc_hd__a21oi_1 _32365_ (.A1(_11541_),
    .A2(net1645),
    .B1(_11542_),
    .Y(_04016_));
 sky130_fd_sc_hd__inv_1 _32366_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[23] ),
    .Y(_11543_));
 sky130_fd_sc_hd__o21ai_0 _32367_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[25] ),
    .A2(net1648),
    .B1(net2092),
    .Y(_11544_));
 sky130_fd_sc_hd__a21oi_1 _32368_ (.A1(_11543_),
    .A2(net1648),
    .B1(_11544_),
    .Y(_04017_));
 sky130_fd_sc_hd__o21ai_0 _32369_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[26] ),
    .A2(net1645),
    .B1(net2110),
    .Y(_11545_));
 sky130_fd_sc_hd__a21oi_1 _32370_ (.A1(_05814_),
    .A2(net1646),
    .B1(_11545_),
    .Y(_04018_));
 sky130_fd_sc_hd__o21ai_0 _32371_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[27] ),
    .A2(net1645),
    .B1(net2105),
    .Y(_11546_));
 sky130_fd_sc_hd__a21oi_1 _32372_ (.A1(_05827_),
    .A2(net1646),
    .B1(_11546_),
    .Y(_04019_));
 sky130_fd_sc_hd__o21ai_0 _32375_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[28] ),
    .A2(net1646),
    .B1(net2105),
    .Y(_11549_));
 sky130_fd_sc_hd__a21oi_1 _32376_ (.A1(_05840_),
    .A2(net1646),
    .B1(_11549_),
    .Y(_04020_));
 sky130_fd_sc_hd__o21ai_0 _32377_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[29] ),
    .A2(net1645),
    .B1(net2104),
    .Y(_11550_));
 sky130_fd_sc_hd__a21oi_1 _32378_ (.A1(_05853_),
    .A2(net1645),
    .B1(_11550_),
    .Y(_04021_));
 sky130_fd_sc_hd__o21ai_0 _32380_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[30] ),
    .A2(net1648),
    .B1(net2097),
    .Y(_11552_));
 sky130_fd_sc_hd__a21oi_1 _32381_ (.A1(_05866_),
    .A2(net1644),
    .B1(_11552_),
    .Y(_04022_));
 sky130_fd_sc_hd__o21ai_0 _32382_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[31] ),
    .A2(net1641),
    .B1(net2032),
    .Y(_11553_));
 sky130_fd_sc_hd__a21oi_1 _32383_ (.A1(_05880_),
    .A2(net1641),
    .B1(_11553_),
    .Y(_04023_));
 sky130_fd_sc_hd__o21ai_0 _32384_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[4] ),
    .A2(net1641),
    .B1(net2034),
    .Y(_11554_));
 sky130_fd_sc_hd__a21oi_1 _32385_ (.A1(_20548_),
    .A2(net1641),
    .B1(_11554_),
    .Y(_04024_));
 sky130_fd_sc_hd__o21ai_0 _32386_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[5] ),
    .A2(net1644),
    .B1(net2043),
    .Y(_11555_));
 sky130_fd_sc_hd__a21oi_1 _32387_ (.A1(_20575_),
    .A2(net1644),
    .B1(_11555_),
    .Y(_04025_));
 sky130_fd_sc_hd__o21ai_0 _32388_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[6] ),
    .A2(net1642),
    .B1(net2043),
    .Y(_11556_));
 sky130_fd_sc_hd__a21oi_1 _32389_ (.A1(_20603_),
    .A2(net1642),
    .B1(_11556_),
    .Y(_04026_));
 sky130_fd_sc_hd__inv_1 _32390_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[5] ),
    .Y(_11557_));
 sky130_fd_sc_hd__o21ai_0 _32391_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[7] ),
    .A2(net1641),
    .B1(net2084),
    .Y(_11558_));
 sky130_fd_sc_hd__a21oi_1 _32392_ (.A1(_11557_),
    .A2(net1641),
    .B1(_11558_),
    .Y(_04027_));
 sky130_fd_sc_hd__o21ai_0 _32393_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[8] ),
    .A2(net1643),
    .B1(net2045),
    .Y(_11559_));
 sky130_fd_sc_hd__a21oi_1 _32394_ (.A1(_20672_),
    .A2(net1643),
    .B1(_11559_),
    .Y(_04028_));
 sky130_fd_sc_hd__inv_1 _32395_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[7] ),
    .Y(_11560_));
 sky130_fd_sc_hd__o21ai_0 _32396_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[9] ),
    .A2(net1643),
    .B1(net2045),
    .Y(_11561_));
 sky130_fd_sc_hd__a21oi_1 _32397_ (.A1(_11560_),
    .A2(net1644),
    .B1(_11561_),
    .Y(_04029_));
 sky130_fd_sc_hd__o21ai_0 _32399_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[10] ),
    .A2(net1643),
    .B1(net2069),
    .Y(_11563_));
 sky130_fd_sc_hd__a21oi_1 _32400_ (.A1(_20714_),
    .A2(net1644),
    .B1(_11563_),
    .Y(_04030_));
 sky130_fd_sc_hd__o21ai_0 _32401_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[11] ),
    .A2(net1641),
    .B1(net2088),
    .Y(_11564_));
 sky130_fd_sc_hd__a21oi_1 _32402_ (.A1(_20737_),
    .A2(net1642),
    .B1(_11564_),
    .Y(_04031_));
 sky130_fd_sc_hd__o21ai_0 _32403_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[0] ),
    .A2(net1642),
    .B1(net2090),
    .Y(_11565_));
 sky130_fd_sc_hd__a21oi_1 _32404_ (.A1(_20388_),
    .A2(net1642),
    .B1(_11565_),
    .Y(_04032_));
 sky130_fd_sc_hd__o21ai_0 _32405_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[1] ),
    .A2(net1642),
    .B1(net2087),
    .Y(_11566_));
 sky130_fd_sc_hd__a21oi_1 _32406_ (.A1(_20438_),
    .A2(net1642),
    .B1(_11566_),
    .Y(_04033_));
 sky130_fd_sc_hd__o21ai_0 _32407_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mtvec_m_select ),
    .A2(net2222),
    .B1(net2085),
    .Y(_11567_));
 sky130_fd_sc_hd__a21oi_1 _32408_ (.A1(net2210),
    .A2(net2221),
    .B1(_11567_),
    .Y(_04034_));
 sky130_fd_sc_hd__inv_1 _32409_ (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec_m_select ),
    .Y(_11568_));
 sky130_fd_sc_hd__o21ai_0 _32411_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mtvec_w_select ),
    .A2(net2251),
    .B1(net2085),
    .Y(_11570_));
 sky130_fd_sc_hd__a21oi_1 _32412_ (.A1(_11568_),
    .A2(net2221),
    .B1(_11570_),
    .Y(_04035_));
 sky130_fd_sc_hd__nor2_1 _32413_ (.A(net2892),
    .B(net671),
    .Y(_11571_));
 sky130_fd_sc_hd__nor2_1 _32414_ (.A(net884),
    .B(_11184_),
    .Y(_11572_));
 sky130_fd_sc_hd__nand3_1 _32415_ (.A(_11186_),
    .B(_11141_),
    .C(_11572_),
    .Y(_11573_));
 sky130_fd_sc_hd__nand2_1 _32416_ (.A(net671),
    .B(_11573_),
    .Y(_11574_));
 sky130_fd_sc_hd__nand2_1 _32417_ (.A(_11574_),
    .B(net2031),
    .Y(_11575_));
 sky130_fd_sc_hd__nor2_4 _32418_ (.A(_11571_),
    .B(_11575_),
    .Y(_04036_));
 sky130_fd_sc_hd__nor2_1 _32419_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.msie.x_data ),
    .B(net1884),
    .Y(_11576_));
 sky130_fd_sc_hd__o21ai_0 _32420_ (.A1(\inst$top.soc.cpu.exception.m_mie.msie ),
    .A2(net2222),
    .B1(net2086),
    .Y(_11577_));
 sky130_fd_sc_hd__nor2_1 _32421_ (.A(_11576_),
    .B(_11577_),
    .Y(_04037_));
 sky130_fd_sc_hd__o21ai_0 _32422_ (.A1(\inst$top.soc.cpu.exception.m_mie[10] ),
    .A2(net2258),
    .B1(net2100),
    .Y(_11578_));
 sky130_fd_sc_hd__a21oi_1 _32423_ (.A1(_05759_),
    .A2(net2258),
    .B1(_11578_),
    .Y(_04038_));
 sky130_fd_sc_hd__o21ai_0 _32425_ (.A1(\inst$top.soc.cpu.exception.m_mie[11] ),
    .A2(net2256),
    .B1(net2096),
    .Y(_11580_));
 sky130_fd_sc_hd__a21oi_1 _32426_ (.A1(_05776_),
    .A2(net2256),
    .B1(_11580_),
    .Y(_04039_));
 sky130_fd_sc_hd__o21ai_0 _32427_ (.A1(\inst$top.soc.cpu.exception.m_mie[12] ),
    .A2(net2253),
    .B1(net2090),
    .Y(_11581_));
 sky130_fd_sc_hd__a21oi_1 _32428_ (.A1(_05796_),
    .A2(net2253),
    .B1(_11581_),
    .Y(_04040_));
 sky130_fd_sc_hd__o21ai_0 _32429_ (.A1(\inst$top.soc.cpu.exception.m_mie[13] ),
    .A2(net2256),
    .B1(net2100),
    .Y(_11582_));
 sky130_fd_sc_hd__a21oi_1 _32430_ (.A1(_05815_),
    .A2(net2257),
    .B1(_11582_),
    .Y(_04041_));
 sky130_fd_sc_hd__o21ai_0 _32433_ (.A1(\inst$top.soc.cpu.exception.m_mie[14] ),
    .A2(net2256),
    .B1(net2095),
    .Y(_11585_));
 sky130_fd_sc_hd__a21oi_1 _32434_ (.A1(_05828_),
    .A2(net2256),
    .B1(_11585_),
    .Y(_04042_));
 sky130_fd_sc_hd__o21ai_0 _32435_ (.A1(\inst$top.soc.cpu.exception.m_mie[15] ),
    .A2(net2233),
    .B1(net2095),
    .Y(_11586_));
 sky130_fd_sc_hd__a21oi_1 _32436_ (.A1(_05841_),
    .A2(net2233),
    .B1(_11586_),
    .Y(_04043_));
 sky130_fd_sc_hd__o21ai_0 _32437_ (.A1(\inst$top.soc.cpu.exception.m_mie[16] ),
    .A2(net2233),
    .B1(net2095),
    .Y(_11587_));
 sky130_fd_sc_hd__a21oi_1 _32438_ (.A1(_05854_),
    .A2(net2233),
    .B1(_11587_),
    .Y(_04044_));
 sky130_fd_sc_hd__o21ai_0 _32439_ (.A1(\inst$top.soc.cpu.exception.m_mie[17] ),
    .A2(net2233),
    .B1(net2096),
    .Y(_11588_));
 sky130_fd_sc_hd__a21oi_1 _32440_ (.A1(_05863_),
    .A2(net2233),
    .B1(_11588_),
    .Y(_04045_));
 sky130_fd_sc_hd__nor2_1 _32441_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[15] ),
    .B(net1884),
    .Y(_11589_));
 sky130_fd_sc_hd__o21ai_0 _32442_ (.A1(\inst$top.soc.cpu.exception.m_mie[18] ),
    .A2(net2251),
    .B1(net2085),
    .Y(_11590_));
 sky130_fd_sc_hd__nor2_1 _32443_ (.A(_11589_),
    .B(_11590_),
    .Y(_04046_));
 sky130_fd_sc_hd__nor2_1 _32445_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mtie.x_data ),
    .B(net1884),
    .Y(_11592_));
 sky130_fd_sc_hd__o21ai_0 _32447_ (.A1(\inst$top.soc.cpu.exception.m_mie.mtie ),
    .A2(net2222),
    .B1(net2086),
    .Y(_11594_));
 sky130_fd_sc_hd__nor2_1 _32448_ (.A(_11592_),
    .B(_11594_),
    .Y(_04047_));
 sky130_fd_sc_hd__nor2_1 _32449_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.meie.x_data ),
    .B(net1884),
    .Y(_11595_));
 sky130_fd_sc_hd__o21ai_0 _32450_ (.A1(\inst$top.soc.cpu.exception.m_mie.meie ),
    .A2(net2224),
    .B1(net2087),
    .Y(_11596_));
 sky130_fd_sc_hd__nor2_1 _32451_ (.A(_11595_),
    .B(_11596_),
    .Y(_04048_));
 sky130_fd_sc_hd__nor2_1 _32452_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[0] ),
    .B(net1884),
    .Y(_11597_));
 sky130_fd_sc_hd__o21ai_0 _32453_ (.A1(\inst$top.soc.cpu.exception.m_mie[3] ),
    .A2(net2222),
    .B1(net2085),
    .Y(_11598_));
 sky130_fd_sc_hd__nor2_1 _32454_ (.A(_11597_),
    .B(_11598_),
    .Y(_04049_));
 sky130_fd_sc_hd__o21ai_0 _32455_ (.A1(\inst$top.soc.cpu.exception.m_mie[4] ),
    .A2(net2255),
    .B1(net2101),
    .Y(_11599_));
 sky130_fd_sc_hd__a21oi_1 _32456_ (.A1(_05631_),
    .A2(net2255),
    .B1(_11599_),
    .Y(_04050_));
 sky130_fd_sc_hd__o21ai_0 _32458_ (.A1(\inst$top.soc.cpu.exception.m_mie[5] ),
    .A2(net2255),
    .B1(net2101),
    .Y(_11601_));
 sky130_fd_sc_hd__a21oi_1 _32459_ (.A1(_05652_),
    .A2(net2255),
    .B1(_11601_),
    .Y(_04051_));
 sky130_fd_sc_hd__o21ai_0 _32460_ (.A1(\inst$top.soc.cpu.exception.m_mie[6] ),
    .A2(net2255),
    .B1(net2098),
    .Y(_11602_));
 sky130_fd_sc_hd__a21oi_1 _32461_ (.A1(_05674_),
    .A2(net2255),
    .B1(_11602_),
    .Y(_04052_));
 sky130_fd_sc_hd__o21ai_0 _32463_ (.A1(\inst$top.soc.cpu.exception.m_mie[7] ),
    .A2(net2253),
    .B1(net2091),
    .Y(_11604_));
 sky130_fd_sc_hd__a21oi_1 _32464_ (.A1(_05699_),
    .A2(net2254),
    .B1(_11604_),
    .Y(_04053_));
 sky130_fd_sc_hd__o21ai_0 _32465_ (.A1(\inst$top.soc.cpu.exception.m_mie[8] ),
    .A2(net2231),
    .B1(net2094),
    .Y(_11605_));
 sky130_fd_sc_hd__a21oi_1 _32466_ (.A1(_05720_),
    .A2(net2231),
    .B1(_11605_),
    .Y(_04054_));
 sky130_fd_sc_hd__o21ai_0 _32467_ (.A1(\inst$top.soc.cpu.exception.m_mie[9] ),
    .A2(net2258),
    .B1(net2099),
    .Y(_11606_));
 sky130_fd_sc_hd__a21oi_1 _32468_ (.A1(_05738_),
    .A2(net2258),
    .B1(_11606_),
    .Y(_04055_));
 sky130_fd_sc_hd__o21ai_0 _32470_ (.A1(\inst$top.soc.cpu.exception.m_mip.msip ),
    .A2(net2224),
    .B1(net2088),
    .Y(_11608_));
 sky130_fd_sc_hd__a21oi_1 _32471_ (.A1(_20510_),
    .A2(net2224),
    .B1(_11608_),
    .Y(_04056_));
 sky130_fd_sc_hd__o21ai_0 _32472_ (.A1(\inst$top.soc.cpu.exception.m_mip[10] ),
    .A2(net2258),
    .B1(net2100),
    .Y(_11609_));
 sky130_fd_sc_hd__a21oi_1 _32473_ (.A1(_05755_),
    .A2(net2258),
    .B1(_11609_),
    .Y(_04057_));
 sky130_fd_sc_hd__nor2_1 _32474_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[8] ),
    .B(net1892),
    .Y(_11610_));
 sky130_fd_sc_hd__o21ai_0 _32475_ (.A1(\inst$top.soc.cpu.exception.m_mip[11] ),
    .A2(net2256),
    .B1(net2096),
    .Y(_11611_));
 sky130_fd_sc_hd__nor2_1 _32476_ (.A(_11610_),
    .B(_11611_),
    .Y(_04058_));
 sky130_fd_sc_hd__nor2_1 _32477_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[9] ),
    .B(net1893),
    .Y(_11612_));
 sky130_fd_sc_hd__o21ai_0 _32478_ (.A1(\inst$top.soc.cpu.exception.m_mip[12] ),
    .A2(net2253),
    .B1(net2090),
    .Y(_11613_));
 sky130_fd_sc_hd__nor2_1 _32479_ (.A(_11612_),
    .B(_11613_),
    .Y(_04059_));
 sky130_fd_sc_hd__nor2_1 _32480_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[10] ),
    .B(net1893),
    .Y(_11614_));
 sky130_fd_sc_hd__o21ai_0 _32481_ (.A1(\inst$top.soc.cpu.exception.m_mip[13] ),
    .A2(net2257),
    .B1(net2099),
    .Y(_11615_));
 sky130_fd_sc_hd__nor2_1 _32482_ (.A(_11614_),
    .B(_11615_),
    .Y(_04060_));
 sky130_fd_sc_hd__nor2_1 _32483_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[11] ),
    .B(net1891),
    .Y(_11616_));
 sky130_fd_sc_hd__o21ai_0 _32485_ (.A1(\inst$top.soc.cpu.exception.m_mip[14] ),
    .A2(net2257),
    .B1(net2096),
    .Y(_11618_));
 sky130_fd_sc_hd__nor2_1 _32486_ (.A(_11616_),
    .B(_11618_),
    .Y(_04061_));
 sky130_fd_sc_hd__nor2_1 _32487_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[12] ),
    .B(net1891),
    .Y(_11619_));
 sky130_fd_sc_hd__o21ai_0 _32488_ (.A1(\inst$top.soc.cpu.exception.m_mip[15] ),
    .A2(net2257),
    .B1(net2095),
    .Y(_11620_));
 sky130_fd_sc_hd__nor2_1 _32489_ (.A(_11619_),
    .B(_11620_),
    .Y(_04062_));
 sky130_fd_sc_hd__o21ai_0 _32490_ (.A1(\inst$top.soc.cpu.exception.m_mip[16] ),
    .A2(net2234),
    .B1(net2095),
    .Y(_11621_));
 sky130_fd_sc_hd__a21oi_1 _32491_ (.A1(_05851_),
    .A2(net2234),
    .B1(_11621_),
    .Y(_04063_));
 sky130_fd_sc_hd__nor2_1 _32492_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[14] ),
    .B(net1891),
    .Y(_11622_));
 sky130_fd_sc_hd__o21ai_0 _32493_ (.A1(\inst$top.soc.cpu.exception.m_mip[17] ),
    .A2(net2233),
    .B1(net2096),
    .Y(_11623_));
 sky130_fd_sc_hd__nor2_1 _32494_ (.A(_11622_),
    .B(_11623_),
    .Y(_04064_));
 sky130_fd_sc_hd__nor2_1 _32495_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[15] ),
    .B(net1884),
    .Y(_11624_));
 sky130_fd_sc_hd__o21ai_0 _32496_ (.A1(\inst$top.soc.cpu.exception.m_mip[18] ),
    .A2(net2251),
    .B1(net2086),
    .Y(_11625_));
 sky130_fd_sc_hd__nor2_1 _32497_ (.A(_11624_),
    .B(_11625_),
    .Y(_04065_));
 sky130_fd_sc_hd__o21ai_0 _32498_ (.A1(\inst$top.soc.cpu.exception.m_mip.mtip ),
    .A2(net2224),
    .B1(net2087),
    .Y(_11626_));
 sky130_fd_sc_hd__a21oi_1 _32499_ (.A1(_20631_),
    .A2(net2224),
    .B1(_11626_),
    .Y(_04066_));
 sky130_fd_sc_hd__o21ai_0 _32500_ (.A1(\inst$top.soc.cpu.exception.m_mip.meip ),
    .A2(net2224),
    .B1(net2087),
    .Y(_11627_));
 sky130_fd_sc_hd__a21oi_1 _32501_ (.A1(_20735_),
    .A2(net2224),
    .B1(_11627_),
    .Y(_04067_));
 sky130_fd_sc_hd__o21ai_0 _32503_ (.A1(\inst$top.soc.cpu.exception.m_mip[3] ),
    .A2(net2224),
    .B1(net2087),
    .Y(_11629_));
 sky130_fd_sc_hd__a21oi_1 _32504_ (.A1(_05608_),
    .A2(net2224),
    .B1(_11629_),
    .Y(_04068_));
 sky130_fd_sc_hd__nor2_1 _32506_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[1] ),
    .B(net1909),
    .Y(_11631_));
 sky130_fd_sc_hd__o21ai_0 _32508_ (.A1(\inst$top.soc.cpu.exception.m_mip[4] ),
    .A2(net2259),
    .B1(net2101),
    .Y(_11633_));
 sky130_fd_sc_hd__nor2_1 _32509_ (.A(_11631_),
    .B(_11633_),
    .Y(_04069_));
 sky130_fd_sc_hd__nor2_1 _32510_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[2] ),
    .B(net1893),
    .Y(_11634_));
 sky130_fd_sc_hd__o21ai_0 _32511_ (.A1(\inst$top.soc.cpu.exception.m_mip[5] ),
    .A2(net2254),
    .B1(net2091),
    .Y(_11635_));
 sky130_fd_sc_hd__nor2_1 _32512_ (.A(_11634_),
    .B(_11635_),
    .Y(_04070_));
 sky130_fd_sc_hd__nor2_1 _32513_ (.A(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[3] ),
    .B(net1893),
    .Y(_11636_));
 sky130_fd_sc_hd__o21ai_0 _32514_ (.A1(\inst$top.soc.cpu.exception.m_mip[6] ),
    .A2(net2259),
    .B1(net2098),
    .Y(_11637_));
 sky130_fd_sc_hd__nor2_1 _32515_ (.A(_11636_),
    .B(_11637_),
    .Y(_04071_));
 sky130_fd_sc_hd__o21ai_0 _32516_ (.A1(\inst$top.soc.cpu.exception.m_mip[7] ),
    .A2(net2254),
    .B1(net2091),
    .Y(_11638_));
 sky130_fd_sc_hd__a21oi_1 _32517_ (.A1(_05696_),
    .A2(net2253),
    .B1(_11638_),
    .Y(_04072_));
 sky130_fd_sc_hd__o21ai_0 _32519_ (.A1(\inst$top.soc.cpu.exception.m_mip[8] ),
    .A2(net2231),
    .B1(net2094),
    .Y(_11640_));
 sky130_fd_sc_hd__a21oi_1 _32520_ (.A1(_05716_),
    .A2(net2231),
    .B1(_11640_),
    .Y(_04073_));
 sky130_fd_sc_hd__o21ai_0 _32521_ (.A1(\inst$top.soc.cpu.exception.m_mip[9] ),
    .A2(net2258),
    .B1(net2099),
    .Y(_11641_));
 sky130_fd_sc_hd__a21oi_1 _32522_ (.A1(_05735_),
    .A2(net2258),
    .B1(_11641_),
    .Y(_04074_));
 sky130_fd_sc_hd__inv_1 _32523_ (.A(net2891),
    .Y(_11642_));
 sky130_fd_sc_hd__o21ai_0 _32528_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mstatus.mie.x_data ),
    .A2(net1884),
    .B1(net2083),
    .Y(_11647_));
 sky130_fd_sc_hd__a21oi_1 _32529_ (.A1(_11642_),
    .A2(net1885),
    .B1(_11647_),
    .Y(_04075_));
 sky130_fd_sc_hd__o21ai_0 _32531_ (.A1(\inst$top.soc.cpu.exception.m_mstatus.mpie ),
    .A2(net2221),
    .B1(net2084),
    .Y(_11649_));
 sky130_fd_sc_hd__a21oi_1 _32532_ (.A1(_20636_),
    .A2(net2220),
    .B1(_11649_),
    .Y(_04076_));
 sky130_fd_sc_hd__o21ai_0 _32535_ (.A1(\inst$top.soc.cpu.exception.w_data$48[0] ),
    .A2(net2254),
    .B1(net2089),
    .Y(_11652_));
 sky130_fd_sc_hd__inv_1 _32536_ (.A(_20142_),
    .Y(_11653_));
 sky130_fd_sc_hd__nor2_1 _32537_ (.A(_20141_),
    .B(_20148_),
    .Y(_11654_));
 sky130_fd_sc_hd__o221ai_1 _32538_ (.A1(_11653_),
    .A2(_20143_),
    .B1(_20152_),
    .B2(_20203_),
    .C1(_11654_),
    .Y(_11655_));
 sky130_fd_sc_hd__nand2_1 _32539_ (.A(_11654_),
    .B(_20142_),
    .Y(_11656_));
 sky130_fd_sc_hd__inv_1 _32540_ (.A(_20153_),
    .Y(_11657_));
 sky130_fd_sc_hd__a31oi_1 _32541_ (.A1(_20143_),
    .A2(_11657_),
    .A3(_20154_),
    .B1(_11656_),
    .Y(_11658_));
 sky130_fd_sc_hd__nor2_1 _32542_ (.A(_11656_),
    .B(_11658_),
    .Y(_11659_));
 sky130_fd_sc_hd__inv_1 _32543_ (.A(_11659_),
    .Y(_11660_));
 sky130_fd_sc_hd__nor2_1 _32544_ (.A(_20205_),
    .B(_11660_),
    .Y(_11661_));
 sky130_fd_sc_hd__inv_1 _32545_ (.A(_11661_),
    .Y(_11662_));
 sky130_fd_sc_hd__nor2_1 _32546_ (.A(_20159_),
    .B(_11662_),
    .Y(_11663_));
 sky130_fd_sc_hd__inv_1 _32547_ (.A(_11663_),
    .Y(_11664_));
 sky130_fd_sc_hd__nor4_1 _32548_ (.A(_20207_),
    .B(_20208_),
    .C(_20169_),
    .D(_20216_),
    .Y(_11665_));
 sky130_fd_sc_hd__nand2_1 _32549_ (.A(_11661_),
    .B(_11665_),
    .Y(_11666_));
 sky130_fd_sc_hd__nand2_1 _32550_ (.A(_11664_),
    .B(_11666_),
    .Y(_11667_));
 sky130_fd_sc_hd__o21ai_0 _32551_ (.A1(_20155_),
    .A2(_11660_),
    .B1(_20199_),
    .Y(_11668_));
 sky130_fd_sc_hd__or3_1 _32552_ (.A(_20207_),
    .B(_20163_),
    .C(_11662_),
    .X(_11669_));
 sky130_fd_sc_hd__inv_1 _32553_ (.A(_20171_),
    .Y(_11670_));
 sky130_fd_sc_hd__inv_1 _32554_ (.A(_20211_),
    .Y(_11671_));
 sky130_fd_sc_hd__nor3_1 _32555_ (.A(_20214_),
    .B(_20175_),
    .C(_11671_),
    .Y(_11672_));
 sky130_fd_sc_hd__a21oi_1 _32556_ (.A1(_11670_),
    .A2(_20211_),
    .B1(_11672_),
    .Y(_11673_));
 sky130_fd_sc_hd__nand4_1 _32557_ (.A(_11669_),
    .B(_20218_),
    .C(net2231),
    .D(_11673_),
    .Y(_11674_));
 sky130_fd_sc_hd__nor4_1 _32558_ (.A(_11655_),
    .B(_11667_),
    .C(_11668_),
    .D(_11674_),
    .Y(_11675_));
 sky130_fd_sc_hd__nor2_1 _32559_ (.A(_11652_),
    .B(_11675_),
    .Y(_04077_));
 sky130_fd_sc_hd__o21ai_0 _32560_ (.A1(_11657_),
    .A2(_20150_),
    .B1(_11654_),
    .Y(_11676_));
 sky130_fd_sc_hd__nor2_1 _32561_ (.A(_20155_),
    .B(_11660_),
    .Y(_11677_));
 sky130_fd_sc_hd__nor3_1 _32562_ (.A(_20158_),
    .B(_11660_),
    .C(_11677_),
    .Y(_11678_));
 sky130_fd_sc_hd__a2111oi_0 _32563_ (.A1(_20167_),
    .A2(_20193_),
    .B1(_11676_),
    .C1(_11678_),
    .D1(_11667_),
    .Y(_11679_));
 sky130_fd_sc_hd__nor4_1 _32565_ (.A(_20168_),
    .B(_20178_),
    .C(_20150_),
    .D(_20166_),
    .Y(_11681_));
 sky130_fd_sc_hd__a21oi_1 _32566_ (.A1(net1381),
    .A2(_20173_),
    .B1(_11681_),
    .Y(_11682_));
 sky130_fd_sc_hd__o21ai_0 _32568_ (.A1(\inst$top.soc.cpu.exception.w_data$48[1] ),
    .A2(net2225),
    .B1(net2087),
    .Y(_11684_));
 sky130_fd_sc_hd__a41oi_1 _32569_ (.A1(_11679_),
    .A2(_20252_),
    .A3(net2236),
    .A4(_11682_),
    .B1(_11684_),
    .Y(_04078_));
 sky130_fd_sc_hd__nor2_1 _32572_ (.A(_11670_),
    .B(_11671_),
    .Y(_11687_));
 sky130_fd_sc_hd__inv_1 _32573_ (.A(_11687_),
    .Y(_11688_));
 sky130_fd_sc_hd__nor2_1 _32574_ (.A(_20174_),
    .B(_11688_),
    .Y(_11689_));
 sky130_fd_sc_hd__nand4_1 _32575_ (.A(_20146_),
    .B(net2891),
    .C(\inst$top.soc.cpu.exception.m_mip.mtip ),
    .D(\inst$top.soc.cpu.exception.m_mie.mtie ),
    .Y(_11690_));
 sky130_fd_sc_hd__nor2_1 _32576_ (.A(_11677_),
    .B(_11678_),
    .Y(_11691_));
 sky130_fd_sc_hd__o311ai_0 _32577_ (.A1(_20150_),
    .A2(_20153_),
    .A3(_20154_),
    .B1(_11690_),
    .C1(_11691_),
    .Y(_11692_));
 sky130_fd_sc_hd__nor3_1 _32578_ (.A(_11689_),
    .B(_11667_),
    .C(_11692_),
    .Y(_11693_));
 sky130_fd_sc_hd__or2_2 _32579_ (.A(_11672_),
    .B(_11681_),
    .X(_11694_));
 sky130_fd_sc_hd__nor2_1 _32580_ (.A(net1885),
    .B(_11694_),
    .Y(_11695_));
 sky130_fd_sc_hd__nand3_1 _32581_ (.A(_11693_),
    .B(_20253_),
    .C(_11695_),
    .Y(_11696_));
 sky130_fd_sc_hd__o211ai_1 _32582_ (.A1(\inst$top.soc.cpu.exception.w_data$48[2] ),
    .A2(net2225),
    .B1(net2088),
    .C1(_11696_),
    .Y(_11697_));
 sky130_fd_sc_hd__inv_2 _32583_ (.A(_11697_),
    .Y(_04079_));
 sky130_fd_sc_hd__nand2_1 _32584_ (.A(_20225_),
    .B(net2217),
    .Y(_11698_));
 sky130_fd_sc_hd__o211ai_1 _32585_ (.A1(\inst$top.soc.cpu.exception.w_data$48[31] ),
    .A2(net2216),
    .B1(net2032),
    .C1(_11698_),
    .Y(_11699_));
 sky130_fd_sc_hd__inv_2 _32586_ (.A(_11699_),
    .Y(_04080_));
 sky130_fd_sc_hd__nand2_1 _32587_ (.A(net1381),
    .B(_20173_),
    .Y(_11700_));
 sky130_fd_sc_hd__nand3b_1 _32588_ (.A_N(_11689_),
    .B(_11669_),
    .C(_11700_),
    .Y(_11701_));
 sky130_fd_sc_hd__nor2_1 _32589_ (.A(_20251_),
    .B(_11701_),
    .Y(_11702_));
 sky130_fd_sc_hd__nand3b_1 _32590_ (.A_N(_20162_),
    .B(_11661_),
    .C(_20159_),
    .Y(_11703_));
 sky130_fd_sc_hd__o21a_1 _32591_ (.A1(_20148_),
    .A2(_20140_),
    .B1(_11703_),
    .X(_11704_));
 sky130_fd_sc_hd__nand4_1 _32592_ (.A(_11702_),
    .B(_11666_),
    .C(_11695_),
    .D(_11704_),
    .Y(_11705_));
 sky130_fd_sc_hd__o211ai_1 _32593_ (.A1(\inst$top.soc.cpu.exception.w_data$48[3] ),
    .A2(net2225),
    .B1(net2089),
    .C1(_11705_),
    .Y(_11706_));
 sky130_fd_sc_hd__inv_2 _32594_ (.A(_11706_),
    .Y(_04081_));
 sky130_fd_sc_hd__nand3_1 _32595_ (.A(_11691_),
    .B(_11664_),
    .C(_11703_),
    .Y(_11707_));
 sky130_fd_sc_hd__nor2_1 _32596_ (.A(_11658_),
    .B(_11694_),
    .Y(_11708_));
 sky130_fd_sc_hd__nand2_1 _32597_ (.A(_11654_),
    .B(_11653_),
    .Y(_11709_));
 sky130_fd_sc_hd__nand3_1 _32598_ (.A(_11708_),
    .B(_11709_),
    .C(_11666_),
    .Y(_11710_));
 sky130_fd_sc_hd__nor3_1 _32599_ (.A(_11707_),
    .B(_11710_),
    .C(_11701_),
    .Y(_11711_));
 sky130_fd_sc_hd__nand2_1 _32601_ (.A(_11711_),
    .B(net2225),
    .Y(_11713_));
 sky130_fd_sc_hd__o211ai_1 _32602_ (.A1(\inst$top.soc.cpu.exception.w_data$48[4] ),
    .A2(net2225),
    .B1(net2034),
    .C1(_11713_),
    .Y(_11714_));
 sky130_fd_sc_hd__inv_2 _32603_ (.A(_11714_),
    .Y(_04082_));
 sky130_fd_sc_hd__inv_1 _32605_ (.A(net1019),
    .Y(_11716_));
 sky130_fd_sc_hd__nand2_1 _32606_ (.A(_11716_),
    .B(\inst$top.soc.cpu.sink__payload$18[180] ),
    .Y(_11717_));
 sky130_fd_sc_hd__nand2_1 _32608_ (.A(net1069),
    .B(\inst$top.soc.cpu.sink__payload$18[109] ),
    .Y(_11719_));
 sky130_fd_sc_hd__nand3_1 _32609_ (.A(net1381),
    .B(_20219_),
    .C(\inst$top.soc.cpu.sink__payload$18[32] ),
    .Y(_11720_));
 sky130_fd_sc_hd__o21ai_0 _32610_ (.A1(\inst$top.soc.cpu.exception.w_data$51[0] ),
    .A2(net2229),
    .B1(net2043),
    .Y(_11721_));
 sky130_fd_sc_hd__a41oi_1 _32611_ (.A1(_11717_),
    .A2(_11719_),
    .A3(net2228),
    .A4(_11720_),
    .B1(_11721_),
    .Y(_04083_));
 sky130_fd_sc_hd__inv_1 _32612_ (.A(_20218_),
    .Y(_11722_));
 sky130_fd_sc_hd__inv_2 _32614_ (.A(\inst$top.soc.cpu.sink__payload$18[102] ),
    .Y(_11724_));
 sky130_fd_sc_hd__inv_1 _32617_ (.A(\inst$top.soc.cpu.sink__payload$18[190] ),
    .Y(_11727_));
 sky130_fd_sc_hd__o22ai_1 _32618_ (.A1(_11724_),
    .A2(net1193),
    .B1(_11727_),
    .B2(net1020),
    .Y(_11728_));
 sky130_fd_sc_hd__a221oi_1 _32619_ (.A1(\inst$top.soc.cpu.sink__payload$18[10] ),
    .A2(net1028),
    .B1(\inst$top.soc.cpu.sink__payload$18[119] ),
    .B2(net1070),
    .C1(_11728_),
    .Y(_11729_));
 sky130_fd_sc_hd__o21ai_0 _32620_ (.A1(\inst$top.soc.cpu.exception.w_data$51[10] ),
    .A2(net2240),
    .B1(net2070),
    .Y(_11730_));
 sky130_fd_sc_hd__a21oi_1 _32621_ (.A1(_11729_),
    .A2(net2240),
    .B1(_11730_),
    .Y(_04084_));
 sky130_fd_sc_hd__inv_1 _32622_ (.A(\inst$top.soc.cpu.sink__payload$18[191] ),
    .Y(_11731_));
 sky130_fd_sc_hd__o22ai_1 _32623_ (.A1(_20271_),
    .A2(net1195),
    .B1(_11731_),
    .B2(net1019),
    .Y(_11732_));
 sky130_fd_sc_hd__a221oi_1 _32624_ (.A1(\inst$top.soc.cpu.sink__payload$18[11] ),
    .A2(net1027),
    .B1(\inst$top.soc.cpu.sink__payload$18[120] ),
    .B2(net1068),
    .C1(_11732_),
    .Y(_11733_));
 sky130_fd_sc_hd__o21ai_0 _32625_ (.A1(\inst$top.soc.cpu.exception.w_data$51[11] ),
    .A2(net2230),
    .B1(net2093),
    .Y(_11734_));
 sky130_fd_sc_hd__a21oi_1 _32626_ (.A1(_11733_),
    .A2(net2230),
    .B1(_11734_),
    .Y(_04085_));
 sky130_fd_sc_hd__inv_2 _32627_ (.A(\inst$top.soc.cpu.sink__payload$18[106] ),
    .Y(_11735_));
 sky130_fd_sc_hd__inv_1 _32628_ (.A(\inst$top.soc.cpu.sink__payload$18[192] ),
    .Y(_11736_));
 sky130_fd_sc_hd__o22ai_1 _32629_ (.A1(_11735_),
    .A2(net1194),
    .B1(_11736_),
    .B2(net1021),
    .Y(_11737_));
 sky130_fd_sc_hd__a221oi_1 _32630_ (.A1(\inst$top.soc.cpu.sink__payload$18[12] ),
    .A2(net1029),
    .B1(\inst$top.soc.cpu.sink__payload$18[121] ),
    .B2(net1071),
    .C1(_11737_),
    .Y(_11738_));
 sky130_fd_sc_hd__o21ai_0 _32631_ (.A1(\inst$top.soc.cpu.exception.w_data$51[12] ),
    .A2(net2232),
    .B1(net2097),
    .Y(_11739_));
 sky130_fd_sc_hd__a21oi_1 _32632_ (.A1(_11738_),
    .A2(net2232),
    .B1(_11739_),
    .Y(_04086_));
 sky130_fd_sc_hd__inv_1 _32633_ (.A(\inst$top.soc.cpu.sink__payload$18[107] ),
    .Y(_11740_));
 sky130_fd_sc_hd__inv_1 _32634_ (.A(\inst$top.soc.cpu.sink__payload$18[193] ),
    .Y(_11741_));
 sky130_fd_sc_hd__o22ai_1 _32635_ (.A1(_11740_),
    .A2(net1193),
    .B1(_11741_),
    .B2(net1020),
    .Y(_11742_));
 sky130_fd_sc_hd__a221oi_1 _32636_ (.A1(\inst$top.soc.cpu.sink__payload$18[13] ),
    .A2(net1028),
    .B1(\inst$top.soc.cpu.sink__payload$18[122] ),
    .B2(net1070),
    .C1(_11742_),
    .Y(_11743_));
 sky130_fd_sc_hd__o21ai_0 _32637_ (.A1(\inst$top.soc.cpu.exception.w_data$51[13] ),
    .A2(net2242),
    .B1(net2104),
    .Y(_11744_));
 sky130_fd_sc_hd__a21oi_1 _32638_ (.A1(_11743_),
    .A2(net2242),
    .B1(_11744_),
    .Y(_04087_));
 sky130_fd_sc_hd__inv_1 _32639_ (.A(\inst$top.soc.cpu.sink__payload$18[108] ),
    .Y(_11745_));
 sky130_fd_sc_hd__inv_1 _32640_ (.A(\inst$top.soc.cpu.sink__payload$18[194] ),
    .Y(_11746_));
 sky130_fd_sc_hd__o22ai_1 _32641_ (.A1(_11745_),
    .A2(net1193),
    .B1(_11746_),
    .B2(net1020),
    .Y(_11747_));
 sky130_fd_sc_hd__a221oi_1 _32642_ (.A1(\inst$top.soc.cpu.sink__payload$18[14] ),
    .A2(net1028),
    .B1(\inst$top.soc.cpu.sink__payload$18[123] ),
    .B2(net1070),
    .C1(_11747_),
    .Y(_11748_));
 sky130_fd_sc_hd__o21ai_0 _32643_ (.A1(\inst$top.soc.cpu.exception.w_data$51[14] ),
    .A2(net2239),
    .B1(net2069),
    .Y(_11749_));
 sky130_fd_sc_hd__a21oi_1 _32644_ (.A1(_11748_),
    .A2(net2239),
    .B1(_11749_),
    .Y(_04088_));
 sky130_fd_sc_hd__inv_1 _32645_ (.A(\inst$top.soc.cpu.sink__payload$18[47] ),
    .Y(_11750_));
 sky130_fd_sc_hd__inv_1 _32646_ (.A(\inst$top.soc.cpu.sink__payload$18[195] ),
    .Y(_11751_));
 sky130_fd_sc_hd__o22ai_1 _32647_ (.A1(_11750_),
    .A2(net1193),
    .B1(_11751_),
    .B2(net1020),
    .Y(_11752_));
 sky130_fd_sc_hd__a221oi_1 _32648_ (.A1(\inst$top.soc.cpu.sink__payload$18[15] ),
    .A2(net1028),
    .B1(\inst$top.soc.cpu.sink__payload$18[124] ),
    .B2(net1070),
    .C1(_11752_),
    .Y(_11753_));
 sky130_fd_sc_hd__o21ai_0 _32650_ (.A1(\inst$top.soc.cpu.exception.w_data$51[15] ),
    .A2(net2240),
    .B1(net2070),
    .Y(_11755_));
 sky130_fd_sc_hd__a21oi_1 _32651_ (.A1(_11753_),
    .A2(net2241),
    .B1(_11755_),
    .Y(_04089_));
 sky130_fd_sc_hd__inv_1 _32652_ (.A(\inst$top.soc.cpu.sink__payload$18[196] ),
    .Y(_11756_));
 sky130_fd_sc_hd__nand3_1 _32653_ (.A(net1381),
    .B(_20219_),
    .C(\inst$top.soc.cpu.sink__payload$18[48] ),
    .Y(_11757_));
 sky130_fd_sc_hd__o21ai_0 _32654_ (.A1(_11756_),
    .A2(net1021),
    .B1(_11757_),
    .Y(_11758_));
 sky130_fd_sc_hd__a221oi_1 _32655_ (.A1(\inst$top.soc.cpu.sink__payload$18[16] ),
    .A2(net1029),
    .B1(\inst$top.soc.cpu.sink__payload$18[125] ),
    .B2(net1071),
    .C1(_11758_),
    .Y(_11759_));
 sky130_fd_sc_hd__o21ai_0 _32656_ (.A1(\inst$top.soc.cpu.exception.w_data$51[16] ),
    .A2(net2232),
    .B1(net2097),
    .Y(_11760_));
 sky130_fd_sc_hd__a21oi_1 _32657_ (.A1(_11759_),
    .A2(net2232),
    .B1(_11760_),
    .Y(_04090_));
 sky130_fd_sc_hd__inv_1 _32659_ (.A(\inst$top.soc.cpu.sink__payload$18[49] ),
    .Y(_11762_));
 sky130_fd_sc_hd__inv_1 _32660_ (.A(\inst$top.soc.cpu.sink__payload$18[197] ),
    .Y(_11763_));
 sky130_fd_sc_hd__o22ai_1 _32661_ (.A1(_11762_),
    .A2(net1194),
    .B1(_11763_),
    .B2(net1021),
    .Y(_11764_));
 sky130_fd_sc_hd__a221oi_1 _32662_ (.A1(\inst$top.soc.cpu.sink__payload$18[17] ),
    .A2(net1029),
    .B1(\inst$top.soc.cpu.sink__payload$18[126] ),
    .B2(net1071),
    .C1(_11764_),
    .Y(_11765_));
 sky130_fd_sc_hd__o21ai_0 _32664_ (.A1(\inst$top.soc.cpu.exception.w_data$51[17] ),
    .A2(net2256),
    .B1(net2096),
    .Y(_11767_));
 sky130_fd_sc_hd__a21oi_1 _32665_ (.A1(_11765_),
    .A2(net2256),
    .B1(_11767_),
    .Y(_04091_));
 sky130_fd_sc_hd__inv_1 _32666_ (.A(\inst$top.soc.cpu.sink__payload$18[50] ),
    .Y(_11768_));
 sky130_fd_sc_hd__inv_1 _32667_ (.A(\inst$top.soc.cpu.sink__payload$18[198] ),
    .Y(_11769_));
 sky130_fd_sc_hd__o22ai_1 _32668_ (.A1(_11768_),
    .A2(net1195),
    .B1(_11769_),
    .B2(net1018),
    .Y(_11770_));
 sky130_fd_sc_hd__a221oi_1 _32669_ (.A1(\inst$top.soc.cpu.sink__payload$18[18] ),
    .A2(net1027),
    .B1(\inst$top.soc.cpu.sink__payload$18[127] ),
    .B2(net1069),
    .C1(_11770_),
    .Y(_11771_));
 sky130_fd_sc_hd__o21ai_0 _32670_ (.A1(\inst$top.soc.cpu.exception.w_data$51[18] ),
    .A2(net2255),
    .B1(net2094),
    .Y(_11772_));
 sky130_fd_sc_hd__a21oi_1 _32671_ (.A1(_11771_),
    .A2(net2256),
    .B1(_11772_),
    .Y(_04092_));
 sky130_fd_sc_hd__inv_1 _32673_ (.A(\inst$top.soc.cpu.sink__payload$18[51] ),
    .Y(_11774_));
 sky130_fd_sc_hd__inv_1 _32674_ (.A(\inst$top.soc.cpu.sink__payload$18[199] ),
    .Y(_11775_));
 sky130_fd_sc_hd__o22ai_1 _32675_ (.A1(_11774_),
    .A2(net1195),
    .B1(_11775_),
    .B2(net1018),
    .Y(_11776_));
 sky130_fd_sc_hd__a221oi_1 _32676_ (.A1(\inst$top.soc.cpu.sink__payload$18[19] ),
    .A2(net1030),
    .B1(\inst$top.soc.cpu.sink__payload$18[128] ),
    .B2(net1069),
    .C1(_11776_),
    .Y(_11777_));
 sky130_fd_sc_hd__o21ai_0 _32678_ (.A1(\inst$top.soc.cpu.exception.w_data$51[19] ),
    .A2(net2256),
    .B1(net2096),
    .Y(_11779_));
 sky130_fd_sc_hd__a21oi_1 _32679_ (.A1(_11777_),
    .A2(net2233),
    .B1(_11779_),
    .Y(_04093_));
 sky130_fd_sc_hd__a22oi_1 _32680_ (.A1(net1068),
    .A2(\inst$top.soc.cpu.sink__payload$18[110] ),
    .B1(_11716_),
    .B2(\inst$top.soc.cpu.sink__payload$18[181] ),
    .Y(_11780_));
 sky130_fd_sc_hd__nand3_1 _32682_ (.A(net1381),
    .B(_20219_),
    .C(\inst$top.soc.cpu.sink__payload$18[33] ),
    .Y(_11782_));
 sky130_fd_sc_hd__o21ai_0 _32683_ (.A1(\inst$top.soc.cpu.exception.w_data$51[1] ),
    .A2(net2227),
    .B1(net2043),
    .Y(_11783_));
 sky130_fd_sc_hd__a31oi_1 _32684_ (.A1(_11780_),
    .A2(net2227),
    .A3(_11782_),
    .B1(_11783_),
    .Y(_04094_));
 sky130_fd_sc_hd__inv_1 _32685_ (.A(\inst$top.soc.cpu.sink__payload$18[52] ),
    .Y(_11784_));
 sky130_fd_sc_hd__inv_1 _32686_ (.A(\inst$top.soc.cpu.sink__payload$18[200] ),
    .Y(_11785_));
 sky130_fd_sc_hd__o22ai_1 _32688_ (.A1(_11784_),
    .A2(net1192),
    .B1(_11785_),
    .B2(net1019),
    .Y(_11787_));
 sky130_fd_sc_hd__a221oi_1 _32689_ (.A1(\inst$top.soc.cpu.sink__payload$18[20] ),
    .A2(net1027),
    .B1(\inst$top.soc.cpu.sink__payload$18[129] ),
    .B2(net1069),
    .C1(_11787_),
    .Y(_11788_));
 sky130_fd_sc_hd__o21ai_0 _32690_ (.A1(\inst$top.soc.cpu.exception.w_data$51[20] ),
    .A2(net2255),
    .B1(net2094),
    .Y(_11789_));
 sky130_fd_sc_hd__a21oi_1 _32691_ (.A1(_11788_),
    .A2(net2255),
    .B1(_11789_),
    .Y(_04095_));
 sky130_fd_sc_hd__inv_1 _32692_ (.A(\inst$top.soc.cpu.sink__payload$18[53] ),
    .Y(_11790_));
 sky130_fd_sc_hd__inv_1 _32694_ (.A(\inst$top.soc.cpu.sink__payload$18[201] ),
    .Y(_11792_));
 sky130_fd_sc_hd__o22ai_1 _32695_ (.A1(_11790_),
    .A2(net1195),
    .B1(_11792_),
    .B2(net1019),
    .Y(_11793_));
 sky130_fd_sc_hd__a221oi_1 _32696_ (.A1(\inst$top.soc.cpu.sink__payload$18[21] ),
    .A2(net1027),
    .B1(\inst$top.soc.cpu.sink__payload$18[130] ),
    .B2(net1069),
    .C1(_11793_),
    .Y(_11794_));
 sky130_fd_sc_hd__o21ai_0 _32697_ (.A1(\inst$top.soc.cpu.exception.w_data$51[21] ),
    .A2(net2230),
    .B1(net2093),
    .Y(_11795_));
 sky130_fd_sc_hd__a21oi_1 _32698_ (.A1(_11794_),
    .A2(net2230),
    .B1(_11795_),
    .Y(_04096_));
 sky130_fd_sc_hd__inv_1 _32699_ (.A(\inst$top.soc.cpu.sink__payload$18[54] ),
    .Y(_11796_));
 sky130_fd_sc_hd__inv_1 _32700_ (.A(\inst$top.soc.cpu.sink__payload$18[202] ),
    .Y(_11797_));
 sky130_fd_sc_hd__o22ai_1 _32701_ (.A1(_11796_),
    .A2(net1194),
    .B1(_11797_),
    .B2(net1021),
    .Y(_11798_));
 sky130_fd_sc_hd__a221oi_1 _32702_ (.A1(\inst$top.soc.cpu.sink__payload$18[22] ),
    .A2(net1028),
    .B1(\inst$top.soc.cpu.sink__payload$18[131] ),
    .B2(net1070),
    .C1(_11798_),
    .Y(_11799_));
 sky130_fd_sc_hd__o21ai_0 _32703_ (.A1(\inst$top.soc.cpu.exception.w_data$51[22] ),
    .A2(net2262),
    .B1(net2105),
    .Y(_11800_));
 sky130_fd_sc_hd__a21oi_1 _32704_ (.A1(_11799_),
    .A2(net2262),
    .B1(_11800_),
    .Y(_04097_));
 sky130_fd_sc_hd__inv_1 _32705_ (.A(\inst$top.soc.cpu.sink__payload$18[55] ),
    .Y(_11801_));
 sky130_fd_sc_hd__inv_1 _32706_ (.A(\inst$top.soc.cpu.sink__payload$18[203] ),
    .Y(_11802_));
 sky130_fd_sc_hd__o22ai_1 _32707_ (.A1(_11801_),
    .A2(net1194),
    .B1(_11802_),
    .B2(net1020),
    .Y(_11803_));
 sky130_fd_sc_hd__a221oi_1 _32708_ (.A1(\inst$top.soc.cpu.sink__payload$18[23] ),
    .A2(net1028),
    .B1(\inst$top.soc.cpu.sink__payload$18[132] ),
    .B2(net1070),
    .C1(_11803_),
    .Y(_11804_));
 sky130_fd_sc_hd__o21ai_0 _32709_ (.A1(\inst$top.soc.cpu.exception.w_data$51[23] ),
    .A2(net2260),
    .B1(net2110),
    .Y(_11805_));
 sky130_fd_sc_hd__a21oi_1 _32710_ (.A1(_11804_),
    .A2(net2260),
    .B1(_11805_),
    .Y(_04098_));
 sky130_fd_sc_hd__inv_1 _32711_ (.A(\inst$top.soc.cpu.sink__payload$18[56] ),
    .Y(_11806_));
 sky130_fd_sc_hd__inv_1 _32712_ (.A(\inst$top.soc.cpu.sink__payload$18[204] ),
    .Y(_11807_));
 sky130_fd_sc_hd__o22ai_1 _32713_ (.A1(_11806_),
    .A2(net1193),
    .B1(_11807_),
    .B2(net1020),
    .Y(_11808_));
 sky130_fd_sc_hd__a221oi_1 _32714_ (.A1(\inst$top.soc.cpu.sink__payload$18[24] ),
    .A2(net1028),
    .B1(\inst$top.soc.cpu.sink__payload$18[133] ),
    .B2(net1070),
    .C1(_11808_),
    .Y(_11809_));
 sky130_fd_sc_hd__o21ai_0 _32715_ (.A1(\inst$top.soc.cpu.exception.w_data$51[24] ),
    .A2(net2242),
    .B1(net2104),
    .Y(_11810_));
 sky130_fd_sc_hd__a21oi_1 _32716_ (.A1(_11809_),
    .A2(net2242),
    .B1(_11810_),
    .Y(_04099_));
 sky130_fd_sc_hd__inv_1 _32717_ (.A(\inst$top.soc.cpu.sink__payload$18[57] ),
    .Y(_11811_));
 sky130_fd_sc_hd__inv_1 _32718_ (.A(\inst$top.soc.cpu.sink__payload$18[205] ),
    .Y(_11812_));
 sky130_fd_sc_hd__o22ai_1 _32719_ (.A1(_11811_),
    .A2(net1192),
    .B1(_11812_),
    .B2(net1018),
    .Y(_11813_));
 sky130_fd_sc_hd__a221oi_1 _32720_ (.A1(\inst$top.soc.cpu.sink__payload$18[25] ),
    .A2(net1027),
    .B1(\inst$top.soc.cpu.sink__payload$18[134] ),
    .B2(net1068),
    .C1(_11813_),
    .Y(_11814_));
 sky130_fd_sc_hd__o21ai_0 _32723_ (.A1(\inst$top.soc.cpu.exception.w_data$51[25] ),
    .A2(net2252),
    .B1(net2086),
    .Y(_11817_));
 sky130_fd_sc_hd__a21oi_1 _32724_ (.A1(_11814_),
    .A2(net2251),
    .B1(_11817_),
    .Y(_04100_));
 sky130_fd_sc_hd__inv_1 _32725_ (.A(\inst$top.soc.cpu.sink__payload$18[58] ),
    .Y(_11818_));
 sky130_fd_sc_hd__inv_1 _32726_ (.A(\inst$top.soc.cpu.sink__payload$18[206] ),
    .Y(_11819_));
 sky130_fd_sc_hd__o22ai_1 _32727_ (.A1(_11818_),
    .A2(net1193),
    .B1(_11819_),
    .B2(net1020),
    .Y(_11820_));
 sky130_fd_sc_hd__a221oi_1 _32728_ (.A1(\inst$top.soc.cpu.sink__payload$18[26] ),
    .A2(net1028),
    .B1(\inst$top.soc.cpu.sink__payload$18[135] ),
    .B2(net1070),
    .C1(_11820_),
    .Y(_11821_));
 sky130_fd_sc_hd__o21ai_0 _32729_ (.A1(\inst$top.soc.cpu.exception.w_data$51[26] ),
    .A2(net2260),
    .B1(net2106),
    .Y(_11822_));
 sky130_fd_sc_hd__a21oi_1 _32730_ (.A1(_11821_),
    .A2(net2260),
    .B1(_11822_),
    .Y(_04101_));
 sky130_fd_sc_hd__inv_1 _32732_ (.A(\inst$top.soc.cpu.sink__payload$18[59] ),
    .Y(_11824_));
 sky130_fd_sc_hd__inv_1 _32733_ (.A(\inst$top.soc.cpu.sink__payload$18[207] ),
    .Y(_11825_));
 sky130_fd_sc_hd__o22ai_1 _32734_ (.A1(_11824_),
    .A2(net1193),
    .B1(_11825_),
    .B2(net1020),
    .Y(_11826_));
 sky130_fd_sc_hd__a221oi_1 _32735_ (.A1(\inst$top.soc.cpu.sink__payload$18[27] ),
    .A2(net1028),
    .B1(\inst$top.soc.cpu.sink__payload$18[136] ),
    .B2(net1071),
    .C1(_11826_),
    .Y(_11827_));
 sky130_fd_sc_hd__o21ai_0 _32737_ (.A1(\inst$top.soc.cpu.exception.w_data$51[27] ),
    .A2(net2260),
    .B1(net2106),
    .Y(_11829_));
 sky130_fd_sc_hd__a21oi_1 _32738_ (.A1(_11827_),
    .A2(net2244),
    .B1(_11829_),
    .Y(_04102_));
 sky130_fd_sc_hd__inv_1 _32739_ (.A(\inst$top.soc.cpu.sink__payload$18[60] ),
    .Y(_11830_));
 sky130_fd_sc_hd__inv_1 _32740_ (.A(\inst$top.soc.cpu.sink__payload$18[208] ),
    .Y(_11831_));
 sky130_fd_sc_hd__o22ai_1 _32741_ (.A1(_11830_),
    .A2(net1193),
    .B1(_11831_),
    .B2(net1020),
    .Y(_11832_));
 sky130_fd_sc_hd__a221oi_1 _32742_ (.A1(\inst$top.soc.cpu.sink__payload$18[28] ),
    .A2(net1028),
    .B1(\inst$top.soc.cpu.sink__payload$18[137] ),
    .B2(net1071),
    .C1(_11832_),
    .Y(_11833_));
 sky130_fd_sc_hd__o21ai_0 _32743_ (.A1(\inst$top.soc.cpu.exception.w_data$51[28] ),
    .A2(net2246),
    .B1(net2105),
    .Y(_11834_));
 sky130_fd_sc_hd__a21oi_1 _32744_ (.A1(_11833_),
    .A2(net2246),
    .B1(_11834_),
    .Y(_04103_));
 sky130_fd_sc_hd__inv_1 _32746_ (.A(\inst$top.soc.cpu.sink__payload$18[61] ),
    .Y(_11836_));
 sky130_fd_sc_hd__inv_1 _32747_ (.A(\inst$top.soc.cpu.sink__payload$18[209] ),
    .Y(_11837_));
 sky130_fd_sc_hd__o22ai_1 _32748_ (.A1(_11836_),
    .A2(net1193),
    .B1(_11837_),
    .B2(net1020),
    .Y(_11838_));
 sky130_fd_sc_hd__a221oi_1 _32749_ (.A1(\inst$top.soc.cpu.sink__payload$18[29] ),
    .A2(net1029),
    .B1(\inst$top.soc.cpu.sink__payload$18[138] ),
    .B2(net1070),
    .C1(_11838_),
    .Y(_11839_));
 sky130_fd_sc_hd__o21ai_0 _32751_ (.A1(\inst$top.soc.cpu.exception.w_data$51[29] ),
    .A2(net2242),
    .B1(net2104),
    .Y(_11841_));
 sky130_fd_sc_hd__a21oi_1 _32752_ (.A1(_11839_),
    .A2(net2242),
    .B1(_11841_),
    .Y(_04104_));
 sky130_fd_sc_hd__inv_1 _32753_ (.A(\inst$top.soc.cpu.sink__payload$18[34] ),
    .Y(_11842_));
 sky130_fd_sc_hd__inv_1 _32754_ (.A(\inst$top.soc.cpu.sink__payload$18[182] ),
    .Y(_11843_));
 sky130_fd_sc_hd__o22ai_1 _32756_ (.A1(_11842_),
    .A2(net1192),
    .B1(_11843_),
    .B2(net1018),
    .Y(_11845_));
 sky130_fd_sc_hd__a221oi_1 _32757_ (.A1(\inst$top.soc.cpu.sink__payload$18[2] ),
    .A2(net1027),
    .B1(\inst$top.soc.cpu.sink__payload$18[111] ),
    .B2(net1068),
    .C1(_11845_),
    .Y(_11846_));
 sky130_fd_sc_hd__o21ai_0 _32758_ (.A1(\inst$top.soc.cpu.exception.w_data$51[2] ),
    .A2(net2218),
    .B1(net2034),
    .Y(_11847_));
 sky130_fd_sc_hd__a21oi_1 _32759_ (.A1(_11846_),
    .A2(net2218),
    .B1(_11847_),
    .Y(_04105_));
 sky130_fd_sc_hd__inv_1 _32760_ (.A(\inst$top.soc.cpu.sink__payload$18[62] ),
    .Y(_11848_));
 sky130_fd_sc_hd__inv_1 _32761_ (.A(\inst$top.soc.cpu.sink__payload$18[210] ),
    .Y(_11849_));
 sky130_fd_sc_hd__o22ai_1 _32762_ (.A1(_11848_),
    .A2(net1193),
    .B1(_11849_),
    .B2(net1021),
    .Y(_11850_));
 sky130_fd_sc_hd__a221oi_1 _32763_ (.A1(\inst$top.soc.cpu.sink__payload$18[30] ),
    .A2(net1029),
    .B1(\inst$top.soc.cpu.sink__payload$18[139] ),
    .B2(net1070),
    .C1(_11850_),
    .Y(_11851_));
 sky130_fd_sc_hd__o21ai_0 _32764_ (.A1(\inst$top.soc.cpu.exception.w_data$51[30] ),
    .A2(net2242),
    .B1(net2104),
    .Y(_11852_));
 sky130_fd_sc_hd__a21oi_1 _32765_ (.A1(_11851_),
    .A2(net2242),
    .B1(_11852_),
    .Y(_04106_));
 sky130_fd_sc_hd__inv_1 _32766_ (.A(\inst$top.soc.cpu.sink__payload$18[63] ),
    .Y(_11853_));
 sky130_fd_sc_hd__inv_1 _32767_ (.A(\inst$top.soc.cpu.sink__payload$18[211] ),
    .Y(_11854_));
 sky130_fd_sc_hd__o22ai_1 _32768_ (.A1(_11853_),
    .A2(net1192),
    .B1(_11854_),
    .B2(net1018),
    .Y(_11855_));
 sky130_fd_sc_hd__a221oi_1 _32769_ (.A1(\inst$top.soc.cpu.sink__payload$18[31] ),
    .A2(net1027),
    .B1(\inst$top.soc.cpu.sink__payload$18[140] ),
    .B2(net1068),
    .C1(_11855_),
    .Y(_11856_));
 sky130_fd_sc_hd__o21ai_0 _32770_ (.A1(\inst$top.soc.cpu.exception.w_data$51[31] ),
    .A2(net2216),
    .B1(net2031),
    .Y(_11857_));
 sky130_fd_sc_hd__a21oi_1 _32771_ (.A1(_11856_),
    .A2(net2216),
    .B1(_11857_),
    .Y(_04107_));
 sky130_fd_sc_hd__inv_1 _32772_ (.A(\inst$top.soc.cpu.sink__payload$18[183] ),
    .Y(_11858_));
 sky130_fd_sc_hd__nand3_1 _32773_ (.A(net1381),
    .B(_20219_),
    .C(\inst$top.soc.cpu.sink__payload$18[35] ),
    .Y(_11859_));
 sky130_fd_sc_hd__o21ai_0 _32774_ (.A1(_11858_),
    .A2(net1018),
    .B1(_11859_),
    .Y(_11860_));
 sky130_fd_sc_hd__a21oi_1 _32775_ (.A1(\inst$top.soc.cpu.sink__payload$18[112] ),
    .A2(net1068),
    .B1(_11860_),
    .Y(_11861_));
 sky130_fd_sc_hd__nand2_1 _32776_ (.A(net1027),
    .B(\inst$top.soc.cpu.sink__payload$18[3] ),
    .Y(_11862_));
 sky130_fd_sc_hd__o21ai_0 _32777_ (.A1(\inst$top.soc.cpu.exception.w_data$51[3] ),
    .A2(net2225),
    .B1(net2088),
    .Y(_11863_));
 sky130_fd_sc_hd__a31oi_1 _32778_ (.A1(_11861_),
    .A2(net2217),
    .A3(_11862_),
    .B1(_11863_),
    .Y(_04108_));
 sky130_fd_sc_hd__inv_1 _32779_ (.A(\inst$top.soc.cpu.sink__payload$18[36] ),
    .Y(_11864_));
 sky130_fd_sc_hd__inv_1 _32780_ (.A(\inst$top.soc.cpu.sink__payload$18[184] ),
    .Y(_11865_));
 sky130_fd_sc_hd__o22ai_1 _32781_ (.A1(_11864_),
    .A2(net1192),
    .B1(_11865_),
    .B2(net1018),
    .Y(_11866_));
 sky130_fd_sc_hd__a221oi_1 _32782_ (.A1(\inst$top.soc.cpu.sink__payload$18[4] ),
    .A2(net1027),
    .B1(\inst$top.soc.cpu.sink__payload$18[113] ),
    .B2(net1068),
    .C1(_11866_),
    .Y(_11867_));
 sky130_fd_sc_hd__o21ai_0 _32783_ (.A1(\inst$top.soc.cpu.exception.w_data$51[4] ),
    .A2(net2217),
    .B1(net2033),
    .Y(_11868_));
 sky130_fd_sc_hd__a21oi_1 _32784_ (.A1(_11867_),
    .A2(net2217),
    .B1(_11868_),
    .Y(_04109_));
 sky130_fd_sc_hd__inv_1 _32785_ (.A(\inst$top.soc.cpu.sink__payload$18[37] ),
    .Y(_11869_));
 sky130_fd_sc_hd__inv_1 _32786_ (.A(\inst$top.soc.cpu.sink__payload$18[185] ),
    .Y(_11870_));
 sky130_fd_sc_hd__o22ai_1 _32787_ (.A1(_11869_),
    .A2(net1192),
    .B1(_11870_),
    .B2(net1019),
    .Y(_11871_));
 sky130_fd_sc_hd__a221oi_1 _32788_ (.A1(\inst$top.soc.cpu.sink__payload$18[5] ),
    .A2(net1030),
    .B1(\inst$top.soc.cpu.sink__payload$18[114] ),
    .B2(net1069),
    .C1(_11871_),
    .Y(_11872_));
 sky130_fd_sc_hd__o21ai_0 _32789_ (.A1(\inst$top.soc.cpu.exception.w_data$51[5] ),
    .A2(net2226),
    .B1(net2043),
    .Y(_11873_));
 sky130_fd_sc_hd__a21oi_1 _32790_ (.A1(_11872_),
    .A2(net2226),
    .B1(_11873_),
    .Y(_04110_));
 sky130_fd_sc_hd__inv_1 _32791_ (.A(\inst$top.soc.cpu.sink__payload$18[38] ),
    .Y(_11874_));
 sky130_fd_sc_hd__inv_1 _32792_ (.A(\inst$top.soc.cpu.sink__payload$18[186] ),
    .Y(_11875_));
 sky130_fd_sc_hd__o22ai_1 _32793_ (.A1(_11874_),
    .A2(net1192),
    .B1(_11875_),
    .B2(net1019),
    .Y(_11876_));
 sky130_fd_sc_hd__a221oi_1 _32794_ (.A1(\inst$top.soc.cpu.sink__payload$18[6] ),
    .A2(net1030),
    .B1(\inst$top.soc.cpu.sink__payload$18[115] ),
    .B2(net1069),
    .C1(_11876_),
    .Y(_11877_));
 sky130_fd_sc_hd__o21ai_0 _32796_ (.A1(\inst$top.soc.cpu.exception.w_data$51[6] ),
    .A2(net2227),
    .B1(net2043),
    .Y(_11879_));
 sky130_fd_sc_hd__a21oi_1 _32797_ (.A1(_11877_),
    .A2(net2226),
    .B1(_11879_),
    .Y(_04111_));
 sky130_fd_sc_hd__inv_2 _32798_ (.A(\inst$top.soc.cpu.sink__payload$18[39] ),
    .Y(_11880_));
 sky130_fd_sc_hd__inv_1 _32799_ (.A(\inst$top.soc.cpu.sink__payload$18[187] ),
    .Y(_11881_));
 sky130_fd_sc_hd__o22ai_1 _32800_ (.A1(_11880_),
    .A2(net1192),
    .B1(_11881_),
    .B2(net1018),
    .Y(_11882_));
 sky130_fd_sc_hd__a221oi_1 _32801_ (.A1(\inst$top.soc.cpu.sink__payload$18[7] ),
    .A2(net1027),
    .B1(\inst$top.soc.cpu.sink__payload$18[116] ),
    .B2(net1068),
    .C1(_11882_),
    .Y(_11883_));
 sky130_fd_sc_hd__o21ai_0 _32802_ (.A1(\inst$top.soc.cpu.exception.w_data$51[7] ),
    .A2(net2216),
    .B1(net2032),
    .Y(_11884_));
 sky130_fd_sc_hd__a21oi_1 _32803_ (.A1(_11883_),
    .A2(net2216),
    .B1(_11884_),
    .Y(_04112_));
 sky130_fd_sc_hd__inv_2 _32804_ (.A(\inst$top.soc.cpu.sink__payload$18[100] ),
    .Y(_11885_));
 sky130_fd_sc_hd__inv_1 _32805_ (.A(\inst$top.soc.cpu.sink__payload$18[188] ),
    .Y(_11886_));
 sky130_fd_sc_hd__o22ai_1 _32806_ (.A1(_11885_),
    .A2(net1194),
    .B1(_11886_),
    .B2(net1021),
    .Y(_11887_));
 sky130_fd_sc_hd__a221oi_1 _32807_ (.A1(\inst$top.soc.cpu.sink__payload$18[8] ),
    .A2(net1029),
    .B1(\inst$top.soc.cpu.sink__payload$18[117] ),
    .B2(net1071),
    .C1(_11887_),
    .Y(_11888_));
 sky130_fd_sc_hd__o21ai_0 _32810_ (.A1(\inst$top.soc.cpu.exception.w_data$51[8] ),
    .A2(net2239),
    .B1(net2068),
    .Y(_11891_));
 sky130_fd_sc_hd__a21oi_1 _32811_ (.A1(_11888_),
    .A2(net2239),
    .B1(_11891_),
    .Y(_04113_));
 sky130_fd_sc_hd__inv_1 _32812_ (.A(\inst$top.soc.cpu.sink__payload$18[189] ),
    .Y(_11892_));
 sky130_fd_sc_hd__o22ai_1 _32813_ (.A1(_20267_),
    .A2(net1194),
    .B1(_11892_),
    .B2(net1021),
    .Y(_11893_));
 sky130_fd_sc_hd__a221oi_1 _32814_ (.A1(\inst$top.soc.cpu.sink__payload$18[9] ),
    .A2(net1029),
    .B1(\inst$top.soc.cpu.sink__payload$18[118] ),
    .B2(net1071),
    .C1(_11893_),
    .Y(_11894_));
 sky130_fd_sc_hd__o21ai_0 _32815_ (.A1(\inst$top.soc.cpu.exception.w_data$51[9] ),
    .A2(net2228),
    .B1(net2044),
    .Y(_11895_));
 sky130_fd_sc_hd__a21oi_1 _32816_ (.A1(_11894_),
    .A2(net2228),
    .B1(_11895_),
    .Y(_04114_));
 sky130_fd_sc_hd__o21ai_0 _32819_ (.A1(\inst$top.soc.cpu.exception.w_mret ),
    .A2(net2220),
    .B1(net2084),
    .Y(_11898_));
 sky130_fd_sc_hd__a21oi_1 _32820_ (.A1(net2540),
    .A2(net2223),
    .B1(_11898_),
    .Y(_04115_));
 sky130_fd_sc_hd__o21ai_0 _32821_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mstatus.mpie.w_data ),
    .A2(net2221),
    .B1(net2084),
    .Y(_11899_));
 sky130_fd_sc_hd__a21oi_1 _32822_ (.A1(_11642_),
    .A2(net2221),
    .B1(_11899_),
    .Y(_04116_));
 sky130_fd_sc_hd__nor2_1 _32823_ (.A(\inst$top.soc.cpu.exception.m_mstatus.mpie ),
    .B(net1883),
    .Y(_11900_));
 sky130_fd_sc_hd__o21ai_0 _32824_ (.A1(\inst$top.soc.cpu.exception.w_mstatus.mpie ),
    .A2(net2220),
    .B1(net2083),
    .Y(_11901_));
 sky130_fd_sc_hd__nor2_1 _32825_ (.A(_11900_),
    .B(_11901_),
    .Y(_04117_));
 sky130_fd_sc_hd__o221ai_1 _32828_ (.A1(\inst$top.soc.cpu.exception.w_trap ),
    .A2(net2217),
    .B1(_11698_),
    .B2(_20254_),
    .C1(net2035),
    .Y(_11904_));
 sky130_fd_sc_hd__inv_2 _32829_ (.A(_11904_),
    .Y(_04118_));
 sky130_fd_sc_hd__nor2_1 _32830_ (.A(\inst$top.soc.cpu.f.source__valid ),
    .B(net666),
    .Y(_11905_));
 sky130_fd_sc_hd__inv_1 _32831_ (.A(_20360_),
    .Y(_11906_));
 sky130_fd_sc_hd__nand2_1 _32832_ (.A(_20364_),
    .B(\inst$top.soc.cpu.d.sink__payload.fence_i ),
    .Y(_11907_));
 sky130_fd_sc_hd__inv_1 _32833_ (.A(net2820),
    .Y(_11908_));
 sky130_fd_sc_hd__a21oi_1 _32834_ (.A1(_11908_),
    .A2(\inst$top.soc.cpu.sink__payload$6[45] ),
    .B1(_20296_),
    .Y(_11909_));
 sky130_fd_sc_hd__inv_1 _32835_ (.A(_11909_),
    .Y(_11910_));
 sky130_fd_sc_hd__a21oi_1 _32836_ (.A1(\inst$top.soc.cpu.sink__payload$6[63] ),
    .A2(net1191),
    .B1(_09367_),
    .Y(_11911_));
 sky130_fd_sc_hd__o21ai_1 _32837_ (.A1(_11910_),
    .A2(_11911_),
    .B1(_20348_),
    .Y(_11912_));
 sky130_fd_sc_hd__nand2_1 _32838_ (.A(net883),
    .B(_11373_),
    .Y(_11913_));
 sky130_fd_sc_hd__inv_1 _32839_ (.A(_11913_),
    .Y(_11914_));
 sky130_fd_sc_hd__nand3_1 _32840_ (.A(_11906_),
    .B(net813),
    .C(net831),
    .Y(_11915_));
 sky130_fd_sc_hd__nand4_1 _32843_ (.A(net740),
    .B(\inst$top.soc.cpu.a.source__valid ),
    .C(net813),
    .D(_20359_),
    .Y(_11918_));
 sky130_fd_sc_hd__nand2_1 _32844_ (.A(net667),
    .B(_11918_),
    .Y(_11919_));
 sky130_fd_sc_hd__nand2_1 _32845_ (.A(_11919_),
    .B(net2030),
    .Y(_11920_));
 sky130_fd_sc_hd__nor2_4 _32846_ (.A(_11905_),
    .B(_11920_),
    .Y(_04119_));
 sky130_fd_sc_hd__nand2_1 _32847_ (.A(net621),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[0] ),
    .Y(_11921_));
 sky130_fd_sc_hd__inv_1 _32848_ (.A(\inst$top.soc.cpu.sink__payload[2] ),
    .Y(_11922_));
 sky130_fd_sc_hd__nand2_1 _32849_ (.A(net740),
    .B(_11922_),
    .Y(_11923_));
 sky130_fd_sc_hd__nand3_1 _32852_ (.A(net790),
    .B(\inst$top.soc.cpu.d_branch_target[2] ),
    .C(net831),
    .Y(_11926_));
 sky130_fd_sc_hd__nand3_1 _32853_ (.A(_11923_),
    .B(_11926_),
    .C(net813),
    .Y(_11927_));
 sky130_fd_sc_hd__inv_1 _32854_ (.A(_02863_),
    .Y(_11928_));
 sky130_fd_sc_hd__o21ai_2 _32855_ (.A1(_11928_),
    .A2(_20227_),
    .B1(\inst$top.soc.cpu.x.source__valid ),
    .Y(_11929_));
 sky130_fd_sc_hd__clkinv_1 _32856_ (.A(net870),
    .Y(_11930_));
 sky130_fd_sc_hd__nor2_1 _32859_ (.A(\inst$top.soc.cpu.sink__payload$6[2] ),
    .B(net813),
    .Y(_11933_));
 sky130_fd_sc_hd__nor2_1 _32860_ (.A(net846),
    .B(_11933_),
    .Y(_11934_));
 sky130_fd_sc_hd__nand2_1 _32861_ (.A(_11927_),
    .B(_11934_),
    .Y(_11935_));
 sky130_fd_sc_hd__nand3_1 _32868_ (.A(net1816),
    .B(\inst$top.soc.cpu.sink__payload$18[182] ),
    .C(net1838),
    .Y(_11942_));
 sky130_fd_sc_hd__o211ai_1 _32869_ (.A1(_20462_),
    .A2(net1816),
    .B1(net2537),
    .C1(_11942_),
    .Y(_11943_));
 sky130_fd_sc_hd__o211ai_1 _32871_ (.A1(net2537),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[0] ),
    .B1(_11943_),
    .C1(net872),
    .Y(_11945_));
 sky130_fd_sc_hd__o21ai_0 _32872_ (.A1(_20472_),
    .A2(net872),
    .B1(_11945_),
    .Y(_11946_));
 sky130_fd_sc_hd__nand2_1 _32874_ (.A(_11946_),
    .B(net846),
    .Y(_11948_));
 sky130_fd_sc_hd__nand2_1 _32875_ (.A(_11935_),
    .B(_11948_),
    .Y(_11949_));
 sky130_fd_sc_hd__nand3_1 _32878_ (.A(_11949_),
    .B(net663),
    .C(net753),
    .Y(_11952_));
 sky130_fd_sc_hd__a21oi_4 _32879_ (.A1(_11921_),
    .A2(_11952_),
    .B1(net2935),
    .Y(_04120_));
 sky130_fd_sc_hd__nand2_1 _32880_ (.A(net626),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[10] ),
    .Y(_11953_));
 sky130_fd_sc_hd__inv_1 _32883_ (.A(\inst$top.soc.cpu.sink__payload[10] ),
    .Y(_11956_));
 sky130_fd_sc_hd__inv_1 _32884_ (.A(\inst$top.soc.cpu.sink__payload[11] ),
    .Y(_11957_));
 sky130_fd_sc_hd__nand2_1 _32885_ (.A(\inst$top.soc.cpu.sink__payload[6] ),
    .B(\inst$top.soc.cpu.sink__payload[7] ),
    .Y(_11958_));
 sky130_fd_sc_hd__nand3_1 _32886_ (.A(_02866_),
    .B(\inst$top.soc.cpu.sink__payload[4] ),
    .C(\inst$top.soc.cpu.sink__payload[5] ),
    .Y(_11959_));
 sky130_fd_sc_hd__nor2_1 _32887_ (.A(_11958_),
    .B(_11959_),
    .Y(_11960_));
 sky130_fd_sc_hd__nand3_1 _32888_ (.A(_11960_),
    .B(\inst$top.soc.cpu.sink__payload[8] ),
    .C(\inst$top.soc.cpu.sink__payload[9] ),
    .Y(_11961_));
 sky130_fd_sc_hd__nor3_1 _32889_ (.A(_11956_),
    .B(_11957_),
    .C(_11961_),
    .Y(_11962_));
 sky130_fd_sc_hd__xor2_1 _32890_ (.A(\inst$top.soc.cpu.sink__payload[12] ),
    .B(_11962_),
    .X(_11963_));
 sky130_fd_sc_hd__nand3_1 _32891_ (.A(net741),
    .B(net815),
    .C(_11963_),
    .Y(_11964_));
 sky130_fd_sc_hd__a21oi_1 _32893_ (.A1(net837),
    .A2(\inst$top.soc.cpu.sink__payload$6[12] ),
    .B1(net849),
    .Y(_11966_));
 sky130_fd_sc_hd__nand2_1 _32895_ (.A(_03322_),
    .B(_03319_),
    .Y(_11968_));
 sky130_fd_sc_hd__inv_1 _32896_ (.A(_03321_),
    .Y(_11969_));
 sky130_fd_sc_hd__nand2_1 _32897_ (.A(_11968_),
    .B(_11969_),
    .Y(_11970_));
 sky130_fd_sc_hd__nand2_1 _32898_ (.A(_03320_),
    .B(_03322_),
    .Y(_11971_));
 sky130_fd_sc_hd__a21oi_1 _32899_ (.A1(_03318_),
    .A2(_03315_),
    .B1(_03317_),
    .Y(_11972_));
 sky130_fd_sc_hd__nor2_1 _32900_ (.A(_11971_),
    .B(_11972_),
    .Y(_11973_));
 sky130_fd_sc_hd__nor2_1 _32901_ (.A(_11970_),
    .B(_11973_),
    .Y(_11974_));
 sky130_fd_sc_hd__a21oi_1 _32902_ (.A1(_03314_),
    .A2(_03311_),
    .B1(_03313_),
    .Y(_11975_));
 sky130_fd_sc_hd__nand3_1 _32903_ (.A(_02546_),
    .B(_03312_),
    .C(_03314_),
    .Y(_11976_));
 sky130_fd_sc_hd__nand2_1 _32904_ (.A(_11975_),
    .B(_11976_),
    .Y(_11977_));
 sky130_fd_sc_hd__nand2_1 _32905_ (.A(_03316_),
    .B(_03318_),
    .Y(_11978_));
 sky130_fd_sc_hd__nor2_1 _32906_ (.A(_11978_),
    .B(_11971_),
    .Y(_11979_));
 sky130_fd_sc_hd__nand2_1 _32907_ (.A(_11977_),
    .B(_11979_),
    .Y(_11980_));
 sky130_fd_sc_hd__nand2_1 _32908_ (.A(_11974_),
    .B(_11980_),
    .Y(_11981_));
 sky130_fd_sc_hd__nand2_1 _32909_ (.A(_03324_),
    .B(_03326_),
    .Y(_11982_));
 sky130_fd_sc_hd__inv_1 _32910_ (.A(_11982_),
    .Y(_11983_));
 sky130_fd_sc_hd__nand2_1 _32911_ (.A(_11981_),
    .B(_11983_),
    .Y(_11984_));
 sky130_fd_sc_hd__a21oi_1 _32912_ (.A1(_03326_),
    .A2(_03323_),
    .B1(_03325_),
    .Y(_11985_));
 sky130_fd_sc_hd__nand2_1 _32913_ (.A(_11984_),
    .B(_11985_),
    .Y(_11986_));
 sky130_fd_sc_hd__xor2_1 _32914_ (.A(_03328_),
    .B(_11986_),
    .X(_11987_));
 sky130_fd_sc_hd__nand3_1 _32915_ (.A(net791),
    .B(net832),
    .C(_11987_),
    .Y(_11988_));
 sky130_fd_sc_hd__nand3_1 _32916_ (.A(_11964_),
    .B(_11966_),
    .C(_11988_),
    .Y(_11989_));
 sky130_fd_sc_hd__nand3_1 _32920_ (.A(net1817),
    .B(\inst$top.soc.cpu.sink__payload$18[192] ),
    .C(net1840),
    .Y(_11993_));
 sky130_fd_sc_hd__o211ai_1 _32921_ (.A1(_20751_),
    .A2(net1817),
    .B1(net2545),
    .C1(_11993_),
    .Y(_11994_));
 sky130_fd_sc_hd__o211ai_1 _32923_ (.A1(net2538),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[10] ),
    .B1(_11994_),
    .C1(net873),
    .Y(_11996_));
 sky130_fd_sc_hd__o211ai_1 _32925_ (.A1(_20760_),
    .A2(net873),
    .B1(_11996_),
    .C1(net848),
    .Y(_11998_));
 sky130_fd_sc_hd__nand2_1 _32926_ (.A(_11989_),
    .B(_11998_),
    .Y(_11999_));
 sky130_fd_sc_hd__inv_1 _32927_ (.A(_11999_),
    .Y(_12000_));
 sky130_fd_sc_hd__nand3_1 _32928_ (.A(_12000_),
    .B(net664),
    .C(net754),
    .Y(_12001_));
 sky130_fd_sc_hd__a21oi_4 _32929_ (.A1(_11953_),
    .A2(_12001_),
    .B1(net2932),
    .Y(_04121_));
 sky130_fd_sc_hd__nand2_1 _32930_ (.A(net628),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[11] ),
    .Y(_12002_));
 sky130_fd_sc_hd__inv_1 _32931_ (.A(\inst$top.soc.cpu.sink__payload[12] ),
    .Y(_12003_));
 sky130_fd_sc_hd__nand2_1 _32932_ (.A(\inst$top.soc.cpu.sink__payload[9] ),
    .B(\inst$top.soc.cpu.sink__payload[10] ),
    .Y(_12004_));
 sky130_fd_sc_hd__nand3_1 _32933_ (.A(\inst$top.soc.cpu.sink__payload[2] ),
    .B(\inst$top.soc.cpu.sink__payload[4] ),
    .C(\inst$top.soc.cpu.sink__payload[3] ),
    .Y(_12005_));
 sky130_fd_sc_hd__inv_1 _32934_ (.A(_12005_),
    .Y(_12006_));
 sky130_fd_sc_hd__nand3_1 _32935_ (.A(_12006_),
    .B(\inst$top.soc.cpu.sink__payload[5] ),
    .C(\inst$top.soc.cpu.sink__payload[6] ),
    .Y(_12007_));
 sky130_fd_sc_hd__nand3b_1 _32936_ (.A_N(_12007_),
    .B(\inst$top.soc.cpu.sink__payload[7] ),
    .C(\inst$top.soc.cpu.sink__payload[8] ),
    .Y(_12008_));
 sky130_fd_sc_hd__nor4_1 _32937_ (.A(_11957_),
    .B(_12003_),
    .C(_12004_),
    .D(_12008_),
    .Y(_12009_));
 sky130_fd_sc_hd__xor2_1 _32938_ (.A(\inst$top.soc.cpu.sink__payload[13] ),
    .B(_12009_),
    .X(_12010_));
 sky130_fd_sc_hd__nand2_1 _32939_ (.A(net742),
    .B(_12010_),
    .Y(_12011_));
 sky130_fd_sc_hd__nand3_1 _32940_ (.A(_02911_),
    .B(_02545_),
    .C(_03312_),
    .Y(_12012_));
 sky130_fd_sc_hd__inv_1 _32941_ (.A(_03311_),
    .Y(_12013_));
 sky130_fd_sc_hd__nand2_1 _32942_ (.A(_03312_),
    .B(_03310_),
    .Y(_12014_));
 sky130_fd_sc_hd__nand3_1 _32943_ (.A(_12012_),
    .B(_12013_),
    .C(_12014_),
    .Y(_12015_));
 sky130_fd_sc_hd__nand2_1 _32944_ (.A(_03314_),
    .B(_03316_),
    .Y(_12016_));
 sky130_fd_sc_hd__inv_1 _32945_ (.A(_12016_),
    .Y(_12017_));
 sky130_fd_sc_hd__nand2_1 _32946_ (.A(_03318_),
    .B(_03320_),
    .Y(_12018_));
 sky130_fd_sc_hd__inv_1 _32947_ (.A(_12018_),
    .Y(_12019_));
 sky130_fd_sc_hd__nand3_1 _32948_ (.A(_12015_),
    .B(_12017_),
    .C(_12019_),
    .Y(_12020_));
 sky130_fd_sc_hd__a21o_1 _32949_ (.A1(_03316_),
    .A2(_03313_),
    .B1(_03315_),
    .X(_12021_));
 sky130_fd_sc_hd__nand2_1 _32950_ (.A(_12021_),
    .B(_12019_),
    .Y(_12022_));
 sky130_fd_sc_hd__a21oi_1 _32951_ (.A1(_03320_),
    .A2(_03317_),
    .B1(_03319_),
    .Y(_12023_));
 sky130_fd_sc_hd__nand3_1 _32952_ (.A(_12020_),
    .B(_12022_),
    .C(_12023_),
    .Y(_12024_));
 sky130_fd_sc_hd__nand2_1 _32953_ (.A(_12024_),
    .B(_03322_),
    .Y(_12025_));
 sky130_fd_sc_hd__nand2_1 _32954_ (.A(_12025_),
    .B(_11969_),
    .Y(_12026_));
 sky130_fd_sc_hd__a21o_1 _32955_ (.A1(_12026_),
    .A2(_03324_),
    .B1(_03323_),
    .X(_12027_));
 sky130_fd_sc_hd__nand3_1 _32956_ (.A(_12027_),
    .B(_03326_),
    .C(_03328_),
    .Y(_12028_));
 sky130_fd_sc_hd__a21oi_1 _32957_ (.A1(_03328_),
    .A2(_03325_),
    .B1(_03327_),
    .Y(_12029_));
 sky130_fd_sc_hd__nand2_1 _32958_ (.A(_12028_),
    .B(_12029_),
    .Y(_12030_));
 sky130_fd_sc_hd__xor2_1 _32959_ (.A(_03330_),
    .B(_12030_),
    .X(_12031_));
 sky130_fd_sc_hd__nand3_1 _32960_ (.A(net792),
    .B(net833),
    .C(_12031_),
    .Y(_12032_));
 sky130_fd_sc_hd__nand3_1 _32961_ (.A(_12011_),
    .B(_12032_),
    .C(net816),
    .Y(_12033_));
 sky130_fd_sc_hd__nor2_1 _32962_ (.A(\inst$top.soc.cpu.sink__payload$6[13] ),
    .B(net816),
    .Y(_12034_));
 sky130_fd_sc_hd__nor2_1 _32963_ (.A(net849),
    .B(_12034_),
    .Y(_12035_));
 sky130_fd_sc_hd__nand2_1 _32964_ (.A(_12033_),
    .B(_12035_),
    .Y(_12036_));
 sky130_fd_sc_hd__nand3_1 _32965_ (.A(net1820),
    .B(\inst$top.soc.cpu.sink__payload$18[193] ),
    .C(net1839),
    .Y(_12037_));
 sky130_fd_sc_hd__o211ai_1 _32966_ (.A1(_20771_),
    .A2(net1818),
    .B1(net2543),
    .C1(_12037_),
    .Y(_12038_));
 sky130_fd_sc_hd__o211ai_1 _32967_ (.A1(net2541),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[11] ),
    .B1(_12038_),
    .C1(net876),
    .Y(_12039_));
 sky130_fd_sc_hd__o21ai_0 _32968_ (.A1(_20778_),
    .A2(net876),
    .B1(_12039_),
    .Y(_12040_));
 sky130_fd_sc_hd__nand2_1 _32969_ (.A(_12040_),
    .B(net849),
    .Y(_12041_));
 sky130_fd_sc_hd__nand2_1 _32970_ (.A(_12036_),
    .B(_12041_),
    .Y(_12042_));
 sky130_fd_sc_hd__nand3_1 _32971_ (.A(_12042_),
    .B(net664),
    .C(net754),
    .Y(_12043_));
 sky130_fd_sc_hd__a21oi_4 _32972_ (.A1(_12002_),
    .A2(_12043_),
    .B1(net2944),
    .Y(_04122_));
 sky130_fd_sc_hd__nand2_1 _32973_ (.A(net627),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[12] ),
    .Y(_12044_));
 sky130_fd_sc_hd__inv_1 _32974_ (.A(\inst$top.soc.cpu.sink__payload[14] ),
    .Y(_12045_));
 sky130_fd_sc_hd__nand3_1 _32975_ (.A(_11962_),
    .B(\inst$top.soc.cpu.sink__payload[12] ),
    .C(\inst$top.soc.cpu.sink__payload[13] ),
    .Y(_12046_));
 sky130_fd_sc_hd__xor2_1 _32976_ (.A(_12045_),
    .B(_12046_),
    .X(_12047_));
 sky130_fd_sc_hd__nand3_1 _32977_ (.A(net742),
    .B(net816),
    .C(_12047_),
    .Y(_12048_));
 sky130_fd_sc_hd__nand2_1 _32978_ (.A(_03328_),
    .B(_03330_),
    .Y(_12049_));
 sky130_fd_sc_hd__inv_1 _32979_ (.A(_12049_),
    .Y(_12050_));
 sky130_fd_sc_hd__a21oi_1 _32980_ (.A1(_03330_),
    .A2(_03327_),
    .B1(_03329_),
    .Y(_12051_));
 sky130_fd_sc_hd__o21ai_0 _32981_ (.A1(_12049_),
    .A2(_11985_),
    .B1(_12051_),
    .Y(_12052_));
 sky130_fd_sc_hd__a31oi_1 _32982_ (.A1(_11981_),
    .A2(_11983_),
    .A3(_12050_),
    .B1(_12052_),
    .Y(_12053_));
 sky130_fd_sc_hd__xnor2_1 _32983_ (.A(_03332_),
    .B(_12053_),
    .Y(_12054_));
 sky130_fd_sc_hd__nand3_1 _32984_ (.A(net792),
    .B(net833),
    .C(_12054_),
    .Y(_12055_));
 sky130_fd_sc_hd__a21oi_1 _32985_ (.A1(net838),
    .A2(\inst$top.soc.cpu.sink__payload$6[14] ),
    .B1(net849),
    .Y(_12056_));
 sky130_fd_sc_hd__nand3_1 _32986_ (.A(_12048_),
    .B(_12055_),
    .C(_12056_),
    .Y(_12057_));
 sky130_fd_sc_hd__nand3_1 _32987_ (.A(net1817),
    .B(\inst$top.soc.cpu.sink__payload$18[194] ),
    .C(net1840),
    .Y(_12058_));
 sky130_fd_sc_hd__o211ai_1 _32988_ (.A1(_20789_),
    .A2(net1817),
    .B1(net2541),
    .C1(_12058_),
    .Y(_12059_));
 sky130_fd_sc_hd__o211ai_1 _32989_ (.A1(net2541),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[12] ),
    .B1(_12059_),
    .C1(net879),
    .Y(_12060_));
 sky130_fd_sc_hd__o211ai_1 _32990_ (.A1(_20796_),
    .A2(net876),
    .B1(_12060_),
    .C1(net851),
    .Y(_12061_));
 sky130_fd_sc_hd__nand2_1 _32991_ (.A(_12057_),
    .B(_12061_),
    .Y(_12062_));
 sky130_fd_sc_hd__inv_1 _32992_ (.A(_12062_),
    .Y(_12063_));
 sky130_fd_sc_hd__nand3_1 _32993_ (.A(_12063_),
    .B(net664),
    .C(net754),
    .Y(_12064_));
 sky130_fd_sc_hd__a21oi_4 _32994_ (.A1(_12044_),
    .A2(_12064_),
    .B1(net2944),
    .Y(_04123_));
 sky130_fd_sc_hd__nand2_1 _32995_ (.A(net628),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[13] ),
    .Y(_12065_));
 sky130_fd_sc_hd__inv_1 _32996_ (.A(\inst$top.soc.cpu.sink__payload[15] ),
    .Y(_12066_));
 sky130_fd_sc_hd__nor2_1 _32997_ (.A(_12004_),
    .B(_12008_),
    .Y(_12067_));
 sky130_fd_sc_hd__inv_1 _32998_ (.A(\inst$top.soc.cpu.sink__payload[13] ),
    .Y(_12068_));
 sky130_fd_sc_hd__nor4_1 _32999_ (.A(_11957_),
    .B(_12003_),
    .C(_12068_),
    .D(_12045_),
    .Y(_12069_));
 sky130_fd_sc_hd__nand2_1 _33000_ (.A(_12067_),
    .B(_12069_),
    .Y(_12070_));
 sky130_fd_sc_hd__xor2_1 _33001_ (.A(_12066_),
    .B(_12070_),
    .X(_12071_));
 sky130_fd_sc_hd__nand3_1 _33002_ (.A(net742),
    .B(net816),
    .C(_12071_),
    .Y(_12072_));
 sky130_fd_sc_hd__a21oi_1 _33003_ (.A1(net838),
    .A2(\inst$top.soc.cpu.sink__payload$6[15] ),
    .B1(net849),
    .Y(_12073_));
 sky130_fd_sc_hd__nand2_1 _33004_ (.A(_03322_),
    .B(_03324_),
    .Y(_12074_));
 sky130_fd_sc_hd__a21oi_1 _33005_ (.A1(_03324_),
    .A2(_03321_),
    .B1(_03323_),
    .Y(_12075_));
 sky130_fd_sc_hd__o21ai_0 _33006_ (.A1(_12074_),
    .A2(_12023_),
    .B1(_12075_),
    .Y(_12076_));
 sky130_fd_sc_hd__nand2_1 _33007_ (.A(_03326_),
    .B(_03328_),
    .Y(_12077_));
 sky130_fd_sc_hd__nand2_1 _33008_ (.A(_03330_),
    .B(_03332_),
    .Y(_12078_));
 sky130_fd_sc_hd__nor2_1 _33009_ (.A(_12077_),
    .B(_12078_),
    .Y(_12079_));
 sky130_fd_sc_hd__a21oi_1 _33010_ (.A1(_03332_),
    .A2(_03329_),
    .B1(_03331_),
    .Y(_12080_));
 sky130_fd_sc_hd__o21ai_0 _33011_ (.A1(_12078_),
    .A2(_12029_),
    .B1(_12080_),
    .Y(_12081_));
 sky130_fd_sc_hd__a21oi_1 _33012_ (.A1(_12076_),
    .A2(_12079_),
    .B1(_12081_),
    .Y(_12082_));
 sky130_fd_sc_hd__a21oi_1 _33013_ (.A1(_12014_),
    .A2(_12013_),
    .B1(_12016_),
    .Y(_12083_));
 sky130_fd_sc_hd__nor2_1 _33014_ (.A(_12021_),
    .B(_12083_),
    .Y(_12084_));
 sky130_fd_sc_hd__nand4_1 _33015_ (.A(_12017_),
    .B(_02911_),
    .C(_02545_),
    .D(_03312_),
    .Y(_12085_));
 sky130_fd_sc_hd__nand2_1 _33016_ (.A(_12084_),
    .B(_12085_),
    .Y(_12086_));
 sky130_fd_sc_hd__nor2_1 _33017_ (.A(_12018_),
    .B(_12074_),
    .Y(_12087_));
 sky130_fd_sc_hd__nand3_1 _33018_ (.A(_12086_),
    .B(_12087_),
    .C(_12079_),
    .Y(_12088_));
 sky130_fd_sc_hd__nand2_1 _33019_ (.A(_12082_),
    .B(_12088_),
    .Y(_12089_));
 sky130_fd_sc_hd__xor2_1 _33020_ (.A(_03334_),
    .B(_12089_),
    .X(_12090_));
 sky130_fd_sc_hd__nand3_1 _33021_ (.A(net792),
    .B(net833),
    .C(_12090_),
    .Y(_12091_));
 sky130_fd_sc_hd__nand3_1 _33022_ (.A(_12072_),
    .B(_12073_),
    .C(_12091_),
    .Y(_12092_));
 sky130_fd_sc_hd__nand3_1 _33024_ (.A(net1820),
    .B(\inst$top.soc.cpu.sink__payload$18[195] ),
    .C(net1839),
    .Y(_12094_));
 sky130_fd_sc_hd__o211ai_1 _33025_ (.A1(_20807_),
    .A2(net1820),
    .B1(net2544),
    .C1(_12094_),
    .Y(_12095_));
 sky130_fd_sc_hd__o211ai_1 _33026_ (.A1(net2544),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[13] ),
    .B1(_12095_),
    .C1(net879),
    .Y(_12096_));
 sky130_fd_sc_hd__o211ai_1 _33027_ (.A1(_20817_),
    .A2(net879),
    .B1(_12096_),
    .C1(net851),
    .Y(_12097_));
 sky130_fd_sc_hd__nand2_1 _33028_ (.A(_12092_),
    .B(_12097_),
    .Y(_12098_));
 sky130_fd_sc_hd__inv_1 _33029_ (.A(_12098_),
    .Y(_12099_));
 sky130_fd_sc_hd__nand3_1 _33030_ (.A(_12099_),
    .B(net664),
    .C(net754),
    .Y(_12100_));
 sky130_fd_sc_hd__a21oi_4 _33031_ (.A1(_12065_),
    .A2(_12100_),
    .B1(net2944),
    .Y(_04124_));
 sky130_fd_sc_hd__nor4_1 _33033_ (.A(_12003_),
    .B(_12068_),
    .C(_12045_),
    .D(_12066_),
    .Y(_12102_));
 sky130_fd_sc_hd__nand2_1 _33034_ (.A(_11962_),
    .B(_12102_),
    .Y(_12103_));
 sky130_fd_sc_hd__inv_1 _33035_ (.A(_12103_),
    .Y(_12104_));
 sky130_fd_sc_hd__nor2_1 _33036_ (.A(\inst$top.soc.cpu.sink__payload[16] ),
    .B(_12104_),
    .Y(_12105_));
 sky130_fd_sc_hd__inv_1 _33037_ (.A(\inst$top.soc.cpu.sink__payload[16] ),
    .Y(_12106_));
 sky130_fd_sc_hd__nor2_1 _33038_ (.A(_12106_),
    .B(_12103_),
    .Y(_12107_));
 sky130_fd_sc_hd__o21ai_0 _33039_ (.A1(_12105_),
    .A2(_12107_),
    .B1(net742),
    .Y(_12108_));
 sky130_fd_sc_hd__nand2_1 _33040_ (.A(_03332_),
    .B(_03334_),
    .Y(_12109_));
 sky130_fd_sc_hd__a21oi_1 _33041_ (.A1(_03334_),
    .A2(_03331_),
    .B1(_03333_),
    .Y(_12110_));
 sky130_fd_sc_hd__o21ai_0 _33042_ (.A1(_12109_),
    .A2(_12051_),
    .B1(_12110_),
    .Y(_12111_));
 sky130_fd_sc_hd__a41oi_1 _33043_ (.A1(_11986_),
    .A2(_03332_),
    .A3(_03334_),
    .A4(_12050_),
    .B1(_12111_),
    .Y(_12112_));
 sky130_fd_sc_hd__xor2_1 _33044_ (.A(_03336_),
    .B(_12112_),
    .X(_12113_));
 sky130_fd_sc_hd__nand3_1 _33045_ (.A(net791),
    .B(net832),
    .C(_12113_),
    .Y(_12114_));
 sky130_fd_sc_hd__nand3_1 _33046_ (.A(_12108_),
    .B(_12114_),
    .C(net815),
    .Y(_12115_));
 sky130_fd_sc_hd__a21oi_1 _33048_ (.A1(net838),
    .A2(\inst$top.soc.cpu.sink__payload$6[16] ),
    .B1(net849),
    .Y(_12117_));
 sky130_fd_sc_hd__nand3_1 _33051_ (.A(net1821),
    .B(\inst$top.soc.cpu.sink__payload$18[196] ),
    .C(net1840),
    .Y(_12120_));
 sky130_fd_sc_hd__o211ai_1 _33052_ (.A1(_05598_),
    .A2(net1821),
    .B1(net2541),
    .C1(_12120_),
    .Y(_12121_));
 sky130_fd_sc_hd__o211ai_1 _33053_ (.A1(net2545),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[14] ),
    .B1(_12121_),
    .C1(net880),
    .Y(_12122_));
 sky130_fd_sc_hd__o21ai_0 _33054_ (.A1(_05605_),
    .A2(net880),
    .B1(_12122_),
    .Y(_12123_));
 sky130_fd_sc_hd__nor2_1 _33055_ (.A(net870),
    .B(_12123_),
    .Y(_12124_));
 sky130_fd_sc_hd__a21oi_1 _33056_ (.A1(_12115_),
    .A2(_12117_),
    .B1(_12124_),
    .Y(_12125_));
 sky130_fd_sc_hd__nand2_1 _33057_ (.A(net676),
    .B(_12125_),
    .Y(_12126_));
 sky130_fd_sc_hd__nand2_1 _33059_ (.A(net627),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[14] ),
    .Y(_12128_));
 sky130_fd_sc_hd__a21oi_4 _33060_ (.A1(_12126_),
    .A2(_12128_),
    .B1(net2932),
    .Y(_04125_));
 sky130_fd_sc_hd__nand2_1 _33061_ (.A(net628),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[15] ),
    .Y(_12129_));
 sky130_fd_sc_hd__inv_1 _33062_ (.A(\inst$top.soc.cpu.sink__payload[17] ),
    .Y(_12130_));
 sky130_fd_sc_hd__nor4_1 _33063_ (.A(_12068_),
    .B(_12045_),
    .C(_12066_),
    .D(_12106_),
    .Y(_12131_));
 sky130_fd_sc_hd__nand2_1 _33064_ (.A(_12009_),
    .B(_12131_),
    .Y(_12132_));
 sky130_fd_sc_hd__xor2_1 _33065_ (.A(_12130_),
    .B(_12132_),
    .X(_12133_));
 sky130_fd_sc_hd__nand2_1 _33066_ (.A(net742),
    .B(_12133_),
    .Y(_12134_));
 sky130_fd_sc_hd__nand4_1 _33067_ (.A(_03330_),
    .B(_03332_),
    .C(_03334_),
    .D(_03336_),
    .Y(_12135_));
 sky130_fd_sc_hd__nor3_1 _33068_ (.A(_12074_),
    .B(_12077_),
    .C(_12135_),
    .Y(_12136_));
 sky130_fd_sc_hd__o21a_1 _33069_ (.A1(_12077_),
    .A2(_12075_),
    .B1(_12029_),
    .X(_12137_));
 sky130_fd_sc_hd__nand2_1 _33070_ (.A(_03334_),
    .B(_03336_),
    .Y(_12138_));
 sky130_fd_sc_hd__a21oi_1 _33071_ (.A1(_03336_),
    .A2(_03333_),
    .B1(_03335_),
    .Y(_12139_));
 sky130_fd_sc_hd__o21ai_0 _33072_ (.A1(_12138_),
    .A2(_12080_),
    .B1(_12139_),
    .Y(_12140_));
 sky130_fd_sc_hd__o21bai_1 _33073_ (.A1(_12135_),
    .A2(_12137_),
    .B1_N(_12140_),
    .Y(_12141_));
 sky130_fd_sc_hd__a21oi_1 _33074_ (.A1(_12024_),
    .A2(_12136_),
    .B1(_12141_),
    .Y(_12142_));
 sky130_fd_sc_hd__xor2_1 _33075_ (.A(_03338_),
    .B(_12142_),
    .X(_12143_));
 sky130_fd_sc_hd__inv_1 _33076_ (.A(_12143_),
    .Y(_12144_));
 sky130_fd_sc_hd__nand3_1 _33077_ (.A(net791),
    .B(net832),
    .C(_12144_),
    .Y(_12145_));
 sky130_fd_sc_hd__nand3_1 _33078_ (.A(_12134_),
    .B(_12145_),
    .C(net815),
    .Y(_12146_));
 sky130_fd_sc_hd__nor2_1 _33079_ (.A(\inst$top.soc.cpu.sink__payload$6[17] ),
    .B(net816),
    .Y(_12147_));
 sky130_fd_sc_hd__nor2_1 _33080_ (.A(net849),
    .B(_12147_),
    .Y(_12148_));
 sky130_fd_sc_hd__nand2_1 _33081_ (.A(_12146_),
    .B(_12148_),
    .Y(_12149_));
 sky130_fd_sc_hd__nand3_1 _33082_ (.A(net1817),
    .B(\inst$top.soc.cpu.sink__payload$18[197] ),
    .C(net1840),
    .Y(_12150_));
 sky130_fd_sc_hd__o211ai_1 _33083_ (.A1(_05622_),
    .A2(net1817),
    .B1(net2541),
    .C1(_12150_),
    .Y(_12151_));
 sky130_fd_sc_hd__o211ai_1 _33084_ (.A1(net2541),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[15] ),
    .B1(_12151_),
    .C1(net876),
    .Y(_12152_));
 sky130_fd_sc_hd__o21ai_0 _33085_ (.A1(_11525_),
    .A2(net876),
    .B1(_12152_),
    .Y(_12153_));
 sky130_fd_sc_hd__nand2_1 _33086_ (.A(_12153_),
    .B(net849),
    .Y(_12154_));
 sky130_fd_sc_hd__nand2_1 _33087_ (.A(_12149_),
    .B(_12154_),
    .Y(_12155_));
 sky130_fd_sc_hd__nand3_1 _33088_ (.A(_12155_),
    .B(net663),
    .C(net753),
    .Y(_12156_));
 sky130_fd_sc_hd__a21oi_4 _33089_ (.A1(_12129_),
    .A2(_12156_),
    .B1(net2932),
    .Y(_04126_));
 sky130_fd_sc_hd__nand2_1 _33091_ (.A(net626),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[16] ),
    .Y(_12158_));
 sky130_fd_sc_hd__nor4_1 _33093_ (.A(_12045_),
    .B(_12066_),
    .C(_12106_),
    .D(_12130_),
    .Y(_12160_));
 sky130_fd_sc_hd__inv_1 _33094_ (.A(_12160_),
    .Y(_12161_));
 sky130_fd_sc_hd__nor2_1 _33095_ (.A(_12161_),
    .B(_12046_),
    .Y(_12162_));
 sky130_fd_sc_hd__xor2_1 _33096_ (.A(\inst$top.soc.cpu.sink__payload[18] ),
    .B(_12162_),
    .X(_12163_));
 sky130_fd_sc_hd__nand3_1 _33097_ (.A(net741),
    .B(net814),
    .C(_12163_),
    .Y(_12164_));
 sky130_fd_sc_hd__nand2_1 _33098_ (.A(_03336_),
    .B(_03338_),
    .Y(_12165_));
 sky130_fd_sc_hd__a21oi_1 _33099_ (.A1(_03338_),
    .A2(_03335_),
    .B1(_03337_),
    .Y(_12166_));
 sky130_fd_sc_hd__o21ai_0 _33100_ (.A1(_12165_),
    .A2(_12112_),
    .B1(_12166_),
    .Y(_12167_));
 sky130_fd_sc_hd__xor2_1 _33101_ (.A(_03340_),
    .B(_12167_),
    .X(_12168_));
 sky130_fd_sc_hd__nand3_1 _33102_ (.A(net790),
    .B(net831),
    .C(_12168_),
    .Y(_12169_));
 sky130_fd_sc_hd__a21oi_1 _33103_ (.A1(net837),
    .A2(\inst$top.soc.cpu.sink__payload$6[18] ),
    .B1(net846),
    .Y(_12170_));
 sky130_fd_sc_hd__nand3_1 _33104_ (.A(_12164_),
    .B(_12169_),
    .C(_12170_),
    .Y(_12171_));
 sky130_fd_sc_hd__nand3_1 _33105_ (.A(net1815),
    .B(\inst$top.soc.cpu.sink__payload$18[198] ),
    .C(net1838),
    .Y(_12172_));
 sky130_fd_sc_hd__o211ai_1 _33106_ (.A1(_05644_),
    .A2(net1815),
    .B1(net2538),
    .C1(_12172_),
    .Y(_12173_));
 sky130_fd_sc_hd__o211ai_1 _33107_ (.A1(net2539),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[16] ),
    .B1(_12173_),
    .C1(net873),
    .Y(_12174_));
 sky130_fd_sc_hd__o211ai_1 _33108_ (.A1(_11527_),
    .A2(net873),
    .B1(_12174_),
    .C1(net848),
    .Y(_12175_));
 sky130_fd_sc_hd__nand2_1 _33109_ (.A(_12171_),
    .B(_12175_),
    .Y(_12176_));
 sky130_fd_sc_hd__inv_1 _33110_ (.A(_12176_),
    .Y(_12177_));
 sky130_fd_sc_hd__nand3_1 _33111_ (.A(_12177_),
    .B(net663),
    .C(net753),
    .Y(_12178_));
 sky130_fd_sc_hd__a21oi_4 _33113_ (.A1(_12158_),
    .A2(_12178_),
    .B1(net2934),
    .Y(_04127_));
 sky130_fd_sc_hd__inv_1 _33114_ (.A(\inst$top.soc.cpu.sink__payload[18] ),
    .Y(_12180_));
 sky130_fd_sc_hd__nor4_1 _33115_ (.A(_12066_),
    .B(_12106_),
    .C(_12130_),
    .D(_12180_),
    .Y(_12181_));
 sky130_fd_sc_hd__nand3_1 _33116_ (.A(_12067_),
    .B(_12069_),
    .C(_12181_),
    .Y(_12182_));
 sky130_fd_sc_hd__inv_1 _33117_ (.A(_12182_),
    .Y(_12183_));
 sky130_fd_sc_hd__nand2_1 _33118_ (.A(_12183_),
    .B(\inst$top.soc.cpu.sink__payload[19] ),
    .Y(_12184_));
 sky130_fd_sc_hd__inv_1 _33119_ (.A(\inst$top.soc.cpu.sink__payload[19] ),
    .Y(_12185_));
 sky130_fd_sc_hd__nand2_1 _33120_ (.A(_12182_),
    .B(_12185_),
    .Y(_12186_));
 sky130_fd_sc_hd__nand2_1 _33121_ (.A(_12184_),
    .B(_12186_),
    .Y(_12187_));
 sky130_fd_sc_hd__nand2_1 _33122_ (.A(net741),
    .B(_12187_),
    .Y(_12188_));
 sky130_fd_sc_hd__nand2_1 _33125_ (.A(_03338_),
    .B(_03340_),
    .Y(_12191_));
 sky130_fd_sc_hd__a21oi_1 _33126_ (.A1(_03340_),
    .A2(_03337_),
    .B1(_03339_),
    .Y(_12192_));
 sky130_fd_sc_hd__o21ai_0 _33127_ (.A1(_12191_),
    .A2(_12142_),
    .B1(_12192_),
    .Y(_12193_));
 sky130_fd_sc_hd__xnor2_1 _33128_ (.A(_03342_),
    .B(_12193_),
    .Y(_12194_));
 sky130_fd_sc_hd__nand3_1 _33129_ (.A(net791),
    .B(net832),
    .C(_12194_),
    .Y(_12195_));
 sky130_fd_sc_hd__nand3_1 _33131_ (.A(_12188_),
    .B(_12195_),
    .C(net814),
    .Y(_12197_));
 sky130_fd_sc_hd__nand2_1 _33132_ (.A(net837),
    .B(\inst$top.soc.cpu.sink__payload$6[19] ),
    .Y(_12198_));
 sky130_fd_sc_hd__nand2_1 _33133_ (.A(_12197_),
    .B(_12198_),
    .Y(_12199_));
 sky130_fd_sc_hd__nand2_1 _33135_ (.A(_12199_),
    .B(net870),
    .Y(_12201_));
 sky130_fd_sc_hd__nand3_1 _33139_ (.A(net1815),
    .B(\inst$top.soc.cpu.sink__payload$18[199] ),
    .C(_02865_),
    .Y(_12205_));
 sky130_fd_sc_hd__o211ai_1 _33140_ (.A1(_05666_),
    .A2(net1821),
    .B1(net2538),
    .C1(_12205_),
    .Y(_12206_));
 sky130_fd_sc_hd__o211ai_1 _33142_ (.A1(net2538),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[17] ),
    .B1(_12206_),
    .C1(net874),
    .Y(_12208_));
 sky130_fd_sc_hd__o21ai_0 _33143_ (.A1(_11529_),
    .A2(net874),
    .B1(_12208_),
    .Y(_12209_));
 sky130_fd_sc_hd__nand2_1 _33145_ (.A(_12209_),
    .B(net847),
    .Y(_12211_));
 sky130_fd_sc_hd__nand2_1 _33146_ (.A(_12201_),
    .B(_12211_),
    .Y(_12212_));
 sky130_fd_sc_hd__nand2_1 _33147_ (.A(net670),
    .B(_12212_),
    .Y(_12213_));
 sky130_fd_sc_hd__nand2_1 _33148_ (.A(net626),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[17] ),
    .Y(_12214_));
 sky130_fd_sc_hd__a21oi_4 _33149_ (.A1(_12213_),
    .A2(_12214_),
    .B1(net2933),
    .Y(_04128_));
 sky130_fd_sc_hd__nand2_1 _33150_ (.A(net621),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[18] ),
    .Y(_12215_));
 sky130_fd_sc_hd__inv_1 _33151_ (.A(\inst$top.soc.cpu.sink__payload[20] ),
    .Y(_12216_));
 sky130_fd_sc_hd__nor4_1 _33152_ (.A(_12106_),
    .B(_12130_),
    .C(_12180_),
    .D(_12185_),
    .Y(_12217_));
 sky130_fd_sc_hd__nand2_1 _33153_ (.A(_12104_),
    .B(_12217_),
    .Y(_12218_));
 sky130_fd_sc_hd__xor2_1 _33154_ (.A(_12216_),
    .B(_12218_),
    .X(_12219_));
 sky130_fd_sc_hd__nand2_1 _33155_ (.A(net741),
    .B(_12219_),
    .Y(_12220_));
 sky130_fd_sc_hd__nand2_1 _33156_ (.A(_03340_),
    .B(_03342_),
    .Y(_12221_));
 sky130_fd_sc_hd__nor4_1 _33157_ (.A(_12049_),
    .B(_12109_),
    .C(_12165_),
    .D(_12221_),
    .Y(_12222_));
 sky130_fd_sc_hd__nand2_1 _33158_ (.A(_03312_),
    .B(_03314_),
    .Y(_12223_));
 sky130_fd_sc_hd__nor2_1 _33159_ (.A(_12223_),
    .B(_11978_),
    .Y(_12224_));
 sky130_fd_sc_hd__nor2_1 _33160_ (.A(_11971_),
    .B(_11982_),
    .Y(_12225_));
 sky130_fd_sc_hd__nand4_1 _33161_ (.A(_12222_),
    .B(_12224_),
    .C(_02546_),
    .D(_12225_),
    .Y(_12226_));
 sky130_fd_sc_hd__nor2_1 _33162_ (.A(_12165_),
    .B(_12221_),
    .Y(_12227_));
 sky130_fd_sc_hd__a21oi_1 _33163_ (.A1(_03342_),
    .A2(_03339_),
    .B1(_03341_),
    .Y(_12228_));
 sky130_fd_sc_hd__o21ai_0 _33164_ (.A1(_12221_),
    .A2(_12166_),
    .B1(_12228_),
    .Y(_12229_));
 sky130_fd_sc_hd__a21oi_1 _33165_ (.A1(_12111_),
    .A2(_12227_),
    .B1(_12229_),
    .Y(_12230_));
 sky130_fd_sc_hd__o21ai_0 _33166_ (.A1(_11978_),
    .A2(_11975_),
    .B1(_11972_),
    .Y(_12231_));
 sky130_fd_sc_hd__nand2_1 _33167_ (.A(_12231_),
    .B(_12225_),
    .Y(_12232_));
 sky130_fd_sc_hd__a21boi_0 _33168_ (.A1(_11970_),
    .A2(_11983_),
    .B1_N(_11985_),
    .Y(_12233_));
 sky130_fd_sc_hd__nand2_1 _33169_ (.A(_12232_),
    .B(_12233_),
    .Y(_12234_));
 sky130_fd_sc_hd__nand2_1 _33170_ (.A(_12234_),
    .B(_12222_),
    .Y(_12235_));
 sky130_fd_sc_hd__nand3_1 _33171_ (.A(_12226_),
    .B(_12230_),
    .C(_12235_),
    .Y(_12236_));
 sky130_fd_sc_hd__xnor2_1 _33172_ (.A(_03344_),
    .B(_12236_),
    .Y(_12237_));
 sky130_fd_sc_hd__inv_1 _33173_ (.A(_12237_),
    .Y(_12238_));
 sky130_fd_sc_hd__nand3_1 _33174_ (.A(net791),
    .B(net832),
    .C(_12238_),
    .Y(_12239_));
 sky130_fd_sc_hd__nand3_1 _33175_ (.A(_12220_),
    .B(_12239_),
    .C(net814),
    .Y(_12240_));
 sky130_fd_sc_hd__nor2_1 _33176_ (.A(\inst$top.soc.cpu.sink__payload$6[20] ),
    .B(net814),
    .Y(_12241_));
 sky130_fd_sc_hd__nor2_1 _33177_ (.A(net847),
    .B(_12241_),
    .Y(_12242_));
 sky130_fd_sc_hd__nand2_1 _33178_ (.A(_12240_),
    .B(_12242_),
    .Y(_12243_));
 sky130_fd_sc_hd__inv_1 _33179_ (.A(\inst$top.soc.cpu.sink__payload$12[20] ),
    .Y(_12244_));
 sky130_fd_sc_hd__nand3_1 _33180_ (.A(net1821),
    .B(\inst$top.soc.cpu.sink__payload$18[200] ),
    .C(net1838),
    .Y(_12245_));
 sky130_fd_sc_hd__o211ai_1 _33181_ (.A1(_12244_),
    .A2(net1815),
    .B1(net2538),
    .C1(_12245_),
    .Y(_12246_));
 sky130_fd_sc_hd__o211ai_1 _33182_ (.A1(net2538),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[18] ),
    .B1(_12246_),
    .C1(net873),
    .Y(_12247_));
 sky130_fd_sc_hd__o21ai_0 _33183_ (.A1(_05695_),
    .A2(net873),
    .B1(_12247_),
    .Y(_12248_));
 sky130_fd_sc_hd__nand2_1 _33184_ (.A(_12248_),
    .B(net847),
    .Y(_12249_));
 sky130_fd_sc_hd__nand2_1 _33185_ (.A(_12243_),
    .B(_12249_),
    .Y(_12250_));
 sky130_fd_sc_hd__nand3_1 _33186_ (.A(_12250_),
    .B(net663),
    .C(net753),
    .Y(_12251_));
 sky130_fd_sc_hd__a21oi_2 _33187_ (.A1(_12215_),
    .A2(_12251_),
    .B1(net2934),
    .Y(_04129_));
 sky130_fd_sc_hd__nand2_1 _33188_ (.A(net626),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[19] ),
    .Y(_12252_));
 sky130_fd_sc_hd__nor2_1 _33189_ (.A(_12216_),
    .B(_12184_),
    .Y(_12253_));
 sky130_fd_sc_hd__xor2_1 _33190_ (.A(\inst$top.soc.cpu.sink__payload[21] ),
    .B(_12253_),
    .X(_12254_));
 sky130_fd_sc_hd__nand2_1 _33191_ (.A(net741),
    .B(_12254_),
    .Y(_12255_));
 sky130_fd_sc_hd__nand2_1 _33192_ (.A(_03342_),
    .B(_03344_),
    .Y(_12256_));
 sky130_fd_sc_hd__a21oi_1 _33193_ (.A1(_03344_),
    .A2(_03341_),
    .B1(_03343_),
    .Y(_12257_));
 sky130_fd_sc_hd__o21ai_0 _33194_ (.A1(_12256_),
    .A2(_12192_),
    .B1(_12257_),
    .Y(_12258_));
 sky130_fd_sc_hd__nor3_1 _33195_ (.A(_12191_),
    .B(_12256_),
    .C(_12142_),
    .Y(_12259_));
 sky130_fd_sc_hd__nor2_1 _33196_ (.A(_12258_),
    .B(_12259_),
    .Y(_12260_));
 sky130_fd_sc_hd__xnor2_1 _33197_ (.A(_03346_),
    .B(_12260_),
    .Y(_12261_));
 sky130_fd_sc_hd__nand3_1 _33198_ (.A(net791),
    .B(net832),
    .C(_12261_),
    .Y(_12262_));
 sky130_fd_sc_hd__nand3_1 _33199_ (.A(_12255_),
    .B(_12262_),
    .C(net814),
    .Y(_12263_));
 sky130_fd_sc_hd__nor2_1 _33200_ (.A(\inst$top.soc.cpu.sink__payload$6[21] ),
    .B(net814),
    .Y(_12264_));
 sky130_fd_sc_hd__nor2_1 _33201_ (.A(net847),
    .B(_12264_),
    .Y(_12265_));
 sky130_fd_sc_hd__nand2_1 _33202_ (.A(_12263_),
    .B(_12265_),
    .Y(_12266_));
 sky130_fd_sc_hd__nand2_1 _33203_ (.A(\inst$top.soc.cpu.sink__payload$12[21] ),
    .B(_02862_),
    .Y(_12267_));
 sky130_fd_sc_hd__o311ai_0 _33204_ (.A1(_02862_),
    .A2(_11792_),
    .A3(_20257_),
    .B1(net2539),
    .C1(_12267_),
    .Y(_12268_));
 sky130_fd_sc_hd__o211ai_1 _33205_ (.A1(net2538),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[19] ),
    .B1(_12268_),
    .C1(net873),
    .Y(_12269_));
 sky130_fd_sc_hd__o21ai_0 _33206_ (.A1(_11534_),
    .A2(net873),
    .B1(_12269_),
    .Y(_12270_));
 sky130_fd_sc_hd__nand2_1 _33207_ (.A(_12270_),
    .B(net847),
    .Y(_12271_));
 sky130_fd_sc_hd__nand2_1 _33208_ (.A(_12266_),
    .B(_12271_),
    .Y(_12272_));
 sky130_fd_sc_hd__nand3_1 _33209_ (.A(_12272_),
    .B(net663),
    .C(net753),
    .Y(_12273_));
 sky130_fd_sc_hd__a21oi_2 _33210_ (.A1(_12252_),
    .A2(_12273_),
    .B1(net2933),
    .Y(_04130_));
 sky130_fd_sc_hd__nand2_1 _33211_ (.A(net621),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[1] ),
    .Y(_12274_));
 sky130_fd_sc_hd__nand2_1 _33212_ (.A(net740),
    .B(_02867_),
    .Y(_12275_));
 sky130_fd_sc_hd__nand3_1 _33213_ (.A(net790),
    .B(\inst$top.soc.cpu.d_branch_target[3] ),
    .C(net831),
    .Y(_12276_));
 sky130_fd_sc_hd__nand3_1 _33214_ (.A(_12275_),
    .B(_12276_),
    .C(net813),
    .Y(_12277_));
 sky130_fd_sc_hd__nor2_1 _33215_ (.A(\inst$top.soc.cpu.sink__payload$6[3] ),
    .B(net813),
    .Y(_12278_));
 sky130_fd_sc_hd__nor2_1 _33216_ (.A(net846),
    .B(_12278_),
    .Y(_12279_));
 sky130_fd_sc_hd__nand2_1 _33217_ (.A(_12277_),
    .B(_12279_),
    .Y(_12280_));
 sky130_fd_sc_hd__nand2_1 _33218_ (.A(\inst$top.soc.cpu.sink__payload$12[3] ),
    .B(_02862_),
    .Y(_12281_));
 sky130_fd_sc_hd__o311ai_0 _33219_ (.A1(_02862_),
    .A2(_11858_),
    .A3(_20257_),
    .B1(net2537),
    .C1(_12281_),
    .Y(_12282_));
 sky130_fd_sc_hd__o211ai_1 _33220_ (.A1(net2540),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[1] ),
    .B1(_12282_),
    .C1(net872),
    .Y(_12283_));
 sky130_fd_sc_hd__o21ai_0 _33221_ (.A1(_20512_),
    .A2(net872),
    .B1(_12283_),
    .Y(_12284_));
 sky130_fd_sc_hd__nand2_1 _33222_ (.A(_12284_),
    .B(net846),
    .Y(_12285_));
 sky130_fd_sc_hd__nand2_1 _33223_ (.A(_12280_),
    .B(_12285_),
    .Y(_12286_));
 sky130_fd_sc_hd__nand3_1 _33224_ (.A(_12286_),
    .B(net663),
    .C(net753),
    .Y(_12287_));
 sky130_fd_sc_hd__a21oi_4 _33225_ (.A1(_12274_),
    .A2(_12287_),
    .B1(net2935),
    .Y(_04131_));
 sky130_fd_sc_hd__nand2_1 _33226_ (.A(net636),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[20] ),
    .Y(_12288_));
 sky130_fd_sc_hd__inv_1 _33227_ (.A(\inst$top.soc.cpu.sink__payload[22] ),
    .Y(_12289_));
 sky130_fd_sc_hd__nand2_1 _33228_ (.A(\inst$top.soc.cpu.sink__payload[20] ),
    .B(\inst$top.soc.cpu.sink__payload[21] ),
    .Y(_12290_));
 sky130_fd_sc_hd__inv_1 _33229_ (.A(_12290_),
    .Y(_12291_));
 sky130_fd_sc_hd__nand4_1 _33230_ (.A(_12162_),
    .B(\inst$top.soc.cpu.sink__payload[18] ),
    .C(\inst$top.soc.cpu.sink__payload[19] ),
    .D(_12291_),
    .Y(_12292_));
 sky130_fd_sc_hd__xor2_1 _33231_ (.A(_12289_),
    .B(_12292_),
    .X(_12293_));
 sky130_fd_sc_hd__nand2_1 _33232_ (.A(net742),
    .B(_12293_),
    .Y(_12294_));
 sky130_fd_sc_hd__nand3_1 _33233_ (.A(_12236_),
    .B(_03344_),
    .C(_03346_),
    .Y(_12295_));
 sky130_fd_sc_hd__a21oi_1 _33234_ (.A1(_03346_),
    .A2(_03343_),
    .B1(_03345_),
    .Y(_12296_));
 sky130_fd_sc_hd__nand2_1 _33235_ (.A(_12295_),
    .B(_12296_),
    .Y(_12297_));
 sky130_fd_sc_hd__xor2_1 _33236_ (.A(_03348_),
    .B(_12297_),
    .X(_12298_));
 sky130_fd_sc_hd__nand3_1 _33237_ (.A(net792),
    .B(net833),
    .C(_12298_),
    .Y(_12299_));
 sky130_fd_sc_hd__nand3_1 _33238_ (.A(_12294_),
    .B(_12299_),
    .C(net816),
    .Y(_12300_));
 sky130_fd_sc_hd__nor2_1 _33239_ (.A(\inst$top.soc.cpu.sink__payload$6[22] ),
    .B(net816),
    .Y(_12301_));
 sky130_fd_sc_hd__nor2_1 _33240_ (.A(net850),
    .B(_12301_),
    .Y(_12302_));
 sky130_fd_sc_hd__nand2_1 _33241_ (.A(_12300_),
    .B(_12302_),
    .Y(_12303_));
 sky130_fd_sc_hd__inv_1 _33242_ (.A(\inst$top.soc.cpu.sink__payload$12[22] ),
    .Y(_12304_));
 sky130_fd_sc_hd__nand3_1 _33243_ (.A(net1818),
    .B(\inst$top.soc.cpu.sink__payload$18[202] ),
    .C(net1839),
    .Y(_12305_));
 sky130_fd_sc_hd__o211ai_1 _33244_ (.A1(_12304_),
    .A2(net1818),
    .B1(net2543),
    .C1(_12305_),
    .Y(_12306_));
 sky130_fd_sc_hd__o211ai_1 _33245_ (.A1(net2543),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[20] ),
    .B1(_12306_),
    .C1(net878),
    .Y(_12307_));
 sky130_fd_sc_hd__o21ai_0 _33246_ (.A1(_05734_),
    .A2(net878),
    .B1(_12307_),
    .Y(_12308_));
 sky130_fd_sc_hd__nand2_1 _33247_ (.A(_12308_),
    .B(net850),
    .Y(_12309_));
 sky130_fd_sc_hd__nand2_1 _33248_ (.A(_12303_),
    .B(_12309_),
    .Y(_12310_));
 sky130_fd_sc_hd__nand3_1 _33249_ (.A(_12310_),
    .B(net664),
    .C(net754),
    .Y(_12311_));
 sky130_fd_sc_hd__a21oi_2 _33250_ (.A1(_12288_),
    .A2(_12311_),
    .B1(net2945),
    .Y(_04132_));
 sky130_fd_sc_hd__inv_1 _33251_ (.A(\inst$top.soc.cpu.sink__payload[23] ),
    .Y(_12312_));
 sky130_fd_sc_hd__nand2_1 _33252_ (.A(\inst$top.soc.cpu.sink__payload[21] ),
    .B(\inst$top.soc.cpu.sink__payload[22] ),
    .Y(_12313_));
 sky130_fd_sc_hd__nor3_1 _33253_ (.A(_12185_),
    .B(_12216_),
    .C(_12313_),
    .Y(_12314_));
 sky130_fd_sc_hd__nand2_1 _33254_ (.A(_12183_),
    .B(_12314_),
    .Y(_12315_));
 sky130_fd_sc_hd__xor2_1 _33255_ (.A(_12312_),
    .B(_12315_),
    .X(_12316_));
 sky130_fd_sc_hd__inv_1 _33256_ (.A(_12316_),
    .Y(_12317_));
 sky130_fd_sc_hd__nand2_1 _33257_ (.A(net743),
    .B(_12317_),
    .Y(_12318_));
 sky130_fd_sc_hd__inv_1 _33258_ (.A(_03350_),
    .Y(_12319_));
 sky130_fd_sc_hd__nand2_1 _33259_ (.A(_03346_),
    .B(_03348_),
    .Y(_12320_));
 sky130_fd_sc_hd__nor2_1 _33260_ (.A(_12256_),
    .B(_12320_),
    .Y(_12321_));
 sky130_fd_sc_hd__a21oi_1 _33261_ (.A1(_03348_),
    .A2(_03345_),
    .B1(_03347_),
    .Y(_12322_));
 sky130_fd_sc_hd__o21ai_0 _33262_ (.A1(_12320_),
    .A2(_12257_),
    .B1(_12322_),
    .Y(_12323_));
 sky130_fd_sc_hd__a21o_1 _33263_ (.A1(_12193_),
    .A2(_12321_),
    .B1(_12323_),
    .X(_12324_));
 sky130_fd_sc_hd__xor2_1 _33264_ (.A(_12319_),
    .B(_12324_),
    .X(_12325_));
 sky130_fd_sc_hd__nand3_1 _33265_ (.A(net793),
    .B(net834),
    .C(_12325_),
    .Y(_12326_));
 sky130_fd_sc_hd__nand3_1 _33266_ (.A(_12318_),
    .B(_12326_),
    .C(net817),
    .Y(_12327_));
 sky130_fd_sc_hd__nand2_1 _33267_ (.A(_20362_),
    .B(\inst$top.soc.cpu.sink__payload$6[23] ),
    .Y(_12328_));
 sky130_fd_sc_hd__nand2_1 _33268_ (.A(_12327_),
    .B(_12328_),
    .Y(_12329_));
 sky130_fd_sc_hd__nand2_1 _33269_ (.A(_12329_),
    .B(net871),
    .Y(_12330_));
 sky130_fd_sc_hd__nand3_1 _33270_ (.A(net1818),
    .B(\inst$top.soc.cpu.sink__payload$18[203] ),
    .C(net1840),
    .Y(_12331_));
 sky130_fd_sc_hd__o211ai_1 _33271_ (.A1(_05749_),
    .A2(net1818),
    .B1(net2543),
    .C1(_12331_),
    .Y(_12332_));
 sky130_fd_sc_hd__o211ai_1 _33272_ (.A1(net2543),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[21] ),
    .B1(_12332_),
    .C1(net878),
    .Y(_12333_));
 sky130_fd_sc_hd__o21ai_0 _33273_ (.A1(_11539_),
    .A2(net878),
    .B1(_12333_),
    .Y(_12334_));
 sky130_fd_sc_hd__nand2_1 _33274_ (.A(_12334_),
    .B(net851),
    .Y(_12335_));
 sky130_fd_sc_hd__nand2_1 _33275_ (.A(_12330_),
    .B(_12335_),
    .Y(_12336_));
 sky130_fd_sc_hd__nand2_1 _33276_ (.A(net677),
    .B(_12336_),
    .Y(_12337_));
 sky130_fd_sc_hd__nand2_1 _33277_ (.A(net636),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[21] ),
    .Y(_12338_));
 sky130_fd_sc_hd__a21oi_4 _33278_ (.A1(_12337_),
    .A2(_12338_),
    .B1(net2944),
    .Y(_04133_));
 sky130_fd_sc_hd__inv_1 _33279_ (.A(\inst$top.soc.cpu.sink__payload[24] ),
    .Y(_12339_));
 sky130_fd_sc_hd__nor4_1 _33280_ (.A(_12289_),
    .B(_12312_),
    .C(_12290_),
    .D(_12218_),
    .Y(_12340_));
 sky130_fd_sc_hd__xor2_1 _33281_ (.A(_12339_),
    .B(_12340_),
    .X(_12341_));
 sky130_fd_sc_hd__nand2_1 _33282_ (.A(net743),
    .B(_12341_),
    .Y(_12342_));
 sky130_fd_sc_hd__inv_1 _33283_ (.A(_03352_),
    .Y(_12343_));
 sky130_fd_sc_hd__nand2_1 _33284_ (.A(_03348_),
    .B(_03350_),
    .Y(_12344_));
 sky130_fd_sc_hd__inv_1 _33285_ (.A(_12344_),
    .Y(_12345_));
 sky130_fd_sc_hd__nand2_1 _33286_ (.A(_12297_),
    .B(_12345_),
    .Y(_12346_));
 sky130_fd_sc_hd__a21oi_1 _33287_ (.A1(_03350_),
    .A2(_03347_),
    .B1(_03349_),
    .Y(_12347_));
 sky130_fd_sc_hd__nand2_1 _33288_ (.A(_12346_),
    .B(_12347_),
    .Y(_12348_));
 sky130_fd_sc_hd__xor2_1 _33289_ (.A(_12343_),
    .B(_12348_),
    .X(_12349_));
 sky130_fd_sc_hd__nand3_1 _33290_ (.A(net793),
    .B(net834),
    .C(_12349_),
    .Y(_12350_));
 sky130_fd_sc_hd__nand3_1 _33291_ (.A(_12342_),
    .B(_12350_),
    .C(net817),
    .Y(_12351_));
 sky130_fd_sc_hd__nand2_1 _33292_ (.A(_20362_),
    .B(\inst$top.soc.cpu.sink__payload$6[24] ),
    .Y(_12352_));
 sky130_fd_sc_hd__nand2_1 _33293_ (.A(_12351_),
    .B(_12352_),
    .Y(_12353_));
 sky130_fd_sc_hd__nand2_1 _33294_ (.A(_12353_),
    .B(net871),
    .Y(_12354_));
 sky130_fd_sc_hd__nand3_1 _33295_ (.A(net1818),
    .B(\inst$top.soc.cpu.sink__payload$18[204] ),
    .C(net1840),
    .Y(_12355_));
 sky130_fd_sc_hd__o211ai_1 _33296_ (.A1(_05768_),
    .A2(net1819),
    .B1(net2543),
    .C1(_12355_),
    .Y(_12356_));
 sky130_fd_sc_hd__o211ai_1 _33297_ (.A1(net2543),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[22] ),
    .B1(_12356_),
    .C1(net877),
    .Y(_12357_));
 sky130_fd_sc_hd__o21ai_0 _33298_ (.A1(_11541_),
    .A2(net877),
    .B1(_12357_),
    .Y(_12358_));
 sky130_fd_sc_hd__nand2_1 _33299_ (.A(_12358_),
    .B(net851),
    .Y(_12359_));
 sky130_fd_sc_hd__nand2_1 _33300_ (.A(_12354_),
    .B(_12359_),
    .Y(_12360_));
 sky130_fd_sc_hd__nand2_1 _33301_ (.A(net677),
    .B(_12360_),
    .Y(_12361_));
 sky130_fd_sc_hd__nand2_1 _33302_ (.A(net635),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[22] ),
    .Y(_12362_));
 sky130_fd_sc_hd__a21oi_4 _33303_ (.A1(_12361_),
    .A2(_12362_),
    .B1(net2945),
    .Y(_04134_));
 sky130_fd_sc_hd__inv_1 _33304_ (.A(\inst$top.soc.cpu.sink__payload[25] ),
    .Y(_12363_));
 sky130_fd_sc_hd__nor3_1 _33305_ (.A(_12312_),
    .B(_12339_),
    .C(_12313_),
    .Y(_12364_));
 sky130_fd_sc_hd__nand2_1 _33306_ (.A(_12253_),
    .B(_12364_),
    .Y(_12365_));
 sky130_fd_sc_hd__xor2_1 _33307_ (.A(_12363_),
    .B(_12365_),
    .X(_12366_));
 sky130_fd_sc_hd__inv_1 _33308_ (.A(_12366_),
    .Y(_12367_));
 sky130_fd_sc_hd__nand2_1 _33309_ (.A(net742),
    .B(_12367_),
    .Y(_12368_));
 sky130_fd_sc_hd__nand2_1 _33310_ (.A(_03350_),
    .B(_03352_),
    .Y(_12369_));
 sky130_fd_sc_hd__nor4_1 _33311_ (.A(_12191_),
    .B(_12256_),
    .C(_12320_),
    .D(_12369_),
    .Y(_12370_));
 sky130_fd_sc_hd__nand2_1 _33312_ (.A(_12141_),
    .B(_12370_),
    .Y(_12371_));
 sky130_fd_sc_hd__nor2_1 _33313_ (.A(_12320_),
    .B(_12369_),
    .Y(_12372_));
 sky130_fd_sc_hd__a21oi_1 _33314_ (.A1(_03352_),
    .A2(_03349_),
    .B1(_03351_),
    .Y(_12373_));
 sky130_fd_sc_hd__o21ai_0 _33315_ (.A1(_12369_),
    .A2(_12322_),
    .B1(_12373_),
    .Y(_12374_));
 sky130_fd_sc_hd__a21oi_1 _33316_ (.A1(_12258_),
    .A2(_12372_),
    .B1(_12374_),
    .Y(_12375_));
 sky130_fd_sc_hd__nand3_1 _33317_ (.A(_12024_),
    .B(_12370_),
    .C(_12136_),
    .Y(_12376_));
 sky130_fd_sc_hd__nand3_1 _33318_ (.A(_12371_),
    .B(_12375_),
    .C(_12376_),
    .Y(_12377_));
 sky130_fd_sc_hd__xnor2_2 _33319_ (.A(_03354_),
    .B(_12377_),
    .Y(_12378_));
 sky130_fd_sc_hd__nand3_1 _33320_ (.A(net792),
    .B(net833),
    .C(_12378_),
    .Y(_12379_));
 sky130_fd_sc_hd__nand3_1 _33321_ (.A(_12368_),
    .B(_12379_),
    .C(net816),
    .Y(_12380_));
 sky130_fd_sc_hd__nand2_1 _33322_ (.A(net838),
    .B(\inst$top.soc.cpu.sink__payload$6[25] ),
    .Y(_12381_));
 sky130_fd_sc_hd__nand2_1 _33323_ (.A(_12380_),
    .B(_12381_),
    .Y(_12382_));
 sky130_fd_sc_hd__nand2_1 _33324_ (.A(_12382_),
    .B(net871),
    .Y(_12383_));
 sky130_fd_sc_hd__inv_1 _33325_ (.A(\inst$top.soc.cpu.sink__payload$12[25] ),
    .Y(_12384_));
 sky130_fd_sc_hd__nand3_1 _33326_ (.A(net1816),
    .B(\inst$top.soc.cpu.sink__payload$18[205] ),
    .C(net1838),
    .Y(_12385_));
 sky130_fd_sc_hd__o211ai_1 _33327_ (.A1(_12384_),
    .A2(net1816),
    .B1(net2540),
    .C1(_12385_),
    .Y(_12386_));
 sky130_fd_sc_hd__o211ai_1 _33328_ (.A1(net2537),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[23] ),
    .B1(_12386_),
    .C1(net875),
    .Y(_12387_));
 sky130_fd_sc_hd__o21ai_0 _33329_ (.A1(_11543_),
    .A2(net875),
    .B1(_12387_),
    .Y(_12388_));
 sky130_fd_sc_hd__nand2_1 _33330_ (.A(_12388_),
    .B(net846),
    .Y(_12389_));
 sky130_fd_sc_hd__nand2_1 _33331_ (.A(_12383_),
    .B(_12389_),
    .Y(_12390_));
 sky130_fd_sc_hd__nand2_1 _33332_ (.A(net676),
    .B(_12390_),
    .Y(_12391_));
 sky130_fd_sc_hd__nand2_1 _33333_ (.A(net627),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[23] ),
    .Y(_12392_));
 sky130_fd_sc_hd__a21oi_4 _33334_ (.A1(_12391_),
    .A2(_12392_),
    .B1(net2944),
    .Y(_04135_));
 sky130_fd_sc_hd__nor4_1 _33335_ (.A(_12289_),
    .B(_12312_),
    .C(_12339_),
    .D(_12363_),
    .Y(_12393_));
 sky130_fd_sc_hd__inv_1 _33336_ (.A(_12393_),
    .Y(_12394_));
 sky130_fd_sc_hd__nor2_1 _33337_ (.A(_12394_),
    .B(_12292_),
    .Y(_12395_));
 sky130_fd_sc_hd__xor2_1 _33338_ (.A(\inst$top.soc.cpu.sink__payload[26] ),
    .B(_12395_),
    .X(_12396_));
 sky130_fd_sc_hd__inv_1 _33339_ (.A(_12396_),
    .Y(_12397_));
 sky130_fd_sc_hd__nand2_1 _33340_ (.A(net743),
    .B(_12397_),
    .Y(_12398_));
 sky130_fd_sc_hd__nand2_1 _33341_ (.A(_03344_),
    .B(_03346_),
    .Y(_12399_));
 sky130_fd_sc_hd__nor2_1 _33342_ (.A(_12221_),
    .B(_12399_),
    .Y(_12400_));
 sky130_fd_sc_hd__nand2_1 _33343_ (.A(_03352_),
    .B(_03354_),
    .Y(_12401_));
 sky130_fd_sc_hd__nor2_1 _33344_ (.A(_12344_),
    .B(_12401_),
    .Y(_12402_));
 sky130_fd_sc_hd__nand2_1 _33345_ (.A(_12400_),
    .B(_12402_),
    .Y(_12403_));
 sky130_fd_sc_hd__nor2_1 _33346_ (.A(_12109_),
    .B(_12165_),
    .Y(_12404_));
 sky130_fd_sc_hd__o21ai_0 _33347_ (.A1(_12165_),
    .A2(_12110_),
    .B1(_12166_),
    .Y(_12405_));
 sky130_fd_sc_hd__a21oi_1 _33348_ (.A1(_12052_),
    .A2(_12404_),
    .B1(_12405_),
    .Y(_12406_));
 sky130_fd_sc_hd__o21ai_0 _33349_ (.A1(_12399_),
    .A2(_12228_),
    .B1(_12296_),
    .Y(_12407_));
 sky130_fd_sc_hd__a21oi_1 _33350_ (.A1(_03354_),
    .A2(_03351_),
    .B1(_03353_),
    .Y(_12408_));
 sky130_fd_sc_hd__o21ai_0 _33351_ (.A1(_12401_),
    .A2(_12347_),
    .B1(_12408_),
    .Y(_12409_));
 sky130_fd_sc_hd__a21oi_1 _33352_ (.A1(_12407_),
    .A2(_12402_),
    .B1(_12409_),
    .Y(_12410_));
 sky130_fd_sc_hd__nor4_1 _33353_ (.A(_11982_),
    .B(_12049_),
    .C(_12109_),
    .D(_12165_),
    .Y(_12411_));
 sky130_fd_sc_hd__nand4_1 _33354_ (.A(_12411_),
    .B(_11981_),
    .C(_12400_),
    .D(_12402_),
    .Y(_12412_));
 sky130_fd_sc_hd__o211ai_1 _33355_ (.A1(_12403_),
    .A2(_12406_),
    .B1(_12410_),
    .C1(_12412_),
    .Y(_12413_));
 sky130_fd_sc_hd__xnor2_1 _33356_ (.A(_03356_),
    .B(_12413_),
    .Y(_12414_));
 sky130_fd_sc_hd__nand3_1 _33357_ (.A(net793),
    .B(net834),
    .C(_12414_),
    .Y(_12415_));
 sky130_fd_sc_hd__nand3_1 _33358_ (.A(_12398_),
    .B(_12415_),
    .C(net817),
    .Y(_12416_));
 sky130_fd_sc_hd__nand2_1 _33359_ (.A(net838),
    .B(\inst$top.soc.cpu.sink__payload$6[26] ),
    .Y(_12417_));
 sky130_fd_sc_hd__nand2_1 _33360_ (.A(_12416_),
    .B(_12417_),
    .Y(_12418_));
 sky130_fd_sc_hd__nand2_1 _33361_ (.A(_12418_),
    .B(net871),
    .Y(_12419_));
 sky130_fd_sc_hd__inv_1 _33362_ (.A(\inst$top.soc.cpu.sink__payload$12[26] ),
    .Y(_12420_));
 sky130_fd_sc_hd__nand3_1 _33363_ (.A(net1820),
    .B(\inst$top.soc.cpu.sink__payload$18[206] ),
    .C(net1839),
    .Y(_12421_));
 sky130_fd_sc_hd__o211ai_1 _33364_ (.A1(_12420_),
    .A2(net1819),
    .B1(net2542),
    .C1(_12421_),
    .Y(_12422_));
 sky130_fd_sc_hd__o211ai_1 _33365_ (.A1(net2542),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[24] ),
    .B1(_12422_),
    .C1(net878),
    .Y(_12423_));
 sky130_fd_sc_hd__o21ai_0 _33366_ (.A1(_05814_),
    .A2(net877),
    .B1(_12423_),
    .Y(_12424_));
 sky130_fd_sc_hd__nand2_1 _33367_ (.A(_12424_),
    .B(net850),
    .Y(_12425_));
 sky130_fd_sc_hd__nand2_1 _33368_ (.A(_12419_),
    .B(_12425_),
    .Y(_12426_));
 sky130_fd_sc_hd__nand2_1 _33369_ (.A(net682),
    .B(_12426_),
    .Y(_12427_));
 sky130_fd_sc_hd__nand2_1 _33370_ (.A(net638),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[24] ),
    .Y(_12428_));
 sky130_fd_sc_hd__a21oi_4 _33371_ (.A1(_12427_),
    .A2(_12428_),
    .B1(net2948),
    .Y(_04136_));
 sky130_fd_sc_hd__nor2_1 _33372_ (.A(_12138_),
    .B(_12191_),
    .Y(_12429_));
 sky130_fd_sc_hd__o21ai_0 _33373_ (.A1(_12191_),
    .A2(_12139_),
    .B1(_12192_),
    .Y(_12430_));
 sky130_fd_sc_hd__a21oi_1 _33374_ (.A1(_12081_),
    .A2(_12429_),
    .B1(_12430_),
    .Y(_12431_));
 sky130_fd_sc_hd__inv_1 _33375_ (.A(_12321_),
    .Y(_12432_));
 sky130_fd_sc_hd__nand2_1 _33376_ (.A(_03354_),
    .B(_03356_),
    .Y(_12433_));
 sky130_fd_sc_hd__nor2_1 _33377_ (.A(_12369_),
    .B(_12433_),
    .Y(_12434_));
 sky130_fd_sc_hd__inv_1 _33378_ (.A(_12434_),
    .Y(_12435_));
 sky130_fd_sc_hd__nor2_1 _33379_ (.A(_12432_),
    .B(_12435_),
    .Y(_12436_));
 sky130_fd_sc_hd__inv_1 _33380_ (.A(_12436_),
    .Y(_12437_));
 sky130_fd_sc_hd__a21oi_1 _33381_ (.A1(_03356_),
    .A2(_03353_),
    .B1(_03355_),
    .Y(_12438_));
 sky130_fd_sc_hd__o21ai_0 _33382_ (.A1(_12433_),
    .A2(_12373_),
    .B1(_12438_),
    .Y(_12439_));
 sky130_fd_sc_hd__a21oi_1 _33383_ (.A1(_12323_),
    .A2(_12434_),
    .B1(_12439_),
    .Y(_12440_));
 sky130_fd_sc_hd__nand4_1 _33384_ (.A(_12027_),
    .B(_12079_),
    .C(_12429_),
    .D(_12436_),
    .Y(_12441_));
 sky130_fd_sc_hd__o211ai_1 _33385_ (.A1(_12431_),
    .A2(_12437_),
    .B1(_12440_),
    .C1(_12441_),
    .Y(_12442_));
 sky130_fd_sc_hd__inv_1 _33386_ (.A(_12442_),
    .Y(_12443_));
 sky130_fd_sc_hd__inv_1 _33387_ (.A(_03358_),
    .Y(_12444_));
 sky130_fd_sc_hd__nand2_1 _33388_ (.A(_12443_),
    .B(_12444_),
    .Y(_12445_));
 sky130_fd_sc_hd__nand2_1 _33389_ (.A(_12442_),
    .B(_03358_),
    .Y(_12446_));
 sky130_fd_sc_hd__nand2_1 _33390_ (.A(_12445_),
    .B(_12446_),
    .Y(_12447_));
 sky130_fd_sc_hd__nand3_1 _33391_ (.A(net793),
    .B(_12447_),
    .C(net833),
    .Y(_12448_));
 sky130_fd_sc_hd__nand4_1 _33392_ (.A(\inst$top.soc.cpu.sink__payload[23] ),
    .B(\inst$top.soc.cpu.sink__payload[24] ),
    .C(\inst$top.soc.cpu.sink__payload[25] ),
    .D(\inst$top.soc.cpu.sink__payload[26] ),
    .Y(_12449_));
 sky130_fd_sc_hd__nor2_1 _33393_ (.A(_12449_),
    .B(_12315_),
    .Y(_12450_));
 sky130_fd_sc_hd__xor2_1 _33394_ (.A(\inst$top.soc.cpu.sink__payload[27] ),
    .B(_12450_),
    .X(_12451_));
 sky130_fd_sc_hd__inv_1 _33395_ (.A(_12451_),
    .Y(_12452_));
 sky130_fd_sc_hd__nand2_1 _33396_ (.A(net743),
    .B(_12452_),
    .Y(_12453_));
 sky130_fd_sc_hd__nand3_1 _33397_ (.A(_12448_),
    .B(_12453_),
    .C(net817),
    .Y(_12454_));
 sky130_fd_sc_hd__nand2_1 _33398_ (.A(net838),
    .B(\inst$top.soc.cpu.sink__payload$6[27] ),
    .Y(_12455_));
 sky130_fd_sc_hd__nand2_1 _33399_ (.A(_12454_),
    .B(_12455_),
    .Y(_12456_));
 sky130_fd_sc_hd__nand2_1 _33400_ (.A(_12456_),
    .B(net871),
    .Y(_12457_));
 sky130_fd_sc_hd__nand3_1 _33401_ (.A(net1820),
    .B(\inst$top.soc.cpu.sink__payload$18[207] ),
    .C(net1839),
    .Y(_12458_));
 sky130_fd_sc_hd__o211ai_1 _33402_ (.A1(_19947_),
    .A2(net1819),
    .B1(net2542),
    .C1(_12458_),
    .Y(_12459_));
 sky130_fd_sc_hd__o211ai_1 _33403_ (.A1(net2542),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[25] ),
    .B1(_12459_),
    .C1(net878),
    .Y(_12460_));
 sky130_fd_sc_hd__o21ai_0 _33404_ (.A1(_05827_),
    .A2(net877),
    .B1(_12460_),
    .Y(_12461_));
 sky130_fd_sc_hd__nand2_1 _33405_ (.A(_12461_),
    .B(net850),
    .Y(_12462_));
 sky130_fd_sc_hd__nand2_1 _33406_ (.A(_12457_),
    .B(_12462_),
    .Y(_12463_));
 sky130_fd_sc_hd__nand2_1 _33407_ (.A(net682),
    .B(_12463_),
    .Y(_12464_));
 sky130_fd_sc_hd__nand2_1 _33408_ (.A(net638),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[25] ),
    .Y(_12465_));
 sky130_fd_sc_hd__a21oi_4 _33410_ (.A1(_12464_),
    .A2(_12465_),
    .B1(net2948),
    .Y(_04137_));
 sky130_fd_sc_hd__nand2_1 _33411_ (.A(\inst$top.soc.cpu.sink__payload[26] ),
    .B(\inst$top.soc.cpu.sink__payload[27] ),
    .Y(_12467_));
 sky130_fd_sc_hd__nor4_1 _33412_ (.A(_12290_),
    .B(_12394_),
    .C(_12467_),
    .D(_12218_),
    .Y(_12468_));
 sky130_fd_sc_hd__xnor2_1 _33413_ (.A(\inst$top.soc.cpu.sink__payload[28] ),
    .B(_12468_),
    .Y(_12469_));
 sky130_fd_sc_hd__nand2_1 _33414_ (.A(net743),
    .B(_12469_),
    .Y(_12470_));
 sky130_fd_sc_hd__inv_1 _33415_ (.A(_03360_),
    .Y(_12471_));
 sky130_fd_sc_hd__nand3_1 _33416_ (.A(_12413_),
    .B(_03356_),
    .C(_03358_),
    .Y(_12472_));
 sky130_fd_sc_hd__a21oi_1 _33417_ (.A1(_03358_),
    .A2(_03355_),
    .B1(_03357_),
    .Y(_12473_));
 sky130_fd_sc_hd__nand2_1 _33418_ (.A(_12472_),
    .B(_12473_),
    .Y(_12474_));
 sky130_fd_sc_hd__xor2_1 _33419_ (.A(_12471_),
    .B(_12474_),
    .X(_12475_));
 sky130_fd_sc_hd__nand3_1 _33420_ (.A(net793),
    .B(net833),
    .C(_12475_),
    .Y(_12476_));
 sky130_fd_sc_hd__nand3_1 _33421_ (.A(_12470_),
    .B(_12476_),
    .C(net817),
    .Y(_12477_));
 sky130_fd_sc_hd__nand2_1 _33422_ (.A(net838),
    .B(\inst$top.soc.cpu.sink__payload$6[28] ),
    .Y(_12478_));
 sky130_fd_sc_hd__nand2_1 _33423_ (.A(_12477_),
    .B(_12478_),
    .Y(_12479_));
 sky130_fd_sc_hd__nand2_1 _33424_ (.A(_12479_),
    .B(net871),
    .Y(_12480_));
 sky130_fd_sc_hd__inv_1 _33425_ (.A(\inst$top.soc.cpu.sink__payload$12[28] ),
    .Y(_12481_));
 sky130_fd_sc_hd__nand3_1 _33426_ (.A(net1818),
    .B(\inst$top.soc.cpu.sink__payload$18[208] ),
    .C(net1839),
    .Y(_12482_));
 sky130_fd_sc_hd__o211ai_1 _33427_ (.A1(_12481_),
    .A2(net1819),
    .B1(net2542),
    .C1(_12482_),
    .Y(_12483_));
 sky130_fd_sc_hd__o211ai_1 _33428_ (.A1(net2542),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[26] ),
    .B1(_12483_),
    .C1(net877),
    .Y(_12484_));
 sky130_fd_sc_hd__o21ai_0 _33429_ (.A1(_05840_),
    .A2(net877),
    .B1(_12484_),
    .Y(_12485_));
 sky130_fd_sc_hd__nand2_1 _33430_ (.A(_12485_),
    .B(net850),
    .Y(_12486_));
 sky130_fd_sc_hd__nand2_1 _33431_ (.A(_12480_),
    .B(_12486_),
    .Y(_12487_));
 sky130_fd_sc_hd__nand2_1 _33432_ (.A(net682),
    .B(_12487_),
    .Y(_12488_));
 sky130_fd_sc_hd__nand2_1 _33433_ (.A(net635),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[26] ),
    .Y(_12489_));
 sky130_fd_sc_hd__a21oi_4 _33434_ (.A1(_12488_),
    .A2(_12489_),
    .B1(net2945),
    .Y(_04138_));
 sky130_fd_sc_hd__nand2_1 _33435_ (.A(\inst$top.soc.cpu.sink__payload[27] ),
    .B(\inst$top.soc.cpu.sink__payload[28] ),
    .Y(_12490_));
 sky130_fd_sc_hd__nor3_1 _33436_ (.A(_12313_),
    .B(_12490_),
    .C(_12449_),
    .Y(_12491_));
 sky130_fd_sc_hd__nand2_1 _33437_ (.A(_12253_),
    .B(_12491_),
    .Y(_12492_));
 sky130_fd_sc_hd__xnor2_1 _33438_ (.A(\inst$top.soc.cpu.sink__payload[29] ),
    .B(_12492_),
    .Y(_12493_));
 sky130_fd_sc_hd__inv_1 _33439_ (.A(_12493_),
    .Y(_12494_));
 sky130_fd_sc_hd__nand2_1 _33440_ (.A(net743),
    .B(_12494_),
    .Y(_12495_));
 sky130_fd_sc_hd__nand2_1 _33441_ (.A(_03358_),
    .B(_03360_),
    .Y(_12496_));
 sky130_fd_sc_hd__nor2_1 _33442_ (.A(_12433_),
    .B(_12496_),
    .Y(_12497_));
 sky130_fd_sc_hd__a21oi_1 _33443_ (.A1(_03360_),
    .A2(_03357_),
    .B1(_03359_),
    .Y(_12498_));
 sky130_fd_sc_hd__o21ai_0 _33444_ (.A1(_12496_),
    .A2(_12438_),
    .B1(_12498_),
    .Y(_12499_));
 sky130_fd_sc_hd__a21oi_1 _33445_ (.A1(_12377_),
    .A2(_12497_),
    .B1(_12499_),
    .Y(_12500_));
 sky130_fd_sc_hd__xor2_1 _33446_ (.A(_03362_),
    .B(_12500_),
    .X(_12501_));
 sky130_fd_sc_hd__nand3_1 _33447_ (.A(net793),
    .B(net833),
    .C(_12501_),
    .Y(_12502_));
 sky130_fd_sc_hd__nand3_1 _33448_ (.A(_12495_),
    .B(_12502_),
    .C(net817),
    .Y(_12503_));
 sky130_fd_sc_hd__nand2_1 _33449_ (.A(net838),
    .B(\inst$top.soc.cpu.sink__payload$6[29] ),
    .Y(_12504_));
 sky130_fd_sc_hd__nand2_1 _33450_ (.A(_12503_),
    .B(_12504_),
    .Y(_12505_));
 sky130_fd_sc_hd__nand2_1 _33451_ (.A(_12505_),
    .B(net871),
    .Y(_12506_));
 sky130_fd_sc_hd__nand3_1 _33452_ (.A(net1818),
    .B(\inst$top.soc.cpu.sink__payload$18[209] ),
    .C(net1839),
    .Y(_12507_));
 sky130_fd_sc_hd__o211ai_1 _33453_ (.A1(_19920_),
    .A2(net1819),
    .B1(net2542),
    .C1(_12507_),
    .Y(_12508_));
 sky130_fd_sc_hd__o211ai_1 _33454_ (.A1(net2542),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[27] ),
    .B1(_12508_),
    .C1(net877),
    .Y(_12509_));
 sky130_fd_sc_hd__o21ai_0 _33455_ (.A1(_05853_),
    .A2(net877),
    .B1(_12509_),
    .Y(_12510_));
 sky130_fd_sc_hd__nand2_1 _33456_ (.A(_12510_),
    .B(net850),
    .Y(_12511_));
 sky130_fd_sc_hd__nand2_1 _33457_ (.A(_12506_),
    .B(_12511_),
    .Y(_12512_));
 sky130_fd_sc_hd__nand2_1 _33458_ (.A(net677),
    .B(_12512_),
    .Y(_12513_));
 sky130_fd_sc_hd__nand2_1 _33459_ (.A(net635),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[27] ),
    .Y(_12514_));
 sky130_fd_sc_hd__a21oi_4 _33460_ (.A1(_12513_),
    .A2(_12514_),
    .B1(net2945),
    .Y(_04139_));
 sky130_fd_sc_hd__inv_1 _33461_ (.A(_12490_),
    .Y(_12515_));
 sky130_fd_sc_hd__nand4_1 _33462_ (.A(_12395_),
    .B(\inst$top.soc.cpu.sink__payload[26] ),
    .C(\inst$top.soc.cpu.sink__payload[29] ),
    .D(_12515_),
    .Y(_12516_));
 sky130_fd_sc_hd__xnor2_1 _33463_ (.A(\inst$top.soc.cpu.sink__payload[30] ),
    .B(_12516_),
    .Y(_12517_));
 sky130_fd_sc_hd__inv_1 _33464_ (.A(_12517_),
    .Y(_12518_));
 sky130_fd_sc_hd__nand2_1 _33465_ (.A(net742),
    .B(_12518_),
    .Y(_12519_));
 sky130_fd_sc_hd__nand2_1 _33466_ (.A(_03356_),
    .B(_03358_),
    .Y(_12520_));
 sky130_fd_sc_hd__nand2_1 _33467_ (.A(_03360_),
    .B(_03362_),
    .Y(_12521_));
 sky130_fd_sc_hd__nor2_1 _33468_ (.A(_12520_),
    .B(_12521_),
    .Y(_12522_));
 sky130_fd_sc_hd__a21oi_1 _33469_ (.A1(_03362_),
    .A2(_03359_),
    .B1(_03361_),
    .Y(_12523_));
 sky130_fd_sc_hd__o21ai_0 _33470_ (.A1(_12521_),
    .A2(_12473_),
    .B1(_12523_),
    .Y(_12524_));
 sky130_fd_sc_hd__a21oi_1 _33471_ (.A1(_12413_),
    .A2(_12522_),
    .B1(_12524_),
    .Y(_12525_));
 sky130_fd_sc_hd__xor2_1 _33472_ (.A(_03364_),
    .B(_12525_),
    .X(_12526_));
 sky130_fd_sc_hd__nand3_1 _33473_ (.A(net792),
    .B(net833),
    .C(_12526_),
    .Y(_12527_));
 sky130_fd_sc_hd__nand3_1 _33474_ (.A(_12519_),
    .B(_12527_),
    .C(net817),
    .Y(_12528_));
 sky130_fd_sc_hd__nand2_1 _33475_ (.A(net838),
    .B(\inst$top.soc.cpu.sink__payload$6[30] ),
    .Y(_12529_));
 sky130_fd_sc_hd__nand2_1 _33476_ (.A(_12528_),
    .B(_12529_),
    .Y(_12530_));
 sky130_fd_sc_hd__nand2_1 _33477_ (.A(_12530_),
    .B(net870),
    .Y(_12531_));
 sky130_fd_sc_hd__nand3_1 _33478_ (.A(net1818),
    .B(\inst$top.soc.cpu.sink__payload$18[210] ),
    .C(net1839),
    .Y(_12532_));
 sky130_fd_sc_hd__o211ai_1 _33479_ (.A1(_19900_),
    .A2(net1818),
    .B1(net2542),
    .C1(_12532_),
    .Y(_12533_));
 sky130_fd_sc_hd__o211ai_1 _33480_ (.A1(net2542),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[28] ),
    .B1(_12533_),
    .C1(net877),
    .Y(_12534_));
 sky130_fd_sc_hd__o21ai_0 _33481_ (.A1(_05866_),
    .A2(net877),
    .B1(_12534_),
    .Y(_12535_));
 sky130_fd_sc_hd__nand2_1 _33482_ (.A(_12535_),
    .B(net850),
    .Y(_12536_));
 sky130_fd_sc_hd__nand2_1 _33483_ (.A(_12531_),
    .B(_12536_),
    .Y(_12537_));
 sky130_fd_sc_hd__nand2_1 _33484_ (.A(net677),
    .B(_12537_),
    .Y(_12538_));
 sky130_fd_sc_hd__nand2_1 _33485_ (.A(net635),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[28] ),
    .Y(_12539_));
 sky130_fd_sc_hd__a21oi_4 _33486_ (.A1(_12538_),
    .A2(_12539_),
    .B1(net2945),
    .Y(_04140_));
 sky130_fd_sc_hd__a21oi_1 _33487_ (.A1(_12430_),
    .A2(_12321_),
    .B1(_12323_),
    .Y(_12540_));
 sky130_fd_sc_hd__inv_1 _33488_ (.A(_03362_),
    .Y(_12541_));
 sky130_fd_sc_hd__inv_1 _33489_ (.A(_03364_),
    .Y(_12542_));
 sky130_fd_sc_hd__nor3_1 _33490_ (.A(_12541_),
    .B(_12542_),
    .C(_12496_),
    .Y(_12543_));
 sky130_fd_sc_hd__nand2_1 _33491_ (.A(_12543_),
    .B(_12434_),
    .Y(_12544_));
 sky130_fd_sc_hd__nor4_1 _33492_ (.A(_12138_),
    .B(_12191_),
    .C(_12432_),
    .D(_12544_),
    .Y(_12545_));
 sky130_fd_sc_hd__nand2_1 _33493_ (.A(_12545_),
    .B(_12089_),
    .Y(_12546_));
 sky130_fd_sc_hd__o21bai_1 _33494_ (.A1(_12541_),
    .A2(_12498_),
    .B1_N(_03361_),
    .Y(_12547_));
 sky130_fd_sc_hd__a221oi_1 _33495_ (.A1(_12547_),
    .A2(_03364_),
    .B1(_12439_),
    .B2(_12543_),
    .C1(_03363_),
    .Y(_12548_));
 sky130_fd_sc_hd__o211ai_1 _33496_ (.A1(_12540_),
    .A2(_12544_),
    .B1(_12546_),
    .C1(_12548_),
    .Y(_12549_));
 sky130_fd_sc_hd__xnor2_1 _33497_ (.A(\inst$top.soc.cpu.sink__payload$6[31] ),
    .B(_11911_),
    .Y(_12550_));
 sky130_fd_sc_hd__xor2_2 _33498_ (.A(_12549_),
    .B(_12550_),
    .X(_12551_));
 sky130_fd_sc_hd__nand3b_1 _33499_ (.A_N(_12551_),
    .B(net790),
    .C(net831),
    .Y(_12552_));
 sky130_fd_sc_hd__nand4_1 _33500_ (.A(_12450_),
    .B(\inst$top.soc.cpu.sink__payload[29] ),
    .C(\inst$top.soc.cpu.sink__payload[30] ),
    .D(_12515_),
    .Y(_12553_));
 sky130_fd_sc_hd__xnor2_1 _33501_ (.A(\inst$top.soc.cpu.sink__payload[31] ),
    .B(_12553_),
    .Y(_12554_));
 sky130_fd_sc_hd__inv_1 _33502_ (.A(_12554_),
    .Y(_12555_));
 sky130_fd_sc_hd__nand2_1 _33503_ (.A(net740),
    .B(_12555_),
    .Y(_12556_));
 sky130_fd_sc_hd__nand3_1 _33504_ (.A(_12552_),
    .B(_12556_),
    .C(net813),
    .Y(_12557_));
 sky130_fd_sc_hd__nand2_1 _33505_ (.A(net837),
    .B(\inst$top.soc.cpu.sink__payload$6[31] ),
    .Y(_12558_));
 sky130_fd_sc_hd__nand2_1 _33506_ (.A(_12557_),
    .B(_12558_),
    .Y(_12559_));
 sky130_fd_sc_hd__nand2_1 _33507_ (.A(_12559_),
    .B(net870),
    .Y(_12560_));
 sky130_fd_sc_hd__nand3_1 _33508_ (.A(net1816),
    .B(\inst$top.soc.cpu.sink__payload$18[211] ),
    .C(net1838),
    .Y(_12561_));
 sky130_fd_sc_hd__o211ai_1 _33509_ (.A1(_19869_),
    .A2(net1816),
    .B1(net2537),
    .C1(_12561_),
    .Y(_12562_));
 sky130_fd_sc_hd__o211ai_1 _33510_ (.A1(net2537),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[29] ),
    .B1(_12562_),
    .C1(net872),
    .Y(_12563_));
 sky130_fd_sc_hd__o21ai_0 _33511_ (.A1(_05880_),
    .A2(net872),
    .B1(_12563_),
    .Y(_12564_));
 sky130_fd_sc_hd__nand2_1 _33512_ (.A(_12564_),
    .B(net848),
    .Y(_12565_));
 sky130_fd_sc_hd__nand2_1 _33513_ (.A(_12560_),
    .B(_12565_),
    .Y(_12566_));
 sky130_fd_sc_hd__nand2_1 _33514_ (.A(net674),
    .B(_12566_),
    .Y(_12567_));
 sky130_fd_sc_hd__nand2_1 _33516_ (.A(net621),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[29] ),
    .Y(_12569_));
 sky130_fd_sc_hd__a21oi_4 _33517_ (.A1(_12567_),
    .A2(_12569_),
    .B1(net2935),
    .Y(_04141_));
 sky130_fd_sc_hd__nand2_1 _33518_ (.A(net621),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[2] ),
    .Y(_12570_));
 sky130_fd_sc_hd__xor2_1 _33519_ (.A(_02866_),
    .B(\inst$top.soc.cpu.sink__payload[4] ),
    .X(_12571_));
 sky130_fd_sc_hd__nand2_1 _33520_ (.A(net740),
    .B(_12571_),
    .Y(_12572_));
 sky130_fd_sc_hd__xor2_1 _33521_ (.A(_02546_),
    .B(_03312_),
    .X(_12573_));
 sky130_fd_sc_hd__nand3_1 _33522_ (.A(net790),
    .B(net831),
    .C(_12573_),
    .Y(_12574_));
 sky130_fd_sc_hd__nand3_1 _33523_ (.A(_12572_),
    .B(_12574_),
    .C(net813),
    .Y(_12575_));
 sky130_fd_sc_hd__nor2_1 _33524_ (.A(\inst$top.soc.cpu.sink__payload$6[4] ),
    .B(net813),
    .Y(_12576_));
 sky130_fd_sc_hd__nor2_1 _33525_ (.A(net846),
    .B(_12576_),
    .Y(_12577_));
 sky130_fd_sc_hd__nand2_1 _33526_ (.A(_12575_),
    .B(_12577_),
    .Y(_12578_));
 sky130_fd_sc_hd__nand2_1 _33527_ (.A(\inst$top.soc.cpu.sink__payload$12[4] ),
    .B(_02862_),
    .Y(_12579_));
 sky130_fd_sc_hd__o311ai_0 _33528_ (.A1(_02862_),
    .A2(_11865_),
    .A3(_20257_),
    .B1(net2537),
    .C1(_12579_),
    .Y(_12580_));
 sky130_fd_sc_hd__o211ai_1 _33529_ (.A1(net2537),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[2] ),
    .B1(_12580_),
    .C1(net872),
    .Y(_12581_));
 sky130_fd_sc_hd__o21ai_0 _33530_ (.A1(_20548_),
    .A2(net872),
    .B1(_12581_),
    .Y(_12582_));
 sky130_fd_sc_hd__nand2_1 _33531_ (.A(_12582_),
    .B(net846),
    .Y(_12583_));
 sky130_fd_sc_hd__nand2_1 _33532_ (.A(_12578_),
    .B(_12583_),
    .Y(_12584_));
 sky130_fd_sc_hd__nand3_1 _33533_ (.A(_12584_),
    .B(net663),
    .C(net753),
    .Y(_12585_));
 sky130_fd_sc_hd__a21oi_4 _33534_ (.A1(_12570_),
    .A2(_12585_),
    .B1(net2935),
    .Y(_04142_));
 sky130_fd_sc_hd__xor2_1 _33535_ (.A(\inst$top.soc.cpu.sink__payload[5] ),
    .B(_12005_),
    .X(_12586_));
 sky130_fd_sc_hd__nand2_1 _33536_ (.A(net740),
    .B(_12586_),
    .Y(_12587_));
 sky130_fd_sc_hd__xnor2_1 _33537_ (.A(_03314_),
    .B(_12015_),
    .Y(_12588_));
 sky130_fd_sc_hd__nand3_1 _33538_ (.A(net790),
    .B(net831),
    .C(_12588_),
    .Y(_12589_));
 sky130_fd_sc_hd__nand3_1 _33539_ (.A(_12587_),
    .B(_12589_),
    .C(net815),
    .Y(_12590_));
 sky130_fd_sc_hd__a21oi_1 _33540_ (.A1(net837),
    .A2(\inst$top.soc.cpu.sink__payload$6[5] ),
    .B1(net847),
    .Y(_12591_));
 sky130_fd_sc_hd__nand3_1 _33541_ (.A(net1815),
    .B(\inst$top.soc.cpu.sink__payload$18[185] ),
    .C(net1838),
    .Y(_12592_));
 sky130_fd_sc_hd__o211ai_1 _33542_ (.A1(_20566_),
    .A2(net1815),
    .B1(net2539),
    .C1(_12592_),
    .Y(_12593_));
 sky130_fd_sc_hd__o211ai_1 _33543_ (.A1(net2539),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[3] ),
    .B1(_12593_),
    .C1(net874),
    .Y(_12594_));
 sky130_fd_sc_hd__o21ai_0 _33544_ (.A1(_20575_),
    .A2(net874),
    .B1(_12594_),
    .Y(_12595_));
 sky130_fd_sc_hd__nor2_1 _33545_ (.A(net870),
    .B(_12595_),
    .Y(_12596_));
 sky130_fd_sc_hd__a21oi_1 _33546_ (.A1(_12590_),
    .A2(_12591_),
    .B1(_12596_),
    .Y(_12597_));
 sky130_fd_sc_hd__nand2_1 _33547_ (.A(net668),
    .B(_12597_),
    .Y(_12598_));
 sky130_fd_sc_hd__nand2_1 _33548_ (.A(net622),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[3] ),
    .Y(_12599_));
 sky130_fd_sc_hd__a21oi_4 _33549_ (.A1(_12598_),
    .A2(_12599_),
    .B1(net2934),
    .Y(_04143_));
 sky130_fd_sc_hd__xor2_1 _33550_ (.A(\inst$top.soc.cpu.sink__payload[6] ),
    .B(_11959_),
    .X(_12600_));
 sky130_fd_sc_hd__nand2_1 _33551_ (.A(net740),
    .B(_12600_),
    .Y(_12601_));
 sky130_fd_sc_hd__xnor2_1 _33552_ (.A(_03316_),
    .B(_11977_),
    .Y(_12602_));
 sky130_fd_sc_hd__nand3_1 _33553_ (.A(net790),
    .B(net831),
    .C(_12602_),
    .Y(_12603_));
 sky130_fd_sc_hd__nand3_1 _33554_ (.A(_12601_),
    .B(_12603_),
    .C(net815),
    .Y(_12604_));
 sky130_fd_sc_hd__a21oi_1 _33555_ (.A1(net837),
    .A2(\inst$top.soc.cpu.sink__payload$6[6] ),
    .B1(net846),
    .Y(_12605_));
 sky130_fd_sc_hd__nand3_1 _33556_ (.A(net1815),
    .B(\inst$top.soc.cpu.sink__payload$18[186] ),
    .C(net1838),
    .Y(_12606_));
 sky130_fd_sc_hd__o211ai_1 _33557_ (.A1(_20594_),
    .A2(net1815),
    .B1(net2539),
    .C1(_12606_),
    .Y(_12607_));
 sky130_fd_sc_hd__o211ai_1 _33558_ (.A1(net2539),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[4] ),
    .B1(_12607_),
    .C1(net874),
    .Y(_12608_));
 sky130_fd_sc_hd__o21ai_0 _33559_ (.A1(_20603_),
    .A2(net874),
    .B1(_12608_),
    .Y(_12609_));
 sky130_fd_sc_hd__nor2_1 _33560_ (.A(net870),
    .B(_12609_),
    .Y(_12610_));
 sky130_fd_sc_hd__a21oi_1 _33561_ (.A1(_12604_),
    .A2(_12605_),
    .B1(_12610_),
    .Y(_12611_));
 sky130_fd_sc_hd__nand2_1 _33562_ (.A(net668),
    .B(_12611_),
    .Y(_12612_));
 sky130_fd_sc_hd__nand2_1 _33563_ (.A(net621),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[4] ),
    .Y(_12613_));
 sky130_fd_sc_hd__a21oi_4 _33564_ (.A1(_12612_),
    .A2(_12613_),
    .B1(net2934),
    .Y(_04144_));
 sky130_fd_sc_hd__xor2_1 _33565_ (.A(\inst$top.soc.cpu.sink__payload[7] ),
    .B(_12007_),
    .X(_12614_));
 sky130_fd_sc_hd__nand2_1 _33566_ (.A(net740),
    .B(_12614_),
    .Y(_12615_));
 sky130_fd_sc_hd__xnor2_1 _33567_ (.A(_03318_),
    .B(_12086_),
    .Y(_12616_));
 sky130_fd_sc_hd__nand3_1 _33568_ (.A(net790),
    .B(net831),
    .C(_12616_),
    .Y(_12617_));
 sky130_fd_sc_hd__nand3_1 _33569_ (.A(_12615_),
    .B(_12617_),
    .C(net813),
    .Y(_12618_));
 sky130_fd_sc_hd__a21oi_1 _33570_ (.A1(net837),
    .A2(\inst$top.soc.cpu.sink__payload$6[7] ),
    .B1(net846),
    .Y(_12619_));
 sky130_fd_sc_hd__nand3_1 _33571_ (.A(net1816),
    .B(\inst$top.soc.cpu.sink__payload$18[187] ),
    .C(net1838),
    .Y(_12620_));
 sky130_fd_sc_hd__o211ai_1 _33572_ (.A1(_20623_),
    .A2(net1816),
    .B1(net2537),
    .C1(_12620_),
    .Y(_12621_));
 sky130_fd_sc_hd__o211ai_1 _33573_ (.A1(net2540),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[5] ),
    .B1(_12621_),
    .C1(net875),
    .Y(_12622_));
 sky130_fd_sc_hd__o21ai_0 _33574_ (.A1(_11557_),
    .A2(net872),
    .B1(_12622_),
    .Y(_12623_));
 sky130_fd_sc_hd__nor2_1 _33575_ (.A(net870),
    .B(_12623_),
    .Y(_12624_));
 sky130_fd_sc_hd__a21oi_1 _33576_ (.A1(_12618_),
    .A2(_12619_),
    .B1(_12624_),
    .Y(_12625_));
 sky130_fd_sc_hd__nand2_1 _33577_ (.A(net668),
    .B(_12625_),
    .Y(_12626_));
 sky130_fd_sc_hd__nand2_1 _33578_ (.A(net621),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[5] ),
    .Y(_12627_));
 sky130_fd_sc_hd__a21oi_4 _33579_ (.A1(_12626_),
    .A2(_12627_),
    .B1(net2943),
    .Y(_04145_));
 sky130_fd_sc_hd__xnor2_1 _33580_ (.A(\inst$top.soc.cpu.sink__payload[8] ),
    .B(_11960_),
    .Y(_12628_));
 sky130_fd_sc_hd__nand2_1 _33581_ (.A(net742),
    .B(_12628_),
    .Y(_12629_));
 sky130_fd_sc_hd__a21oi_1 _33582_ (.A1(_02546_),
    .A2(_12224_),
    .B1(_12231_),
    .Y(_12630_));
 sky130_fd_sc_hd__xor2_1 _33583_ (.A(_03320_),
    .B(_12630_),
    .X(_12631_));
 sky130_fd_sc_hd__nand3_1 _33584_ (.A(net790),
    .B(net832),
    .C(_12631_),
    .Y(_12632_));
 sky130_fd_sc_hd__nand3_1 _33585_ (.A(_12629_),
    .B(_12632_),
    .C(net814),
    .Y(_12633_));
 sky130_fd_sc_hd__a21oi_1 _33586_ (.A1(net837),
    .A2(\inst$top.soc.cpu.sink__payload$6[8] ),
    .B1(net850),
    .Y(_12634_));
 sky130_fd_sc_hd__nand3_1 _33587_ (.A(net1817),
    .B(\inst$top.soc.cpu.sink__payload$18[188] ),
    .C(net1840),
    .Y(_12635_));
 sky130_fd_sc_hd__o211ai_1 _33588_ (.A1(_20664_),
    .A2(net1817),
    .B1(net2541),
    .C1(_12635_),
    .Y(_12636_));
 sky130_fd_sc_hd__o211ai_1 _33589_ (.A1(net2541),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[6] ),
    .B1(_12636_),
    .C1(net876),
    .Y(_12637_));
 sky130_fd_sc_hd__o21ai_0 _33590_ (.A1(_20672_),
    .A2(net876),
    .B1(_12637_),
    .Y(_12638_));
 sky130_fd_sc_hd__nor2_1 _33591_ (.A(net870),
    .B(_12638_),
    .Y(_12639_));
 sky130_fd_sc_hd__a21oi_1 _33592_ (.A1(_12633_),
    .A2(_12634_),
    .B1(_12639_),
    .Y(_12640_));
 sky130_fd_sc_hd__nand2_1 _33593_ (.A(net675),
    .B(_12640_),
    .Y(_12641_));
 sky130_fd_sc_hd__nand2_1 _33594_ (.A(net626),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[6] ),
    .Y(_12642_));
 sky130_fd_sc_hd__a21oi_4 _33595_ (.A1(_12641_),
    .A2(_12642_),
    .B1(net2932),
    .Y(_04146_));
 sky130_fd_sc_hd__xor2_1 _33596_ (.A(\inst$top.soc.cpu.sink__payload[9] ),
    .B(_12008_),
    .X(_12643_));
 sky130_fd_sc_hd__nand2_1 _33597_ (.A(net740),
    .B(_12643_),
    .Y(_12644_));
 sky130_fd_sc_hd__xnor2_1 _33598_ (.A(_03322_),
    .B(_12024_),
    .Y(_12645_));
 sky130_fd_sc_hd__nand3_1 _33599_ (.A(net790),
    .B(net832),
    .C(_12645_),
    .Y(_12646_));
 sky130_fd_sc_hd__nand3_1 _33600_ (.A(_12644_),
    .B(_12646_),
    .C(net814),
    .Y(_12647_));
 sky130_fd_sc_hd__a21oi_1 _33601_ (.A1(net837),
    .A2(\inst$top.soc.cpu.sink__payload$6[9] ),
    .B1(net850),
    .Y(_12648_));
 sky130_fd_sc_hd__nand3_1 _33602_ (.A(net1817),
    .B(\inst$top.soc.cpu.sink__payload$18[189] ),
    .C(net1840),
    .Y(_12649_));
 sky130_fd_sc_hd__o211ai_1 _33603_ (.A1(_20685_),
    .A2(net1817),
    .B1(net2541),
    .C1(_12649_),
    .Y(_12650_));
 sky130_fd_sc_hd__o211ai_1 _33604_ (.A1(net2541),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[7] ),
    .B1(_12650_),
    .C1(net876),
    .Y(_12651_));
 sky130_fd_sc_hd__o21ai_0 _33605_ (.A1(_11560_),
    .A2(net876),
    .B1(_12651_),
    .Y(_12652_));
 sky130_fd_sc_hd__nor2_1 _33606_ (.A(net870),
    .B(_12652_),
    .Y(_12653_));
 sky130_fd_sc_hd__a21oi_1 _33607_ (.A1(_12647_),
    .A2(_12648_),
    .B1(_12653_),
    .Y(_12654_));
 sky130_fd_sc_hd__nand2_1 _33608_ (.A(net675),
    .B(_12654_),
    .Y(_12655_));
 sky130_fd_sc_hd__nand2_1 _33609_ (.A(net626),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[7] ),
    .Y(_12656_));
 sky130_fd_sc_hd__a21oi_4 _33611_ (.A1(_12655_),
    .A2(_12656_),
    .B1(net2933),
    .Y(_04147_));
 sky130_fd_sc_hd__nand2_1 _33612_ (.A(net627),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[8] ),
    .Y(_12658_));
 sky130_fd_sc_hd__xor2_1 _33613_ (.A(_11956_),
    .B(_11961_),
    .X(_12659_));
 sky130_fd_sc_hd__nand2_1 _33614_ (.A(net742),
    .B(_12659_),
    .Y(_12660_));
 sky130_fd_sc_hd__xor2_1 _33615_ (.A(_03324_),
    .B(_11981_),
    .X(_12661_));
 sky130_fd_sc_hd__nand3_1 _33616_ (.A(net792),
    .B(net833),
    .C(_12661_),
    .Y(_12662_));
 sky130_fd_sc_hd__nand3_1 _33617_ (.A(_12660_),
    .B(_12662_),
    .C(net816),
    .Y(_12663_));
 sky130_fd_sc_hd__nor2_1 _33618_ (.A(\inst$top.soc.cpu.sink__payload$6[10] ),
    .B(net816),
    .Y(_12664_));
 sky130_fd_sc_hd__nor2_1 _33619_ (.A(net849),
    .B(_12664_),
    .Y(_12665_));
 sky130_fd_sc_hd__nand2_1 _33620_ (.A(_12663_),
    .B(_12665_),
    .Y(_12666_));
 sky130_fd_sc_hd__nand3_1 _33621_ (.A(net1820),
    .B(\inst$top.soc.cpu.sink__payload$18[190] ),
    .C(net1839),
    .Y(_12667_));
 sky130_fd_sc_hd__o211ai_1 _33622_ (.A1(_20705_),
    .A2(net1820),
    .B1(net2544),
    .C1(_12667_),
    .Y(_12668_));
 sky130_fd_sc_hd__o211ai_1 _33623_ (.A1(net2543),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[8] ),
    .B1(_12668_),
    .C1(net878),
    .Y(_12669_));
 sky130_fd_sc_hd__o21ai_0 _33624_ (.A1(_20714_),
    .A2(net876),
    .B1(_12669_),
    .Y(_12670_));
 sky130_fd_sc_hd__nand2_1 _33625_ (.A(_12670_),
    .B(net849),
    .Y(_12671_));
 sky130_fd_sc_hd__nand2_1 _33626_ (.A(_12666_),
    .B(_12671_),
    .Y(_12672_));
 sky130_fd_sc_hd__nand3_1 _33627_ (.A(_12672_),
    .B(net663),
    .C(net753),
    .Y(_12673_));
 sky130_fd_sc_hd__a21oi_4 _33628_ (.A1(_12658_),
    .A2(_12673_),
    .B1(net2933),
    .Y(_04148_));
 sky130_fd_sc_hd__nand2_1 _33629_ (.A(net621),
    .B(\inst$top.soc.cpu.fetch.ibus__adr[9] ),
    .Y(_12674_));
 sky130_fd_sc_hd__xor2_1 _33630_ (.A(\inst$top.soc.cpu.sink__payload[11] ),
    .B(_12067_),
    .X(_12675_));
 sky130_fd_sc_hd__nand2_1 _33631_ (.A(net740),
    .B(_12675_),
    .Y(_12676_));
 sky130_fd_sc_hd__xor2_1 _33632_ (.A(_03326_),
    .B(_12027_),
    .X(_12677_));
 sky130_fd_sc_hd__nand3_1 _33633_ (.A(net791),
    .B(net832),
    .C(_12677_),
    .Y(_12678_));
 sky130_fd_sc_hd__nand3_1 _33634_ (.A(_12676_),
    .B(_12678_),
    .C(net814),
    .Y(_12679_));
 sky130_fd_sc_hd__nor2_1 _33635_ (.A(\inst$top.soc.cpu.sink__payload$6[11] ),
    .B(net814),
    .Y(_12680_));
 sky130_fd_sc_hd__nor2_1 _33636_ (.A(net847),
    .B(_12680_),
    .Y(_12681_));
 sky130_fd_sc_hd__nand2_1 _33637_ (.A(_12679_),
    .B(_12681_),
    .Y(_12682_));
 sky130_fd_sc_hd__nand3_1 _33638_ (.A(net1815),
    .B(\inst$top.soc.cpu.sink__payload$18[191] ),
    .C(net1838),
    .Y(_12683_));
 sky130_fd_sc_hd__o211ai_1 _33639_ (.A1(_20726_),
    .A2(net1815),
    .B1(net2538),
    .C1(_12683_),
    .Y(_12684_));
 sky130_fd_sc_hd__o211ai_1 _33640_ (.A1(net2538),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[9] ),
    .B1(_12684_),
    .C1(net873),
    .Y(_12685_));
 sky130_fd_sc_hd__o21ai_0 _33641_ (.A1(_20737_),
    .A2(net873),
    .B1(_12685_),
    .Y(_12686_));
 sky130_fd_sc_hd__nand2_1 _33642_ (.A(_12686_),
    .B(net847),
    .Y(_12687_));
 sky130_fd_sc_hd__nand2_1 _33643_ (.A(_12682_),
    .B(_12687_),
    .Y(_12688_));
 sky130_fd_sc_hd__nand3_1 _33644_ (.A(_12688_),
    .B(net663),
    .C(net753),
    .Y(_12689_));
 sky130_fd_sc_hd__a21oi_4 _33645_ (.A1(_12674_),
    .A2(_12689_),
    .B1(net2934),
    .Y(_04149_));
 sky130_fd_sc_hd__nor2_1 _33647_ (.A(\inst$top.soc.sram.wb_bus__ack ),
    .B(\inst$top.soc.wb_to_csr.wb_bus__ack ),
    .Y(_12691_));
 sky130_fd_sc_hd__inv_1 _33648_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__ack ),
    .Y(_12692_));
 sky130_fd_sc_hd__nand2_1 _33649_ (.A(_12691_),
    .B(_12692_),
    .Y(_12693_));
 sky130_fd_sc_hd__nand2_1 _33650_ (.A(_12693_),
    .B(_19847_),
    .Y(_12694_));
 sky130_fd_sc_hd__nand2_1 _33651_ (.A(_12694_),
    .B(\inst$top.soc.cpu.fetch.ibus__cyc ),
    .Y(_12695_));
 sky130_fd_sc_hd__a21oi_2 _33652_ (.A1(net639),
    .A2(_12695_),
    .B1(net2949),
    .Y(_04150_));
 sky130_fd_sc_hd__nand2_1 _33653_ (.A(_12693_),
    .B(_09341_),
    .Y(_12696_));
 sky130_fd_sc_hd__nand2_1 _33655_ (.A(net1802),
    .B(\inst$top.soc.cpu.fetch.ibus__stb ),
    .Y(_12698_));
 sky130_fd_sc_hd__a21oi_2 _33656_ (.A1(net639),
    .A2(_12698_),
    .B1(net2951),
    .Y(_04151_));
 sky130_fd_sc_hd__inv_1 _33658_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[0] ),
    .Y(_12700_));
 sky130_fd_sc_hd__inv_1 _33659_ (.A(_09280_),
    .Y(_12701_));
 sky130_fd_sc_hd__nor2_1 _33660_ (.A(_09311_),
    .B(_12701_),
    .Y(_12702_));
 sky130_fd_sc_hd__nand3_1 _33661_ (.A(_12702_),
    .B(_09308_),
    .C(_09304_),
    .Y(_12703_));
 sky130_fd_sc_hd__nor3_1 _33663_ (.A(_09304_),
    .B(_09280_),
    .C(_09277_),
    .Y(_12705_));
 sky130_fd_sc_hd__nor2_1 _33664_ (.A(_09311_),
    .B(_09308_),
    .Y(_12706_));
 sky130_fd_sc_hd__and2_1 _33665_ (.A(_12705_),
    .B(_12706_),
    .X(_12707_));
 sky130_fd_sc_hd__nand2_1 _33668_ (.A(net1082),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[0] ),
    .Y(_12710_));
 sky130_fd_sc_hd__nand2_1 _33670_ (.A(net858),
    .B(\inst$top.soc.sram.read_port__data[0] ),
    .Y(_12712_));
 sky130_fd_sc_hd__o211ai_1 _33671_ (.A1(_12700_),
    .A2(net1084),
    .B1(_12710_),
    .C1(_12712_),
    .Y(_12713_));
 sky130_fd_sc_hd__inv_1 _33673_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[0] ),
    .Y(_12715_));
 sky130_fd_sc_hd__a21oi_1 _33674_ (.A1(net1799),
    .A2(_12715_),
    .B1(net2948),
    .Y(_12716_));
 sky130_fd_sc_hd__o21ai_0 _33675_ (.A1(net1800),
    .A2(_12713_),
    .B1(_12716_),
    .Y(_12717_));
 sky130_fd_sc_hd__inv_2 _33676_ (.A(_12717_),
    .Y(_04152_));
 sky130_fd_sc_hd__inv_1 _33677_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[10] ),
    .Y(_12718_));
 sky130_fd_sc_hd__inv_1 _33679_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[10] ),
    .Y(_12720_));
 sky130_fd_sc_hd__clkinv_1 _33680_ (.A(net1082),
    .Y(_12721_));
 sky130_fd_sc_hd__nand2_1 _33683_ (.A(net859),
    .B(\inst$top.soc.sram.read_port__data[10] ),
    .Y(_12724_));
 sky130_fd_sc_hd__o221ai_1 _33684_ (.A1(_12718_),
    .A2(net1086),
    .B1(_12720_),
    .B2(net1026),
    .C1(_12724_),
    .Y(_12725_));
 sky130_fd_sc_hd__inv_1 _33685_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[10] ),
    .Y(_12726_));
 sky130_fd_sc_hd__a21oi_1 _33686_ (.A1(net1803),
    .A2(_12726_),
    .B1(net2980),
    .Y(_12727_));
 sky130_fd_sc_hd__o21ai_0 _33687_ (.A1(net1803),
    .A2(_12725_),
    .B1(_12727_),
    .Y(_12728_));
 sky130_fd_sc_hd__inv_2 _33688_ (.A(_12728_),
    .Y(_04153_));
 sky130_fd_sc_hd__inv_1 _33689_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[11] ),
    .Y(_12729_));
 sky130_fd_sc_hd__inv_1 _33690_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[11] ),
    .Y(_12730_));
 sky130_fd_sc_hd__nand2_1 _33691_ (.A(net861),
    .B(\inst$top.soc.sram.read_port__data[11] ),
    .Y(_12731_));
 sky130_fd_sc_hd__o221ai_1 _33692_ (.A1(_12729_),
    .A2(net1085),
    .B1(_12730_),
    .B2(net1025),
    .C1(_12731_),
    .Y(_12732_));
 sky130_fd_sc_hd__inv_1 _33693_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[11] ),
    .Y(_12733_));
 sky130_fd_sc_hd__a21oi_1 _33694_ (.A1(net1804),
    .A2(_12733_),
    .B1(net2980),
    .Y(_12734_));
 sky130_fd_sc_hd__o21ai_0 _33695_ (.A1(net1804),
    .A2(_12732_),
    .B1(_12734_),
    .Y(_12735_));
 sky130_fd_sc_hd__inv_2 _33696_ (.A(_12735_),
    .Y(_04154_));
 sky130_fd_sc_hd__inv_1 _33697_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[12] ),
    .Y(_12736_));
 sky130_fd_sc_hd__nand2_1 _33698_ (.A(net1083),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[12] ),
    .Y(_12737_));
 sky130_fd_sc_hd__nand2_1 _33699_ (.A(net860),
    .B(\inst$top.soc.sram.read_port__data[12] ),
    .Y(_12738_));
 sky130_fd_sc_hd__o211ai_1 _33700_ (.A1(_12736_),
    .A2(net1085),
    .B1(_12737_),
    .C1(_12738_),
    .Y(_12739_));
 sky130_fd_sc_hd__inv_1 _33701_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[12] ),
    .Y(_12740_));
 sky130_fd_sc_hd__a21oi_1 _33702_ (.A1(net1803),
    .A2(_12740_),
    .B1(net2982),
    .Y(_12741_));
 sky130_fd_sc_hd__o21ai_0 _33703_ (.A1(net1803),
    .A2(_12739_),
    .B1(_12741_),
    .Y(_12742_));
 sky130_fd_sc_hd__inv_2 _33704_ (.A(_12742_),
    .Y(_04155_));
 sky130_fd_sc_hd__inv_1 _33705_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[13] ),
    .Y(_12743_));
 sky130_fd_sc_hd__nand2_1 _33706_ (.A(net1083),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[13] ),
    .Y(_12744_));
 sky130_fd_sc_hd__nand2_1 _33707_ (.A(net859),
    .B(\inst$top.soc.sram.read_port__data[13] ),
    .Y(_12745_));
 sky130_fd_sc_hd__o211ai_1 _33708_ (.A1(_12743_),
    .A2(net1086),
    .B1(_12744_),
    .C1(_12745_),
    .Y(_12746_));
 sky130_fd_sc_hd__inv_1 _33709_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[13] ),
    .Y(_12747_));
 sky130_fd_sc_hd__a21oi_1 _33710_ (.A1(net1803),
    .A2(_12747_),
    .B1(net2982),
    .Y(_12748_));
 sky130_fd_sc_hd__o21ai_0 _33711_ (.A1(net1803),
    .A2(_12746_),
    .B1(_12748_),
    .Y(_12749_));
 sky130_fd_sc_hd__inv_2 _33712_ (.A(_12749_),
    .Y(_04156_));
 sky130_fd_sc_hd__inv_1 _33713_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[14] ),
    .Y(_12750_));
 sky130_fd_sc_hd__inv_1 _33714_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[14] ),
    .Y(_12751_));
 sky130_fd_sc_hd__nand2_1 _33715_ (.A(net860),
    .B(\inst$top.soc.sram.read_port__data[14] ),
    .Y(_12752_));
 sky130_fd_sc_hd__o221ai_2 _33716_ (.A1(_12750_),
    .A2(net1085),
    .B1(_12751_),
    .B2(net1025),
    .C1(_12752_),
    .Y(_12753_));
 sky130_fd_sc_hd__inv_1 _33717_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[14] ),
    .Y(_12754_));
 sky130_fd_sc_hd__a21oi_1 _33719_ (.A1(net1801),
    .A2(_12754_),
    .B1(net2949),
    .Y(_12756_));
 sky130_fd_sc_hd__o21ai_0 _33720_ (.A1(net1801),
    .A2(_12753_),
    .B1(_12756_),
    .Y(_12757_));
 sky130_fd_sc_hd__inv_2 _33721_ (.A(_12757_),
    .Y(_04157_));
 sky130_fd_sc_hd__inv_1 _33722_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[15] ),
    .Y(_12758_));
 sky130_fd_sc_hd__inv_1 _33723_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[15] ),
    .Y(_12759_));
 sky130_fd_sc_hd__nand2_1 _33724_ (.A(net860),
    .B(\inst$top.soc.sram.read_port__data[15] ),
    .Y(_12760_));
 sky130_fd_sc_hd__o221ai_1 _33725_ (.A1(_12758_),
    .A2(net1085),
    .B1(_12759_),
    .B2(net1025),
    .C1(_12760_),
    .Y(_12761_));
 sky130_fd_sc_hd__inv_1 _33726_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[15] ),
    .Y(_12762_));
 sky130_fd_sc_hd__a21oi_1 _33727_ (.A1(net1805),
    .A2(_12762_),
    .B1(net2988),
    .Y(_12763_));
 sky130_fd_sc_hd__o21ai_0 _33728_ (.A1(net1805),
    .A2(_12761_),
    .B1(_12763_),
    .Y(_12764_));
 sky130_fd_sc_hd__inv_2 _33729_ (.A(_12764_),
    .Y(_04158_));
 sky130_fd_sc_hd__inv_1 _33730_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[16] ),
    .Y(_12765_));
 sky130_fd_sc_hd__inv_1 _33731_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[16] ),
    .Y(_12766_));
 sky130_fd_sc_hd__nand2_1 _33732_ (.A(net860),
    .B(\inst$top.soc.sram.read_port__data[16] ),
    .Y(_12767_));
 sky130_fd_sc_hd__o221ai_2 _33733_ (.A1(_12765_),
    .A2(net1086),
    .B1(_12766_),
    .B2(net1026),
    .C1(_12767_),
    .Y(_12768_));
 sky130_fd_sc_hd__inv_1 _33734_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[16] ),
    .Y(_12769_));
 sky130_fd_sc_hd__a21oi_1 _33735_ (.A1(net1806),
    .A2(_12769_),
    .B1(net2989),
    .Y(_12770_));
 sky130_fd_sc_hd__o21ai_0 _33736_ (.A1(net1806),
    .A2(_12768_),
    .B1(_12770_),
    .Y(_12771_));
 sky130_fd_sc_hd__inv_2 _33737_ (.A(_12771_),
    .Y(_04159_));
 sky130_fd_sc_hd__inv_1 _33738_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[17] ),
    .Y(_12772_));
 sky130_fd_sc_hd__inv_1 _33739_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[17] ),
    .Y(_12773_));
 sky130_fd_sc_hd__nand2_1 _33740_ (.A(net860),
    .B(\inst$top.soc.sram.read_port__data[17] ),
    .Y(_12774_));
 sky130_fd_sc_hd__o221ai_2 _33741_ (.A1(_12772_),
    .A2(net1086),
    .B1(_12773_),
    .B2(net1026),
    .C1(_12774_),
    .Y(_12775_));
 sky130_fd_sc_hd__inv_1 _33743_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[17] ),
    .Y(_12777_));
 sky130_fd_sc_hd__a21oi_1 _33744_ (.A1(net1806),
    .A2(_12777_),
    .B1(net2989),
    .Y(_12778_));
 sky130_fd_sc_hd__o21ai_0 _33745_ (.A1(net1806),
    .A2(_12775_),
    .B1(_12778_),
    .Y(_12779_));
 sky130_fd_sc_hd__inv_2 _33746_ (.A(_12779_),
    .Y(_04160_));
 sky130_fd_sc_hd__inv_1 _33747_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[18] ),
    .Y(_12780_));
 sky130_fd_sc_hd__inv_1 _33748_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[18] ),
    .Y(_12781_));
 sky130_fd_sc_hd__nand2_1 _33749_ (.A(net862),
    .B(\inst$top.soc.sram.read_port__data[18] ),
    .Y(_12782_));
 sky130_fd_sc_hd__o221ai_1 _33750_ (.A1(_12780_),
    .A2(net1086),
    .B1(_12781_),
    .B2(net1026),
    .C1(_12782_),
    .Y(_12783_));
 sky130_fd_sc_hd__inv_1 _33751_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[18] ),
    .Y(_12784_));
 sky130_fd_sc_hd__a21oi_1 _33752_ (.A1(net1805),
    .A2(_12784_),
    .B1(net2981),
    .Y(_12785_));
 sky130_fd_sc_hd__o21ai_0 _33753_ (.A1(net1804),
    .A2(_12783_),
    .B1(_12785_),
    .Y(_12786_));
 sky130_fd_sc_hd__inv_2 _33754_ (.A(_12786_),
    .Y(_04161_));
 sky130_fd_sc_hd__inv_1 _33756_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[19] ),
    .Y(_12788_));
 sky130_fd_sc_hd__inv_1 _33758_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[19] ),
    .Y(_12790_));
 sky130_fd_sc_hd__nand2_1 _33760_ (.A(net861),
    .B(\inst$top.soc.sram.read_port__data[19] ),
    .Y(_12792_));
 sky130_fd_sc_hd__o221ai_1 _33761_ (.A1(_12788_),
    .A2(net1087),
    .B1(_12790_),
    .B2(net1026),
    .C1(_12792_),
    .Y(_12793_));
 sky130_fd_sc_hd__inv_1 _33762_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[19] ),
    .Y(_12794_));
 sky130_fd_sc_hd__a21oi_1 _33763_ (.A1(net1805),
    .A2(_12794_),
    .B1(net2988),
    .Y(_12795_));
 sky130_fd_sc_hd__o21ai_0 _33764_ (.A1(net1805),
    .A2(_12793_),
    .B1(_12795_),
    .Y(_12796_));
 sky130_fd_sc_hd__inv_2 _33765_ (.A(_12796_),
    .Y(_04162_));
 sky130_fd_sc_hd__inv_1 _33766_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[1] ),
    .Y(_12797_));
 sky130_fd_sc_hd__nand2_1 _33767_ (.A(net1082),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[1] ),
    .Y(_12798_));
 sky130_fd_sc_hd__nand2_1 _33768_ (.A(net858),
    .B(\inst$top.soc.sram.read_port__data[1] ),
    .Y(_12799_));
 sky130_fd_sc_hd__o211ai_1 _33769_ (.A1(_12797_),
    .A2(net1084),
    .B1(_12798_),
    .C1(_12799_),
    .Y(_12800_));
 sky130_fd_sc_hd__inv_1 _33770_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[1] ),
    .Y(_12801_));
 sky130_fd_sc_hd__a21oi_1 _33771_ (.A1(net1799),
    .A2(_12801_),
    .B1(net2948),
    .Y(_12802_));
 sky130_fd_sc_hd__o21ai_0 _33772_ (.A1(net1799),
    .A2(_12800_),
    .B1(_12802_),
    .Y(_12803_));
 sky130_fd_sc_hd__inv_2 _33773_ (.A(_12803_),
    .Y(_04163_));
 sky130_fd_sc_hd__inv_1 _33774_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[20] ),
    .Y(_12804_));
 sky130_fd_sc_hd__inv_1 _33775_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[20] ),
    .Y(_12805_));
 sky130_fd_sc_hd__nand2_1 _33776_ (.A(net862),
    .B(\inst$top.soc.sram.read_port__data[20] ),
    .Y(_12806_));
 sky130_fd_sc_hd__o221ai_1 _33777_ (.A1(_12804_),
    .A2(net1086),
    .B1(_12805_),
    .B2(net1026),
    .C1(_12806_),
    .Y(_12807_));
 sky130_fd_sc_hd__inv_1 _33778_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[20] ),
    .Y(_12808_));
 sky130_fd_sc_hd__a21oi_1 _33779_ (.A1(net1804),
    .A2(_12808_),
    .B1(net2981),
    .Y(_12809_));
 sky130_fd_sc_hd__o21ai_0 _33780_ (.A1(net1804),
    .A2(_12807_),
    .B1(_12809_),
    .Y(_12810_));
 sky130_fd_sc_hd__inv_2 _33781_ (.A(_12810_),
    .Y(_04164_));
 sky130_fd_sc_hd__inv_1 _33782_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[21] ),
    .Y(_12811_));
 sky130_fd_sc_hd__inv_1 _33783_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[21] ),
    .Y(_12812_));
 sky130_fd_sc_hd__nand2_1 _33784_ (.A(net861),
    .B(\inst$top.soc.sram.read_port__data[21] ),
    .Y(_12813_));
 sky130_fd_sc_hd__o221ai_1 _33785_ (.A1(_12811_),
    .A2(net1086),
    .B1(_12812_),
    .B2(net1026),
    .C1(_12813_),
    .Y(_12814_));
 sky130_fd_sc_hd__inv_1 _33786_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[21] ),
    .Y(_12815_));
 sky130_fd_sc_hd__a21oi_1 _33787_ (.A1(net1805),
    .A2(_12815_),
    .B1(net2988),
    .Y(_12816_));
 sky130_fd_sc_hd__o21ai_0 _33788_ (.A1(net1805),
    .A2(_12814_),
    .B1(_12816_),
    .Y(_12817_));
 sky130_fd_sc_hd__inv_2 _33789_ (.A(_12817_),
    .Y(_04165_));
 sky130_fd_sc_hd__inv_1 _33790_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[22] ),
    .Y(_12818_));
 sky130_fd_sc_hd__inv_1 _33791_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[22] ),
    .Y(_12819_));
 sky130_fd_sc_hd__nand2_1 _33792_ (.A(net861),
    .B(\inst$top.soc.sram.read_port__data[22] ),
    .Y(_12820_));
 sky130_fd_sc_hd__o221ai_1 _33793_ (.A1(_12818_),
    .A2(net1086),
    .B1(_12819_),
    .B2(net1026),
    .C1(_12820_),
    .Y(_12821_));
 sky130_fd_sc_hd__inv_1 _33794_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[22] ),
    .Y(_12822_));
 sky130_fd_sc_hd__a21oi_1 _33795_ (.A1(net1806),
    .A2(_12822_),
    .B1(net2989),
    .Y(_12823_));
 sky130_fd_sc_hd__o21ai_0 _33796_ (.A1(net1806),
    .A2(_12821_),
    .B1(_12823_),
    .Y(_12824_));
 sky130_fd_sc_hd__inv_2 _33797_ (.A(_12824_),
    .Y(_04166_));
 sky130_fd_sc_hd__inv_1 _33798_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[23] ),
    .Y(_12825_));
 sky130_fd_sc_hd__inv_1 _33799_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[23] ),
    .Y(_12826_));
 sky130_fd_sc_hd__nand2_1 _33800_ (.A(net861),
    .B(\inst$top.soc.sram.read_port__data[23] ),
    .Y(_12827_));
 sky130_fd_sc_hd__o221ai_2 _33801_ (.A1(_12825_),
    .A2(net1086),
    .B1(_12826_),
    .B2(net1026),
    .C1(_12827_),
    .Y(_12828_));
 sky130_fd_sc_hd__inv_1 _33802_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[23] ),
    .Y(_12829_));
 sky130_fd_sc_hd__a21oi_1 _33804_ (.A1(net1803),
    .A2(_12829_),
    .B1(net2982),
    .Y(_12831_));
 sky130_fd_sc_hd__o21ai_0 _33805_ (.A1(net1803),
    .A2(_12828_),
    .B1(_12831_),
    .Y(_12832_));
 sky130_fd_sc_hd__inv_2 _33806_ (.A(_12832_),
    .Y(_04167_));
 sky130_fd_sc_hd__inv_1 _33807_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[24] ),
    .Y(_12833_));
 sky130_fd_sc_hd__nand2_1 _33808_ (.A(net1082),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[24] ),
    .Y(_12834_));
 sky130_fd_sc_hd__nand2_1 _33809_ (.A(net858),
    .B(\inst$top.soc.sram.read_port__data[24] ),
    .Y(_12835_));
 sky130_fd_sc_hd__o211ai_1 _33810_ (.A1(_12833_),
    .A2(net1084),
    .B1(_12834_),
    .C1(_12835_),
    .Y(_12836_));
 sky130_fd_sc_hd__inv_1 _33811_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[24] ),
    .Y(_12837_));
 sky130_fd_sc_hd__a21oi_1 _33812_ (.A1(net1800),
    .A2(_12837_),
    .B1(net2948),
    .Y(_12838_));
 sky130_fd_sc_hd__o21ai_0 _33813_ (.A1(net1800),
    .A2(net3038),
    .B1(_12838_),
    .Y(_12839_));
 sky130_fd_sc_hd__inv_2 _33814_ (.A(_12839_),
    .Y(_04168_));
 sky130_fd_sc_hd__inv_1 _33815_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[25] ),
    .Y(_12840_));
 sky130_fd_sc_hd__nand2_1 _33816_ (.A(net1083),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[25] ),
    .Y(_12841_));
 sky130_fd_sc_hd__nand2_1 _33817_ (.A(net858),
    .B(\inst$top.soc.sram.read_port__data[25] ),
    .Y(_12842_));
 sky130_fd_sc_hd__o211ai_1 _33818_ (.A1(_12840_),
    .A2(net1085),
    .B1(_12841_),
    .C1(_12842_),
    .Y(_12843_));
 sky130_fd_sc_hd__inv_1 _33819_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[25] ),
    .Y(_12844_));
 sky130_fd_sc_hd__a21oi_1 _33820_ (.A1(net1799),
    .A2(_12844_),
    .B1(net2949),
    .Y(_12845_));
 sky130_fd_sc_hd__o21ai_0 _33821_ (.A1(net1801),
    .A2(_12843_),
    .B1(_12845_),
    .Y(_12846_));
 sky130_fd_sc_hd__inv_2 _33822_ (.A(_12846_),
    .Y(_04169_));
 sky130_fd_sc_hd__inv_1 _33823_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[26] ),
    .Y(_12847_));
 sky130_fd_sc_hd__nand2_1 _33824_ (.A(net1082),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[26] ),
    .Y(_12848_));
 sky130_fd_sc_hd__nand2_1 _33825_ (.A(net858),
    .B(\inst$top.soc.sram.read_port__data[26] ),
    .Y(_12849_));
 sky130_fd_sc_hd__o211ai_1 _33826_ (.A1(_12847_),
    .A2(net1084),
    .B1(_12848_),
    .C1(_12849_),
    .Y(_12850_));
 sky130_fd_sc_hd__inv_1 _33828_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[26] ),
    .Y(_12852_));
 sky130_fd_sc_hd__a21oi_1 _33829_ (.A1(net1800),
    .A2(_12852_),
    .B1(net2949),
    .Y(_12853_));
 sky130_fd_sc_hd__o21ai_0 _33830_ (.A1(net1799),
    .A2(net3037),
    .B1(_12853_),
    .Y(_12854_));
 sky130_fd_sc_hd__inv_2 _33831_ (.A(_12854_),
    .Y(_04170_));
 sky130_fd_sc_hd__inv_1 _33832_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[27] ),
    .Y(_12855_));
 sky130_fd_sc_hd__nand2_1 _33833_ (.A(net1082),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[27] ),
    .Y(_12856_));
 sky130_fd_sc_hd__nand2_1 _33834_ (.A(net858),
    .B(\inst$top.soc.sram.read_port__data[27] ),
    .Y(_12857_));
 sky130_fd_sc_hd__o211ai_1 _33835_ (.A1(_12855_),
    .A2(net1084),
    .B1(_12856_),
    .C1(_12857_),
    .Y(_12858_));
 sky130_fd_sc_hd__inv_1 _33836_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[27] ),
    .Y(_12859_));
 sky130_fd_sc_hd__a21oi_1 _33837_ (.A1(net1799),
    .A2(_12859_),
    .B1(net2948),
    .Y(_12860_));
 sky130_fd_sc_hd__o21ai_0 _33838_ (.A1(net1799),
    .A2(_12858_),
    .B1(_12860_),
    .Y(_12861_));
 sky130_fd_sc_hd__inv_2 _33839_ (.A(_12861_),
    .Y(_04171_));
 sky130_fd_sc_hd__inv_1 _33841_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[28] ),
    .Y(_12863_));
 sky130_fd_sc_hd__nand2_1 _33842_ (.A(net1082),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[28] ),
    .Y(_12864_));
 sky130_fd_sc_hd__nand2_1 _33843_ (.A(net858),
    .B(\inst$top.soc.sram.read_port__data[28] ),
    .Y(_12865_));
 sky130_fd_sc_hd__o211ai_1 _33844_ (.A1(_12863_),
    .A2(net1084),
    .B1(_12864_),
    .C1(_12865_),
    .Y(_12866_));
 sky130_fd_sc_hd__inv_1 _33845_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[28] ),
    .Y(_12867_));
 sky130_fd_sc_hd__a21oi_1 _33846_ (.A1(net1800),
    .A2(_12867_),
    .B1(net2949),
    .Y(_12868_));
 sky130_fd_sc_hd__o21ai_0 _33847_ (.A1(net1800),
    .A2(_12866_),
    .B1(_12868_),
    .Y(_12869_));
 sky130_fd_sc_hd__inv_2 _33848_ (.A(_12869_),
    .Y(_04172_));
 sky130_fd_sc_hd__inv_1 _33849_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[29] ),
    .Y(_12870_));
 sky130_fd_sc_hd__nand2_1 _33850_ (.A(net1083),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[29] ),
    .Y(_12871_));
 sky130_fd_sc_hd__nand2_1 _33851_ (.A(net860),
    .B(\inst$top.soc.sram.read_port__data[29] ),
    .Y(_12872_));
 sky130_fd_sc_hd__o211ai_1 _33852_ (.A1(_12870_),
    .A2(net1085),
    .B1(_12871_),
    .C1(_12872_),
    .Y(_12873_));
 sky130_fd_sc_hd__inv_1 _33853_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[29] ),
    .Y(_12874_));
 sky130_fd_sc_hd__a21oi_1 _33854_ (.A1(net1801),
    .A2(_12874_),
    .B1(net2950),
    .Y(_12875_));
 sky130_fd_sc_hd__o21ai_0 _33855_ (.A1(net1801),
    .A2(net3041),
    .B1(_12875_),
    .Y(_12876_));
 sky130_fd_sc_hd__inv_2 _33856_ (.A(_12876_),
    .Y(_04173_));
 sky130_fd_sc_hd__inv_1 _33857_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[2] ),
    .Y(_12877_));
 sky130_fd_sc_hd__inv_1 _33858_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[2] ),
    .Y(_12878_));
 sky130_fd_sc_hd__nand2_1 _33859_ (.A(net859),
    .B(\inst$top.soc.sram.read_port__data[2] ),
    .Y(_12879_));
 sky130_fd_sc_hd__o221ai_1 _33860_ (.A1(_12877_),
    .A2(net1084),
    .B1(_12878_),
    .B2(net1025),
    .C1(_12879_),
    .Y(_12880_));
 sky130_fd_sc_hd__inv_1 _33861_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[2] ),
    .Y(_12881_));
 sky130_fd_sc_hd__a21oi_1 _33862_ (.A1(net1799),
    .A2(_12881_),
    .B1(net2948),
    .Y(_12882_));
 sky130_fd_sc_hd__o21ai_0 _33863_ (.A1(net1799),
    .A2(_12880_),
    .B1(_12882_),
    .Y(_12883_));
 sky130_fd_sc_hd__inv_2 _33864_ (.A(_12883_),
    .Y(_04174_));
 sky130_fd_sc_hd__inv_1 _33865_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[30] ),
    .Y(_12884_));
 sky130_fd_sc_hd__nand2_1 _33866_ (.A(net1083),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[30] ),
    .Y(_12885_));
 sky130_fd_sc_hd__nand2_1 _33867_ (.A(net859),
    .B(\inst$top.soc.sram.read_port__data[30] ),
    .Y(_12886_));
 sky130_fd_sc_hd__o211ai_1 _33868_ (.A1(_12884_),
    .A2(net1087),
    .B1(_12885_),
    .C1(_12886_),
    .Y(_12887_));
 sky130_fd_sc_hd__inv_1 _33869_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[30] ),
    .Y(_12888_));
 sky130_fd_sc_hd__a21oi_1 _33870_ (.A1(net1799),
    .A2(_12888_),
    .B1(net2949),
    .Y(_12889_));
 sky130_fd_sc_hd__o21ai_0 _33871_ (.A1(net1800),
    .A2(net3040),
    .B1(_12889_),
    .Y(_12890_));
 sky130_fd_sc_hd__inv_2 _33872_ (.A(_12890_),
    .Y(_04175_));
 sky130_fd_sc_hd__inv_1 _33873_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[31] ),
    .Y(_12891_));
 sky130_fd_sc_hd__inv_1 _33874_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[31] ),
    .Y(_12892_));
 sky130_fd_sc_hd__nand2_1 _33875_ (.A(net860),
    .B(\inst$top.soc.sram.read_port__data[31] ),
    .Y(_12893_));
 sky130_fd_sc_hd__o221ai_1 _33876_ (.A1(_12891_),
    .A2(net1085),
    .B1(_12892_),
    .B2(net1025),
    .C1(_12893_),
    .Y(_12894_));
 sky130_fd_sc_hd__inv_1 _33877_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[31] ),
    .Y(_12895_));
 sky130_fd_sc_hd__a21oi_1 _33878_ (.A1(_12696_),
    .A2(_12895_),
    .B1(net2949),
    .Y(_12896_));
 sky130_fd_sc_hd__o21ai_0 _33879_ (.A1(net1802),
    .A2(_12894_),
    .B1(_12896_),
    .Y(_12897_));
 sky130_fd_sc_hd__inv_2 _33880_ (.A(_12897_),
    .Y(_04176_));
 sky130_fd_sc_hd__inv_1 _33881_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[3] ),
    .Y(_12898_));
 sky130_fd_sc_hd__inv_1 _33882_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[3] ),
    .Y(_12899_));
 sky130_fd_sc_hd__nand2_1 _33883_ (.A(net858),
    .B(\inst$top.soc.sram.read_port__data[3] ),
    .Y(_12900_));
 sky130_fd_sc_hd__o221ai_1 _33884_ (.A1(_12898_),
    .A2(net1084),
    .B1(_12899_),
    .B2(net1025),
    .C1(_12900_),
    .Y(_12901_));
 sky130_fd_sc_hd__inv_1 _33885_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[3] ),
    .Y(_12902_));
 sky130_fd_sc_hd__a21oi_1 _33887_ (.A1(net1801),
    .A2(_12902_),
    .B1(net2949),
    .Y(_12904_));
 sky130_fd_sc_hd__o21ai_0 _33888_ (.A1(net1801),
    .A2(_12901_),
    .B1(_12904_),
    .Y(_12905_));
 sky130_fd_sc_hd__inv_2 _33889_ (.A(_12905_),
    .Y(_04177_));
 sky130_fd_sc_hd__inv_1 _33890_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[4] ),
    .Y(_12906_));
 sky130_fd_sc_hd__inv_1 _33891_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[4] ),
    .Y(_12907_));
 sky130_fd_sc_hd__nand2_1 _33892_ (.A(net858),
    .B(\inst$top.soc.sram.read_port__data[4] ),
    .Y(_12908_));
 sky130_fd_sc_hd__o221ai_1 _33893_ (.A1(_12906_),
    .A2(net1084),
    .B1(_12907_),
    .B2(net1025),
    .C1(_12908_),
    .Y(_12909_));
 sky130_fd_sc_hd__inv_1 _33894_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[4] ),
    .Y(_12910_));
 sky130_fd_sc_hd__a21oi_1 _33895_ (.A1(net1802),
    .A2(_12910_),
    .B1(net2950),
    .Y(_12911_));
 sky130_fd_sc_hd__o21ai_0 _33896_ (.A1(net1802),
    .A2(_12909_),
    .B1(_12911_),
    .Y(_12912_));
 sky130_fd_sc_hd__inv_2 _33897_ (.A(_12912_),
    .Y(_04178_));
 sky130_fd_sc_hd__inv_1 _33898_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[5] ),
    .Y(_12913_));
 sky130_fd_sc_hd__inv_1 _33899_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[5] ),
    .Y(_12914_));
 sky130_fd_sc_hd__nand2_1 _33900_ (.A(net859),
    .B(\inst$top.soc.sram.read_port__data[5] ),
    .Y(_12915_));
 sky130_fd_sc_hd__o221ai_2 _33901_ (.A1(_12913_),
    .A2(net1087),
    .B1(_12914_),
    .B2(net1025),
    .C1(_12915_),
    .Y(_12916_));
 sky130_fd_sc_hd__inv_1 _33902_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[5] ),
    .Y(_12917_));
 sky130_fd_sc_hd__a21oi_1 _33903_ (.A1(net1801),
    .A2(_12917_),
    .B1(net2950),
    .Y(_12918_));
 sky130_fd_sc_hd__o21ai_0 _33904_ (.A1(net1801),
    .A2(_12916_),
    .B1(_12918_),
    .Y(_12919_));
 sky130_fd_sc_hd__inv_2 _33905_ (.A(_12919_),
    .Y(_04179_));
 sky130_fd_sc_hd__inv_1 _33906_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[6] ),
    .Y(_12920_));
 sky130_fd_sc_hd__inv_1 _33907_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[6] ),
    .Y(_12921_));
 sky130_fd_sc_hd__nand2_1 _33908_ (.A(net858),
    .B(\inst$top.soc.sram.read_port__data[6] ),
    .Y(_12922_));
 sky130_fd_sc_hd__o221ai_2 _33909_ (.A1(_12920_),
    .A2(net1084),
    .B1(_12921_),
    .B2(net1025),
    .C1(_12922_),
    .Y(_12923_));
 sky130_fd_sc_hd__inv_1 _33910_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[6] ),
    .Y(_12924_));
 sky130_fd_sc_hd__a21oi_1 _33911_ (.A1(net1801),
    .A2(_12924_),
    .B1(net2950),
    .Y(_12925_));
 sky130_fd_sc_hd__o21ai_0 _33912_ (.A1(net1802),
    .A2(_12923_),
    .B1(_12925_),
    .Y(_12926_));
 sky130_fd_sc_hd__inv_2 _33913_ (.A(_12926_),
    .Y(_04180_));
 sky130_fd_sc_hd__inv_1 _33914_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[7] ),
    .Y(_12927_));
 sky130_fd_sc_hd__inv_1 _33915_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[7] ),
    .Y(_12928_));
 sky130_fd_sc_hd__nand2_1 _33916_ (.A(net860),
    .B(\inst$top.soc.sram.read_port__data[7] ),
    .Y(_12929_));
 sky130_fd_sc_hd__o221ai_1 _33917_ (.A1(_12927_),
    .A2(net1085),
    .B1(_12928_),
    .B2(net1025),
    .C1(_12929_),
    .Y(_12930_));
 sky130_fd_sc_hd__inv_1 _33918_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[7] ),
    .Y(_12931_));
 sky130_fd_sc_hd__a21oi_1 _33919_ (.A1(net1804),
    .A2(_12931_),
    .B1(net2988),
    .Y(_12932_));
 sky130_fd_sc_hd__o21ai_0 _33920_ (.A1(net1805),
    .A2(net3039),
    .B1(_12932_),
    .Y(_12933_));
 sky130_fd_sc_hd__inv_2 _33921_ (.A(_12933_),
    .Y(_04181_));
 sky130_fd_sc_hd__inv_1 _33922_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[8] ),
    .Y(_12934_));
 sky130_fd_sc_hd__nand2_1 _33923_ (.A(net1083),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[8] ),
    .Y(_12935_));
 sky130_fd_sc_hd__nand2_1 _33924_ (.A(net860),
    .B(\inst$top.soc.sram.read_port__data[8] ),
    .Y(_12936_));
 sky130_fd_sc_hd__o211ai_1 _33925_ (.A1(_12934_),
    .A2(net1085),
    .B1(_12935_),
    .C1(_12936_),
    .Y(_12937_));
 sky130_fd_sc_hd__inv_1 _33926_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[8] ),
    .Y(_12938_));
 sky130_fd_sc_hd__a21oi_1 _33927_ (.A1(net1804),
    .A2(_12938_),
    .B1(net2980),
    .Y(_12939_));
 sky130_fd_sc_hd__o21ai_0 _33928_ (.A1(net1804),
    .A2(_12937_),
    .B1(_12939_),
    .Y(_12940_));
 sky130_fd_sc_hd__inv_2 _33929_ (.A(_12940_),
    .Y(_04182_));
 sky130_fd_sc_hd__inv_1 _33930_ (.A(\inst$top.soc.wb_to_csr.wb_bus__dat_r[9] ),
    .Y(_12941_));
 sky130_fd_sc_hd__nand2_1 _33931_ (.A(net1082),
    .B(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[9] ),
    .Y(_12942_));
 sky130_fd_sc_hd__nand2_1 _33932_ (.A(net860),
    .B(\inst$top.soc.sram.read_port__data[9] ),
    .Y(_12943_));
 sky130_fd_sc_hd__o211ai_1 _33933_ (.A1(_12941_),
    .A2(net1086),
    .B1(_12942_),
    .C1(_12943_),
    .Y(_12944_));
 sky130_fd_sc_hd__inv_1 _33934_ (.A(\inst$top.soc.cpu.fetch.ibus_rdata[9] ),
    .Y(_12945_));
 sky130_fd_sc_hd__a21oi_1 _33935_ (.A1(net1804),
    .A2(_12945_),
    .B1(net2980),
    .Y(_12946_));
 sky130_fd_sc_hd__o21ai_0 _33936_ (.A1(net1804),
    .A2(_12944_),
    .B1(_12946_),
    .Y(_12947_));
 sky130_fd_sc_hd__inv_2 _33937_ (.A(_12947_),
    .Y(_04183_));
 sky130_fd_sc_hd__nor2_1 _33938_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[0] ),
    .B(net704),
    .Y(_12948_));
 sky130_fd_sc_hd__xor2_1 _33939_ (.A(\inst$top.soc.cpu.sink__payload$24[32] ),
    .B(net2754),
    .X(_12949_));
 sky130_fd_sc_hd__o22ai_1 _33940_ (.A1(net2718),
    .A2(_19831_),
    .B1(_19833_),
    .B2(net2700),
    .Y(_12950_));
 sky130_fd_sc_hd__nand2_1 _33941_ (.A(_19834_),
    .B(net2695),
    .Y(_12951_));
 sky130_fd_sc_hd__o22ai_1 _33942_ (.A1(net2689),
    .A2(_19826_),
    .B1(_19834_),
    .B2(net2695),
    .Y(_12952_));
 sky130_fd_sc_hd__a221oi_1 _33943_ (.A1(_19831_),
    .A2(net2718),
    .B1(_19826_),
    .B2(net2689),
    .C1(_12952_),
    .Y(_12953_));
 sky130_fd_sc_hd__o2111ai_1 _33944_ (.A1(\inst$top.soc.cpu.sink__payload$24[34] ),
    .A2(net2417),
    .B1(_19830_),
    .C1(_12951_),
    .D1(_12953_),
    .Y(_12954_));
 sky130_fd_sc_hd__nor3_1 _33945_ (.A(_12949_),
    .B(_12950_),
    .C(_12954_),
    .Y(_12955_));
 sky130_fd_sc_hd__nand4_1 _33946_ (.A(_20331_),
    .B(_20334_),
    .C(_20342_),
    .D(_12955_),
    .Y(_12956_));
 sky130_fd_sc_hd__clkinv_1 _33947_ (.A(_12956_),
    .Y(_12957_));
 sky130_fd_sc_hd__nor2_2 _33949_ (.A(_20347_),
    .B(_20331_),
    .Y(_12959_));
 sky130_fd_sc_hd__inv_1 _33950_ (.A(net786),
    .Y(_12960_));
 sky130_fd_sc_hd__clkinv_1 _33951_ (.A(net2862),
    .Y(_12961_));
 sky130_fd_sc_hd__o21ai_0 _33953_ (.A1(net2848),
    .A2(_03083_),
    .B1(_20397_),
    .Y(_12963_));
 sky130_fd_sc_hd__o21ai_0 _33956_ (.A1(net2849),
    .A2(net2842),
    .B1(_09917_),
    .Y(_12966_));
 sky130_fd_sc_hd__inv_1 _33957_ (.A(_12966_),
    .Y(_12967_));
 sky130_fd_sc_hd__nand2_1 _33959_ (.A(\inst$top.soc.cpu.sink__payload$12[144] ),
    .B(\inst$top.soc.cpu.sink__payload$12[143] ),
    .Y(_12969_));
 sky130_fd_sc_hd__nor2_1 _33960_ (.A(net2849),
    .B(\inst$top.soc.cpu.d.sink__payload.csr_fmt_i ),
    .Y(_12970_));
 sky130_fd_sc_hd__nor2_1 _33961_ (.A(_12969_),
    .B(_12970_),
    .Y(_12971_));
 sky130_fd_sc_hd__nor2_1 _33963_ (.A(\inst$top.soc.cpu.sink__payload$12[143] ),
    .B(_09912_),
    .Y(_12973_));
 sky130_fd_sc_hd__inv_1 _33964_ (.A(_12973_),
    .Y(_12974_));
 sky130_fd_sc_hd__nor2_1 _33965_ (.A(_12970_),
    .B(_12974_),
    .Y(_12975_));
 sky130_fd_sc_hd__inv_1 _33966_ (.A(_12975_),
    .Y(_12976_));
 sky130_fd_sc_hd__nor2_1 _33967_ (.A(_03090_),
    .B(net1231),
    .Y(_12977_));
 sky130_fd_sc_hd__a221oi_1 _33968_ (.A1(net1798),
    .A2(_03087_),
    .B1(net1871),
    .B2(_03086_),
    .C1(_12977_),
    .Y(_12978_));
 sky130_fd_sc_hd__inv_1 _33969_ (.A(_12978_),
    .Y(_12979_));
 sky130_fd_sc_hd__nor2_1 _33970_ (.A(net2019),
    .B(_12979_),
    .Y(_12980_));
 sky130_fd_sc_hd__a211oi_1 _33971_ (.A1(net2019),
    .A2(_12963_),
    .B1(net2855),
    .C1(_12980_),
    .Y(_12981_));
 sky130_fd_sc_hd__inv_1 _33972_ (.A(_12981_),
    .Y(_12982_));
 sky130_fd_sc_hd__nand3_1 _33973_ (.A(_20331_),
    .B(_20334_),
    .C(_20343_),
    .Y(_12983_));
 sky130_fd_sc_hd__clkinv_1 _33974_ (.A(net785),
    .Y(_12984_));
 sky130_fd_sc_hd__nor2_1 _33977_ (.A(\inst$top.soc.cpu.sink__payload$18[109] ),
    .B(net2834),
    .Y(_12987_));
 sky130_fd_sc_hd__inv_1 _33980_ (.A(\inst$top.soc.cpu.shifter.m_result$7[31] ),
    .Y(_12990_));
 sky130_fd_sc_hd__o21ai_0 _33982_ (.A1(net2871),
    .A2(_12990_),
    .B1(net2840),
    .Y(_12992_));
 sky130_fd_sc_hd__a21oi_1 _33983_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[0] ),
    .A2(net2871),
    .B1(_12992_),
    .Y(_12993_));
 sky130_fd_sc_hd__inv_2 _33984_ (.A(\inst$top.soc.cpu.d.sink__payload$6.divide ),
    .Y(_12994_));
 sky130_fd_sc_hd__o21ai_0 _33986_ (.A1(_12987_),
    .A2(_12993_),
    .B1(net2013),
    .Y(_12996_));
 sky130_fd_sc_hd__inv_1 _33987_ (.A(net2829),
    .Y(_12997_));
 sky130_fd_sc_hd__a21oi_1 _33991_ (.A1(net2923),
    .A2(\inst$top.soc.cpu.divider.remainder[0] ),
    .B1(net2012),
    .Y(_13001_));
 sky130_fd_sc_hd__o21ai_2 _33992_ (.A1(net2922),
    .A2(_02846_),
    .B1(_13001_),
    .Y(_13002_));
 sky130_fd_sc_hd__nand3_1 _33993_ (.A(_12996_),
    .B(_12997_),
    .C(_13002_),
    .Y(_13003_));
 sky130_fd_sc_hd__nand2_1 _33995_ (.A(\inst$top.soc.cpu.d.sink__payload$6.condition_met ),
    .B(net2829),
    .Y(_13005_));
 sky130_fd_sc_hd__nand2_1 _33996_ (.A(_13003_),
    .B(_13005_),
    .Y(_13006_));
 sky130_fd_sc_hd__nand2_1 _33997_ (.A(_12984_),
    .B(_13006_),
    .Y(_13007_));
 sky130_fd_sc_hd__o21ai_0 _33998_ (.A1(net736),
    .A2(_12982_),
    .B1(_13007_),
    .Y(_13008_));
 sky130_fd_sc_hd__a21oi_1 _33999_ (.A1(net737),
    .A2(net1064),
    .B1(_13008_),
    .Y(_13009_));
 sky130_fd_sc_hd__nand2_1 _34000_ (.A(net704),
    .B(_13009_),
    .Y(_13010_));
 sky130_fd_sc_hd__nand2_1 _34001_ (.A(_13010_),
    .B(net2152),
    .Y(_13011_));
 sky130_fd_sc_hd__nor2_4 _34002_ (.A(_12948_),
    .B(_13011_),
    .Y(_04184_));
 sky130_fd_sc_hd__nor2_1 _34004_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[10] ),
    .B(net709),
    .Y(_13013_));
 sky130_fd_sc_hd__inv_1 _34006_ (.A(\inst$top.soc.cpu.sink__payload$18[119] ),
    .Y(_13015_));
 sky130_fd_sc_hd__nor2_1 _34007_ (.A(net2835),
    .B(_13015_),
    .Y(_13016_));
 sky130_fd_sc_hd__inv_1 _34009_ (.A(\inst$top.soc.cpu.shifter.m_result$7[10] ),
    .Y(_13018_));
 sky130_fd_sc_hd__o21ai_0 _34010_ (.A1(net2870),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[21] ),
    .B1(net2835),
    .Y(_13019_));
 sky130_fd_sc_hd__a21oi_1 _34011_ (.A1(net2870),
    .A2(_13018_),
    .B1(_13019_),
    .Y(_13020_));
 sky130_fd_sc_hd__o21ai_0 _34013_ (.A1(_13016_),
    .A2(_13020_),
    .B1(net2014),
    .Y(_13022_));
 sky130_fd_sc_hd__a21oi_1 _34014_ (.A1(_10333_),
    .A2(net2916),
    .B1(net2009),
    .Y(_13023_));
 sky130_fd_sc_hd__o21ai_2 _34015_ (.A1(net2916),
    .A2(\inst$top.soc.cpu.divider.quotient[10] ),
    .B1(_13023_),
    .Y(_13024_));
 sky130_fd_sc_hd__a21oi_1 _34017_ (.A1(_13022_),
    .A2(_13024_),
    .B1(net2830),
    .Y(_13026_));
 sky130_fd_sc_hd__inv_1 _34018_ (.A(_13026_),
    .Y(_13027_));
 sky130_fd_sc_hd__nand2_1 _34021_ (.A(\inst$top.soc.cpu.sink__payload$12[9] ),
    .B(\inst$top.soc.cpu.sink__payload$12[8] ),
    .Y(_13030_));
 sky130_fd_sc_hd__nand2_1 _34022_ (.A(\inst$top.soc.cpu.sink__payload$12[4] ),
    .B(_03112_),
    .Y(_13031_));
 sky130_fd_sc_hd__nand2_1 _34023_ (.A(\inst$top.soc.cpu.sink__payload$12[6] ),
    .B(\inst$top.soc.cpu.sink__payload$12[5] ),
    .Y(_13032_));
 sky130_fd_sc_hd__nor3_1 _34024_ (.A(_20623_),
    .B(_13031_),
    .C(_13032_),
    .Y(_13033_));
 sky130_fd_sc_hd__inv_1 _34025_ (.A(_13033_),
    .Y(_13034_));
 sky130_fd_sc_hd__nor2_1 _34026_ (.A(_13030_),
    .B(_13034_),
    .Y(_13035_));
 sky130_fd_sc_hd__nor2_1 _34027_ (.A(_20705_),
    .B(_13035_),
    .Y(_13036_));
 sky130_fd_sc_hd__nand2_1 _34028_ (.A(_13035_),
    .B(_20705_),
    .Y(_13037_));
 sky130_fd_sc_hd__nand2_1 _34030_ (.A(_13037_),
    .B(net2853),
    .Y(_13039_));
 sky130_fd_sc_hd__inv_1 _34031_ (.A(_03033_),
    .Y(_13040_));
 sky130_fd_sc_hd__inv_1 _34032_ (.A(net2865),
    .Y(_13041_));
 sky130_fd_sc_hd__nand2_1 _34033_ (.A(_03049_),
    .B(_03054_),
    .Y(_13042_));
 sky130_fd_sc_hd__inv_1 _34034_ (.A(_13042_),
    .Y(_13043_));
 sky130_fd_sc_hd__nand3_1 _34035_ (.A(_13043_),
    .B(_03039_),
    .C(_03044_),
    .Y(_13044_));
 sky130_fd_sc_hd__a21oi_1 _34036_ (.A1(_03070_),
    .A2(_03075_),
    .B1(_03069_),
    .Y(_13045_));
 sky130_fd_sc_hd__nand3b_1 _34037_ (.A_N(_00170_),
    .B(_03070_),
    .C(_03076_),
    .Y(_13046_));
 sky130_fd_sc_hd__nand2_1 _34038_ (.A(_13045_),
    .B(_13046_),
    .Y(_13047_));
 sky130_fd_sc_hd__nand2_1 _34039_ (.A(_03060_),
    .B(_03065_),
    .Y(_13048_));
 sky130_fd_sc_hd__inv_1 _34040_ (.A(_13048_),
    .Y(_13049_));
 sky130_fd_sc_hd__nand2_1 _34041_ (.A(_03060_),
    .B(_03064_),
    .Y(_13050_));
 sky130_fd_sc_hd__inv_1 _34042_ (.A(_03059_),
    .Y(_13051_));
 sky130_fd_sc_hd__nand2_1 _34043_ (.A(_13050_),
    .B(_13051_),
    .Y(_13052_));
 sky130_fd_sc_hd__a21oi_1 _34044_ (.A1(_13047_),
    .A2(_13049_),
    .B1(_13052_),
    .Y(_13053_));
 sky130_fd_sc_hd__nand2_1 _34045_ (.A(_03039_),
    .B(_03044_),
    .Y(_13054_));
 sky130_fd_sc_hd__a21oi_1 _34046_ (.A1(_03049_),
    .A2(_03053_),
    .B1(_03048_),
    .Y(_13055_));
 sky130_fd_sc_hd__a21oi_1 _34047_ (.A1(_03039_),
    .A2(_03043_),
    .B1(_03038_),
    .Y(_13056_));
 sky130_fd_sc_hd__o21ai_0 _34048_ (.A1(_13054_),
    .A2(_13055_),
    .B1(_13056_),
    .Y(_13057_));
 sky130_fd_sc_hd__o21bai_1 _34049_ (.A1(_13044_),
    .A2(_13053_),
    .B1_N(_13057_),
    .Y(_13058_));
 sky130_fd_sc_hd__nor2_1 _34050_ (.A(_03060_),
    .B(_03065_),
    .Y(_13059_));
 sky130_fd_sc_hd__inv_1 _34051_ (.A(_13059_),
    .Y(_13060_));
 sky130_fd_sc_hd__inv_1 _34052_ (.A(_03070_),
    .Y(_13061_));
 sky130_fd_sc_hd__a21oi_2 _34053_ (.A1(_13061_),
    .A2(_03078_),
    .B1(_03072_),
    .Y(_13062_));
 sky130_fd_sc_hd__inv_1 _34054_ (.A(_03060_),
    .Y(_13063_));
 sky130_fd_sc_hd__a21oi_1 _34055_ (.A1(_13063_),
    .A2(_00230_),
    .B1(_00273_),
    .Y(_13064_));
 sky130_fd_sc_hd__o21ai_0 _34056_ (.A1(_13060_),
    .A2(_13062_),
    .B1(_13064_),
    .Y(_13065_));
 sky130_fd_sc_hd__nor2_1 _34057_ (.A(_03039_),
    .B(_03044_),
    .Y(_13066_));
 sky130_fd_sc_hd__nor2_1 _34058_ (.A(_03049_),
    .B(_03054_),
    .Y(_13067_));
 sky130_fd_sc_hd__nand2_1 _34059_ (.A(_13066_),
    .B(_13067_),
    .Y(_13068_));
 sky130_fd_sc_hd__inv_1 _34060_ (.A(_13068_),
    .Y(_13069_));
 sky130_fd_sc_hd__nand2_1 _34061_ (.A(_13065_),
    .B(_13069_),
    .Y(_13070_));
 sky130_fd_sc_hd__inv_1 _34062_ (.A(_03076_),
    .Y(_13071_));
 sky130_fd_sc_hd__nand3_1 _34063_ (.A(_13059_),
    .B(_13061_),
    .C(_13071_),
    .Y(_13072_));
 sky130_fd_sc_hd__nor2_1 _34064_ (.A(_13068_),
    .B(_13072_),
    .Y(_13073_));
 sky130_fd_sc_hd__inv_1 _34065_ (.A(_00165_),
    .Y(_13074_));
 sky130_fd_sc_hd__nand2_1 _34066_ (.A(_13073_),
    .B(_13074_),
    .Y(_13075_));
 sky130_fd_sc_hd__inv_1 _34067_ (.A(_00391_),
    .Y(_13076_));
 sky130_fd_sc_hd__o21ai_0 _34068_ (.A1(_03049_),
    .A2(_00325_),
    .B1(_13076_),
    .Y(_13077_));
 sky130_fd_sc_hd__o21bai_1 _34069_ (.A1(_03039_),
    .A2(_00464_),
    .B1_N(_00531_),
    .Y(_13078_));
 sky130_fd_sc_hd__a21oi_1 _34070_ (.A1(_13077_),
    .A2(_13066_),
    .B1(_13078_),
    .Y(_13079_));
 sky130_fd_sc_hd__nand3_1 _34071_ (.A(_13070_),
    .B(_13075_),
    .C(_13079_),
    .Y(_13080_));
 sky130_fd_sc_hd__nand2_1 _34072_ (.A(_13080_),
    .B(net2008),
    .Y(_13081_));
 sky130_fd_sc_hd__o21ai_2 _34073_ (.A1(net2006),
    .A2(_13058_),
    .B1(_13081_),
    .Y(_13082_));
 sky130_fd_sc_hd__or2_2 _34074_ (.A(_13040_),
    .B(_13082_),
    .X(_13083_));
 sky130_fd_sc_hd__nand2_1 _34075_ (.A(_13082_),
    .B(_13040_),
    .Y(_13084_));
 sky130_fd_sc_hd__nand3_1 _34076_ (.A(_13083_),
    .B(net2214),
    .C(_13084_),
    .Y(_13085_));
 sky130_fd_sc_hd__nand2_1 _34077_ (.A(_13085_),
    .B(_20721_),
    .Y(_13086_));
 sky130_fd_sc_hd__nand2_1 _34078_ (.A(_13086_),
    .B(net2019),
    .Y(_13087_));
 sky130_fd_sc_hd__nand2_1 _34080_ (.A(net1797),
    .B(_03159_),
    .Y(_13089_));
 sky130_fd_sc_hd__nand2_1 _34081_ (.A(net1870),
    .B(_03158_),
    .Y(_13090_));
 sky130_fd_sc_hd__o211ai_1 _34082_ (.A1(_03162_),
    .A2(net1231),
    .B1(_13089_),
    .C1(_13090_),
    .Y(_13091_));
 sky130_fd_sc_hd__a21oi_1 _34083_ (.A1(_13091_),
    .A2(net2861),
    .B1(net2855),
    .Y(_13092_));
 sky130_fd_sc_hd__nand2_1 _34084_ (.A(_13087_),
    .B(_13092_),
    .Y(_13093_));
 sky130_fd_sc_hd__o21a_1 _34085_ (.A1(_13036_),
    .A2(_13039_),
    .B1(_13093_),
    .X(_13094_));
 sky130_fd_sc_hd__inv_1 _34086_ (.A(_13094_),
    .Y(_13095_));
 sky130_fd_sc_hd__o22ai_1 _34087_ (.A1(_13027_),
    .A2(net783),
    .B1(net736),
    .B2(_13095_),
    .Y(_13096_));
 sky130_fd_sc_hd__a21oi_1 _34088_ (.A1(net737),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[10] ),
    .B1(_13096_),
    .Y(_13097_));
 sky130_fd_sc_hd__nand2_1 _34089_ (.A(net709),
    .B(_13097_),
    .Y(_13098_));
 sky130_fd_sc_hd__nand2_1 _34090_ (.A(_13098_),
    .B(net2156),
    .Y(_13099_));
 sky130_fd_sc_hd__nor2_2 _34091_ (.A(_13013_),
    .B(_13099_),
    .Y(_04185_));
 sky130_fd_sc_hd__nor2_1 _34092_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[11] ),
    .B(net702),
    .Y(_13100_));
 sky130_fd_sc_hd__inv_1 _34093_ (.A(\inst$top.soc.cpu.sink__payload$18[120] ),
    .Y(_13101_));
 sky130_fd_sc_hd__inv_1 _34094_ (.A(net2871),
    .Y(_13102_));
 sky130_fd_sc_hd__nor2_1 _34096_ (.A(\inst$top.soc.cpu.shifter.m_result$7[11] ),
    .B(net2002),
    .Y(_13104_));
 sky130_fd_sc_hd__o21ai_0 _34097_ (.A1(net2869),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[20] ),
    .B1(net2841),
    .Y(_13105_));
 sky130_fd_sc_hd__o22ai_1 _34098_ (.A1(_13101_),
    .A2(net2833),
    .B1(_13104_),
    .B2(_13105_),
    .Y(_13106_));
 sky130_fd_sc_hd__nand2_1 _34099_ (.A(_13106_),
    .B(net2014),
    .Y(_13107_));
 sky130_fd_sc_hd__a21oi_1 _34102_ (.A1(_10375_),
    .A2(net2917),
    .B1(net2009),
    .Y(_13110_));
 sky130_fd_sc_hd__o21ai_4 _34103_ (.A1(net2917),
    .A2(\inst$top.soc.cpu.divider.quotient[11] ),
    .B1(_13110_),
    .Y(_13111_));
 sky130_fd_sc_hd__a21oi_1 _34104_ (.A1(_13107_),
    .A2(_13111_),
    .B1(net2830),
    .Y(_13112_));
 sky130_fd_sc_hd__inv_1 _34105_ (.A(_13112_),
    .Y(_13113_));
 sky130_fd_sc_hd__nand2_1 _34106_ (.A(\inst$top.soc.cpu.sink__payload$12[8] ),
    .B(\inst$top.soc.cpu.sink__payload$12[7] ),
    .Y(_13114_));
 sky130_fd_sc_hd__nor3_1 _34107_ (.A(_20705_),
    .B(_20685_),
    .C(_13114_),
    .Y(_13115_));
 sky130_fd_sc_hd__nand3_1 _34108_ (.A(\inst$top.soc.cpu.sink__payload$12[4] ),
    .B(\inst$top.soc.cpu.sink__payload$12[3] ),
    .C(\inst$top.soc.cpu.sink__payload$12[2] ),
    .Y(_13116_));
 sky130_fd_sc_hd__nor2_1 _34109_ (.A(_13032_),
    .B(_13116_),
    .Y(_13117_));
 sky130_fd_sc_hd__nand2_1 _34110_ (.A(_13115_),
    .B(_13117_),
    .Y(_13118_));
 sky130_fd_sc_hd__nor2_1 _34111_ (.A(_20726_),
    .B(_13118_),
    .Y(_13119_));
 sky130_fd_sc_hd__nand2_1 _34112_ (.A(_13118_),
    .B(_20726_),
    .Y(_13120_));
 sky130_fd_sc_hd__nand2_1 _34114_ (.A(_13120_),
    .B(net2853),
    .Y(_13122_));
 sky130_fd_sc_hd__nand2_1 _34117_ (.A(net1797),
    .B(_03166_),
    .Y(_13125_));
 sky130_fd_sc_hd__nand2_1 _34119_ (.A(net1870),
    .B(_03165_),
    .Y(_13127_));
 sky130_fd_sc_hd__o211ai_1 _34120_ (.A1(_03169_),
    .A2(net1231),
    .B1(_13125_),
    .C1(_13127_),
    .Y(_13128_));
 sky130_fd_sc_hd__inv_1 _34121_ (.A(net2852),
    .Y(_13129_));
 sky130_fd_sc_hd__o21ai_0 _34123_ (.A1(net2018),
    .A2(_13128_),
    .B1(_13129_),
    .Y(_13131_));
 sky130_fd_sc_hd__nor2_1 _34125_ (.A(_03054_),
    .B(_03060_),
    .Y(_13133_));
 sky130_fd_sc_hd__inv_1 _34126_ (.A(_13133_),
    .Y(_13134_));
 sky130_fd_sc_hd__inv_1 _34127_ (.A(_03065_),
    .Y(_13135_));
 sky130_fd_sc_hd__a21oi_1 _34128_ (.A1(_13135_),
    .A2(_03072_),
    .B1(_00230_),
    .Y(_13136_));
 sky130_fd_sc_hd__inv_1 _34129_ (.A(_03054_),
    .Y(_13137_));
 sky130_fd_sc_hd__a21oi_1 _34130_ (.A1(_13137_),
    .A2(_00273_),
    .B1(_03056_),
    .Y(_13138_));
 sky130_fd_sc_hd__o21ai_0 _34131_ (.A1(_13134_),
    .A2(_13136_),
    .B1(_13138_),
    .Y(_13139_));
 sky130_fd_sc_hd__nor2_1 _34132_ (.A(_03033_),
    .B(_03039_),
    .Y(_13140_));
 sky130_fd_sc_hd__inv_1 _34133_ (.A(_13140_),
    .Y(_13141_));
 sky130_fd_sc_hd__nor2_1 _34134_ (.A(_03044_),
    .B(_03049_),
    .Y(_13142_));
 sky130_fd_sc_hd__inv_1 _34135_ (.A(_13142_),
    .Y(_13143_));
 sky130_fd_sc_hd__nor2_1 _34136_ (.A(_13141_),
    .B(_13143_),
    .Y(_13144_));
 sky130_fd_sc_hd__o21ai_0 _34137_ (.A1(_03044_),
    .A2(_13076_),
    .B1(_00464_),
    .Y(_13145_));
 sky130_fd_sc_hd__nand2_1 _34138_ (.A(_13145_),
    .B(_13140_),
    .Y(_13146_));
 sky130_fd_sc_hd__a21oi_1 _34139_ (.A1(_13040_),
    .A2(_00531_),
    .B1(_03035_),
    .Y(_13147_));
 sky130_fd_sc_hd__nand2_1 _34140_ (.A(_13146_),
    .B(_13147_),
    .Y(_13148_));
 sky130_fd_sc_hd__a21oi_1 _34141_ (.A1(_13139_),
    .A2(_13144_),
    .B1(_13148_),
    .Y(_13149_));
 sky130_fd_sc_hd__nor2_1 _34142_ (.A(_03065_),
    .B(_03070_),
    .Y(_13150_));
 sky130_fd_sc_hd__nand2_1 _34143_ (.A(_13133_),
    .B(_13150_),
    .Y(_13151_));
 sky130_fd_sc_hd__inv_1 _34144_ (.A(_13144_),
    .Y(_13152_));
 sky130_fd_sc_hd__nor2_1 _34145_ (.A(_13151_),
    .B(_13152_),
    .Y(_13153_));
 sky130_fd_sc_hd__inv_1 _34146_ (.A(_03080_),
    .Y(_13154_));
 sky130_fd_sc_hd__a21oi_1 _34147_ (.A1(_13154_),
    .A2(\inst$top.soc.cpu.multiplier.x_prod[0] ),
    .B1(_03081_),
    .Y(_13155_));
 sky130_fd_sc_hd__o21ai_0 _34148_ (.A1(_03076_),
    .A2(_13155_),
    .B1(_00192_),
    .Y(_13156_));
 sky130_fd_sc_hd__nand2_1 _34149_ (.A(_13153_),
    .B(_13156_),
    .Y(_13157_));
 sky130_fd_sc_hd__nand2_1 _34150_ (.A(_13149_),
    .B(_13157_),
    .Y(_13158_));
 sky130_fd_sc_hd__a21o_1 _34151_ (.A1(_03076_),
    .A2(_03079_),
    .B1(_03075_),
    .X(_13159_));
 sky130_fd_sc_hd__nand2_1 _34152_ (.A(_03065_),
    .B(_03070_),
    .Y(_13160_));
 sky130_fd_sc_hd__inv_1 _34153_ (.A(_13160_),
    .Y(_13161_));
 sky130_fd_sc_hd__nand2_1 _34154_ (.A(_13159_),
    .B(_13161_),
    .Y(_13162_));
 sky130_fd_sc_hd__a21oi_1 _34155_ (.A1(_03065_),
    .A2(_03069_),
    .B1(_03064_),
    .Y(_13163_));
 sky130_fd_sc_hd__nand2_1 _34156_ (.A(_13162_),
    .B(_13163_),
    .Y(_13164_));
 sky130_fd_sc_hd__nand2_1 _34157_ (.A(_03044_),
    .B(_03049_),
    .Y(_13165_));
 sky130_fd_sc_hd__inv_1 _34158_ (.A(_13165_),
    .Y(_13166_));
 sky130_fd_sc_hd__nand2_1 _34159_ (.A(_03054_),
    .B(_03060_),
    .Y(_13167_));
 sky130_fd_sc_hd__inv_1 _34160_ (.A(_13167_),
    .Y(_13168_));
 sky130_fd_sc_hd__nand3_1 _34161_ (.A(_13164_),
    .B(_13166_),
    .C(_13168_),
    .Y(_13169_));
 sky130_fd_sc_hd__a21oi_1 _34162_ (.A1(_03054_),
    .A2(_03059_),
    .B1(_03053_),
    .Y(_13170_));
 sky130_fd_sc_hd__inv_1 _34163_ (.A(_13170_),
    .Y(_13171_));
 sky130_fd_sc_hd__a21o_1 _34164_ (.A1(_03044_),
    .A2(_03048_),
    .B1(_03043_),
    .X(_13172_));
 sky130_fd_sc_hd__a21oi_1 _34165_ (.A1(_13171_),
    .A2(_13166_),
    .B1(_13172_),
    .Y(_13173_));
 sky130_fd_sc_hd__nand2_1 _34166_ (.A(_03076_),
    .B(_03080_),
    .Y(_13174_));
 sky130_fd_sc_hd__nand2_1 _34167_ (.A(_13166_),
    .B(_13168_),
    .Y(_13175_));
 sky130_fd_sc_hd__nor3_1 _34168_ (.A(_13174_),
    .B(_13160_),
    .C(_13175_),
    .Y(_13176_));
 sky130_fd_sc_hd__inv_1 _34169_ (.A(_00169_),
    .Y(_13177_));
 sky130_fd_sc_hd__nand2_1 _34170_ (.A(_13176_),
    .B(_13177_),
    .Y(_13178_));
 sky130_fd_sc_hd__nand3_1 _34171_ (.A(_13169_),
    .B(_13173_),
    .C(_13178_),
    .Y(_13179_));
 sky130_fd_sc_hd__nand2_1 _34172_ (.A(_03033_),
    .B(_03039_),
    .Y(_13180_));
 sky130_fd_sc_hd__inv_1 _34173_ (.A(_13180_),
    .Y(_13181_));
 sky130_fd_sc_hd__nand2_1 _34174_ (.A(_13179_),
    .B(_13181_),
    .Y(_13182_));
 sky130_fd_sc_hd__a21oi_1 _34175_ (.A1(_03033_),
    .A2(_03038_),
    .B1(_03032_),
    .Y(_13183_));
 sky130_fd_sc_hd__nand2_1 _34176_ (.A(_13182_),
    .B(_13183_),
    .Y(_13184_));
 sky130_fd_sc_hd__nand2_1 _34177_ (.A(_13184_),
    .B(net2867),
    .Y(_13185_));
 sky130_fd_sc_hd__o21ai_0 _34178_ (.A1(net2867),
    .A2(_13158_),
    .B1(_13185_),
    .Y(_13186_));
 sky130_fd_sc_hd__xor2_4 _34179_ (.A(_03027_),
    .B(_13186_),
    .X(_13187_));
 sky130_fd_sc_hd__nand2_1 _34180_ (.A(_20747_),
    .B(net2018),
    .Y(_13188_));
 sky130_fd_sc_hd__a21oi_1 _34181_ (.A1(_13187_),
    .A2(net2214),
    .B1(_13188_),
    .Y(_13189_));
 sky130_fd_sc_hd__o22ai_1 _34182_ (.A1(_13119_),
    .A2(_13122_),
    .B1(_13131_),
    .B2(_13189_),
    .Y(_13190_));
 sky130_fd_sc_hd__nand2_1 _34184_ (.A(_13190_),
    .B(net787),
    .Y(_13192_));
 sky130_fd_sc_hd__nand2_1 _34185_ (.A(net738),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[11] ),
    .Y(_13193_));
 sky130_fd_sc_hd__o211ai_1 _34186_ (.A1(net784),
    .A2(_13113_),
    .B1(_13192_),
    .C1(_13193_),
    .Y(_13194_));
 sky130_fd_sc_hd__o21ai_1 _34187_ (.A1(_13194_),
    .A2(net654),
    .B1(net2155),
    .Y(_13195_));
 sky130_fd_sc_hd__nor2_4 _34188_ (.A(_13100_),
    .B(_13195_),
    .Y(_04186_));
 sky130_fd_sc_hd__nor2_1 _34189_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[12] ),
    .B(net713),
    .Y(_13196_));
 sky130_fd_sc_hd__nor2_1 _34191_ (.A(_03027_),
    .B(_03033_),
    .Y(_13198_));
 sky130_fd_sc_hd__nand2_1 _34192_ (.A(_13080_),
    .B(_13198_),
    .Y(_13199_));
 sky130_fd_sc_hd__inv_1 _34193_ (.A(_03027_),
    .Y(_13200_));
 sky130_fd_sc_hd__a21oi_1 _34194_ (.A1(_13200_),
    .A2(_03035_),
    .B1(_03029_),
    .Y(_13201_));
 sky130_fd_sc_hd__nand2_1 _34195_ (.A(_13199_),
    .B(_13201_),
    .Y(_13202_));
 sky130_fd_sc_hd__nand2_1 _34196_ (.A(_13052_),
    .B(_13043_),
    .Y(_13203_));
 sky130_fd_sc_hd__nand2_1 _34197_ (.A(_13203_),
    .B(_13055_),
    .Y(_13204_));
 sky130_fd_sc_hd__nand2_1 _34198_ (.A(_03027_),
    .B(_03033_),
    .Y(_13205_));
 sky130_fd_sc_hd__nor2_1 _34199_ (.A(_13054_),
    .B(_13205_),
    .Y(_13206_));
 sky130_fd_sc_hd__nand2_1 _34200_ (.A(_03027_),
    .B(_03032_),
    .Y(_13207_));
 sky130_fd_sc_hd__inv_1 _34201_ (.A(_03026_),
    .Y(_13208_));
 sky130_fd_sc_hd__nand2_1 _34202_ (.A(_13207_),
    .B(_13208_),
    .Y(_13209_));
 sky130_fd_sc_hd__o21bai_1 _34203_ (.A1(_13205_),
    .A2(_13056_),
    .B1_N(_13209_),
    .Y(_13210_));
 sky130_fd_sc_hd__a21oi_1 _34204_ (.A1(_13204_),
    .A2(_13206_),
    .B1(_13210_),
    .Y(_13211_));
 sky130_fd_sc_hd__nand4_1 _34205_ (.A(_13047_),
    .B(_13049_),
    .C(_13043_),
    .D(_13206_),
    .Y(_13212_));
 sky130_fd_sc_hd__nand2_1 _34206_ (.A(_13211_),
    .B(_13212_),
    .Y(_13213_));
 sky130_fd_sc_hd__nand2_1 _34207_ (.A(_13213_),
    .B(net2868),
    .Y(_13214_));
 sky130_fd_sc_hd__o21ai_0 _34208_ (.A1(net2868),
    .A2(_13202_),
    .B1(_13214_),
    .Y(_13215_));
 sky130_fd_sc_hd__xor2_4 _34209_ (.A(_03022_),
    .B(_13215_),
    .X(_13216_));
 sky130_fd_sc_hd__inv_1 _34210_ (.A(_13216_),
    .Y(_13217_));
 sky130_fd_sc_hd__o21ai_0 _34211_ (.A1(net2846),
    .A2(_13217_),
    .B1(_20766_),
    .Y(_13218_));
 sky130_fd_sc_hd__nand2_1 _34212_ (.A(_13218_),
    .B(net2017),
    .Y(_13219_));
 sky130_fd_sc_hd__nand2_1 _34213_ (.A(net1796),
    .B(_03173_),
    .Y(_13220_));
 sky130_fd_sc_hd__nand2_1 _34214_ (.A(net1869),
    .B(_03172_),
    .Y(_13221_));
 sky130_fd_sc_hd__o211ai_1 _34215_ (.A1(_03176_),
    .A2(net1230),
    .B1(_13220_),
    .C1(_13221_),
    .Y(_13222_));
 sky130_fd_sc_hd__a21oi_1 _34217_ (.A1(_13222_),
    .A2(net2861),
    .B1(net2853),
    .Y(_13224_));
 sky130_fd_sc_hd__nand3_1 _34218_ (.A(_13035_),
    .B(\inst$top.soc.cpu.sink__payload$12[11] ),
    .C(\inst$top.soc.cpu.sink__payload$12[10] ),
    .Y(_13225_));
 sky130_fd_sc_hd__o21ai_0 _34219_ (.A1(\inst$top.soc.cpu.sink__payload$12[12] ),
    .A2(_13225_),
    .B1(net2851),
    .Y(_13226_));
 sky130_fd_sc_hd__a21oi_1 _34220_ (.A1(\inst$top.soc.cpu.sink__payload$12[12] ),
    .A2(_13225_),
    .B1(_13226_),
    .Y(_13227_));
 sky130_fd_sc_hd__a21oi_4 _34221_ (.A1(_13219_),
    .A2(_13224_),
    .B1(_13227_),
    .Y(_13228_));
 sky130_fd_sc_hd__inv_1 _34222_ (.A(\inst$top.soc.cpu.sink__payload$18[121] ),
    .Y(_13229_));
 sky130_fd_sc_hd__nor2_1 _34224_ (.A(\inst$top.soc.cpu.shifter.m_result$7[12] ),
    .B(net2003),
    .Y(_13231_));
 sky130_fd_sc_hd__o21ai_0 _34225_ (.A1(net2872),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[19] ),
    .B1(net2837),
    .Y(_13232_));
 sky130_fd_sc_hd__o22ai_1 _34226_ (.A1(_13229_),
    .A2(net2837),
    .B1(_13231_),
    .B2(_13232_),
    .Y(_13233_));
 sky130_fd_sc_hd__nand2_1 _34228_ (.A(_13233_),
    .B(net2015),
    .Y(_13235_));
 sky130_fd_sc_hd__a21oi_1 _34229_ (.A1(_10400_),
    .A2(net2916),
    .B1(net2009),
    .Y(_13236_));
 sky130_fd_sc_hd__o21ai_2 _34230_ (.A1(net2916),
    .A2(\inst$top.soc.cpu.divider.quotient[12] ),
    .B1(_13236_),
    .Y(_13237_));
 sky130_fd_sc_hd__a21oi_1 _34231_ (.A1(_13235_),
    .A2(net1794),
    .B1(net2831),
    .Y(_13238_));
 sky130_fd_sc_hd__inv_1 _34232_ (.A(_13238_),
    .Y(_13239_));
 sky130_fd_sc_hd__inv_1 _34233_ (.A(net988),
    .Y(_13240_));
 sky130_fd_sc_hd__o22ai_1 _34234_ (.A1(_13239_),
    .A2(net785),
    .B1(_13240_),
    .B2(_12956_),
    .Y(_13241_));
 sky130_fd_sc_hd__a21oi_1 _34235_ (.A1(_12959_),
    .A2(_13228_),
    .B1(_13241_),
    .Y(_13242_));
 sky130_fd_sc_hd__nand2_1 _34236_ (.A(net713),
    .B(_13242_),
    .Y(_13243_));
 sky130_fd_sc_hd__nand2_1 _34237_ (.A(_13243_),
    .B(net2173),
    .Y(_13244_));
 sky130_fd_sc_hd__nor2_2 _34238_ (.A(_13196_),
    .B(_13244_),
    .Y(_04187_));
 sky130_fd_sc_hd__nor2_1 _34239_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[13] ),
    .B(net710),
    .Y(_13245_));
 sky130_fd_sc_hd__inv_1 _34240_ (.A(\inst$top.soc.cpu.sink__payload$18[122] ),
    .Y(_13246_));
 sky130_fd_sc_hd__nor2_1 _34241_ (.A(\inst$top.soc.cpu.shifter.m_result$7[13] ),
    .B(net2004),
    .Y(_13247_));
 sky130_fd_sc_hd__o21ai_0 _34242_ (.A1(net2873),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[18] ),
    .B1(net2836),
    .Y(_13248_));
 sky130_fd_sc_hd__o22ai_1 _34243_ (.A1(_13246_),
    .A2(net2836),
    .B1(_13247_),
    .B2(_13248_),
    .Y(_13249_));
 sky130_fd_sc_hd__nand2_1 _34245_ (.A(_13249_),
    .B(net2015),
    .Y(_13251_));
 sky130_fd_sc_hd__a21oi_1 _34246_ (.A1(_10411_),
    .A2(net2916),
    .B1(net2009),
    .Y(_13252_));
 sky130_fd_sc_hd__o21ai_2 _34247_ (.A1(net2916),
    .A2(\inst$top.soc.cpu.divider.quotient[13] ),
    .B1(_13252_),
    .Y(_13253_));
 sky130_fd_sc_hd__a21oi_1 _34248_ (.A1(_13251_),
    .A2(net1793),
    .B1(net2830),
    .Y(_13254_));
 sky130_fd_sc_hd__inv_1 _34249_ (.A(_13254_),
    .Y(_13255_));
 sky130_fd_sc_hd__o21bai_1 _34251_ (.A1(_00169_),
    .A2(_13174_),
    .B1_N(_13159_),
    .Y(_13257_));
 sky130_fd_sc_hd__nand2_1 _34252_ (.A(_13257_),
    .B(_13161_),
    .Y(_13258_));
 sky130_fd_sc_hd__nand2_1 _34253_ (.A(_13258_),
    .B(_13163_),
    .Y(_13259_));
 sky130_fd_sc_hd__nand2_1 _34254_ (.A(_03022_),
    .B(_03027_),
    .Y(_13260_));
 sky130_fd_sc_hd__nor2_1 _34255_ (.A(_13180_),
    .B(_13260_),
    .Y(_13261_));
 sky130_fd_sc_hd__inv_1 _34256_ (.A(_13261_),
    .Y(_13262_));
 sky130_fd_sc_hd__nor2_1 _34257_ (.A(_13175_),
    .B(_13262_),
    .Y(_13263_));
 sky130_fd_sc_hd__a21oi_1 _34258_ (.A1(_03022_),
    .A2(_03026_),
    .B1(_03021_),
    .Y(_13264_));
 sky130_fd_sc_hd__o21ai_0 _34259_ (.A1(_13260_),
    .A2(_13183_),
    .B1(_13264_),
    .Y(_13265_));
 sky130_fd_sc_hd__o21bai_1 _34260_ (.A1(_13262_),
    .A2(_13173_),
    .B1_N(_13265_),
    .Y(_13266_));
 sky130_fd_sc_hd__a21o_1 _34261_ (.A1(_13259_),
    .A2(_13263_),
    .B1(_13266_),
    .X(_13267_));
 sky130_fd_sc_hd__nor2_1 _34262_ (.A(_03022_),
    .B(_03027_),
    .Y(_13268_));
 sky130_fd_sc_hd__nand2_1 _34263_ (.A(_13158_),
    .B(_13268_),
    .Y(_13269_));
 sky130_fd_sc_hd__inv_1 _34264_ (.A(_03022_),
    .Y(_13270_));
 sky130_fd_sc_hd__a21oi_1 _34265_ (.A1(_13270_),
    .A2(_03029_),
    .B1(_00826_),
    .Y(_13271_));
 sky130_fd_sc_hd__nand2_1 _34266_ (.A(_13269_),
    .B(_13271_),
    .Y(_13272_));
 sky130_fd_sc_hd__nand2_1 _34267_ (.A(_13272_),
    .B(net2006),
    .Y(_13273_));
 sky130_fd_sc_hd__o21ai_0 _34268_ (.A1(net2006),
    .A2(_13267_),
    .B1(_13273_),
    .Y(_13274_));
 sky130_fd_sc_hd__inv_1 _34269_ (.A(_13274_),
    .Y(_13275_));
 sky130_fd_sc_hd__inv_1 _34270_ (.A(_03016_),
    .Y(_13276_));
 sky130_fd_sc_hd__nand2_1 _34271_ (.A(_13275_),
    .B(_13276_),
    .Y(_13277_));
 sky130_fd_sc_hd__nand2_1 _34272_ (.A(_13274_),
    .B(_03016_),
    .Y(_13278_));
 sky130_fd_sc_hd__nand3_1 _34273_ (.A(_13277_),
    .B(net2214),
    .C(_13278_),
    .Y(_13279_));
 sky130_fd_sc_hd__nand2_1 _34274_ (.A(_13279_),
    .B(_20785_),
    .Y(_13280_));
 sky130_fd_sc_hd__nand2_1 _34275_ (.A(_13280_),
    .B(net2019),
    .Y(_13281_));
 sky130_fd_sc_hd__nand2_1 _34276_ (.A(net1795),
    .B(_03180_),
    .Y(_13282_));
 sky130_fd_sc_hd__nand2_1 _34277_ (.A(net1868),
    .B(_03179_),
    .Y(_13283_));
 sky130_fd_sc_hd__o211ai_1 _34278_ (.A1(_03183_),
    .A2(net1229),
    .B1(_13282_),
    .C1(_13283_),
    .Y(_13284_));
 sky130_fd_sc_hd__a21oi_1 _34280_ (.A1(_13284_),
    .A2(net2863),
    .B1(net2855),
    .Y(_13286_));
 sky130_fd_sc_hd__nor4_1 _34281_ (.A(_20751_),
    .B(_20726_),
    .C(_20705_),
    .D(_20685_),
    .Y(_13287_));
 sky130_fd_sc_hd__inv_1 _34282_ (.A(_13117_),
    .Y(_13288_));
 sky130_fd_sc_hd__nor2_1 _34283_ (.A(_13114_),
    .B(_13288_),
    .Y(_13289_));
 sky130_fd_sc_hd__nand2_1 _34284_ (.A(_13287_),
    .B(_13289_),
    .Y(_13290_));
 sky130_fd_sc_hd__inv_1 _34285_ (.A(_13290_),
    .Y(_13291_));
 sky130_fd_sc_hd__nand2_1 _34286_ (.A(_13291_),
    .B(_20771_),
    .Y(_13292_));
 sky130_fd_sc_hd__nand2_1 _34287_ (.A(_13290_),
    .B(\inst$top.soc.cpu.sink__payload$12[13] ),
    .Y(_13293_));
 sky130_fd_sc_hd__nand3_1 _34288_ (.A(_13292_),
    .B(net2851),
    .C(_13293_),
    .Y(_13294_));
 sky130_fd_sc_hd__a21boi_1 _34289_ (.A1(_13281_),
    .A2(_13286_),
    .B1_N(_13294_),
    .Y(_13295_));
 sky130_fd_sc_hd__nand2_1 _34290_ (.A(net602),
    .B(net787),
    .Y(_13296_));
 sky130_fd_sc_hd__o21ai_0 _34291_ (.A1(net784),
    .A2(_13255_),
    .B1(_13296_),
    .Y(_13297_));
 sky130_fd_sc_hd__a21oi_1 _34292_ (.A1(net738),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[13] ),
    .B1(_13297_),
    .Y(_13298_));
 sky130_fd_sc_hd__nand2_1 _34293_ (.A(net709),
    .B(_13298_),
    .Y(_13299_));
 sky130_fd_sc_hd__nand2_1 _34294_ (.A(_13299_),
    .B(net2156),
    .Y(_13300_));
 sky130_fd_sc_hd__nor2_2 _34295_ (.A(_13245_),
    .B(_13300_),
    .Y(_04188_));
 sky130_fd_sc_hd__nor2_1 _34296_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[14] ),
    .B(net710),
    .Y(_13301_));
 sky130_fd_sc_hd__nor2_1 _34298_ (.A(_03022_),
    .B(_13276_),
    .Y(_13303_));
 sky130_fd_sc_hd__nand2_1 _34299_ (.A(_13202_),
    .B(_13303_),
    .Y(_13304_));
 sky130_fd_sc_hd__inv_1 _34300_ (.A(_00826_),
    .Y(_13305_));
 sky130_fd_sc_hd__o21ai_0 _34301_ (.A1(_13305_),
    .A2(_13276_),
    .B1(_00940_),
    .Y(_13306_));
 sky130_fd_sc_hd__inv_1 _34302_ (.A(_13306_),
    .Y(_13307_));
 sky130_fd_sc_hd__nand2_1 _34303_ (.A(_13304_),
    .B(_13307_),
    .Y(_13308_));
 sky130_fd_sc_hd__nand2_1 _34305_ (.A(_13308_),
    .B(net2008),
    .Y(_13310_));
 sky130_fd_sc_hd__nor2_1 _34306_ (.A(_03016_),
    .B(_13270_),
    .Y(_13311_));
 sky130_fd_sc_hd__inv_1 _34307_ (.A(_13311_),
    .Y(_13312_));
 sky130_fd_sc_hd__nor2_1 _34308_ (.A(_13205_),
    .B(_13312_),
    .Y(_13313_));
 sky130_fd_sc_hd__a21o_1 _34309_ (.A1(_13276_),
    .A2(_03021_),
    .B1(_03018_),
    .X(_13314_));
 sky130_fd_sc_hd__a21oi_1 _34310_ (.A1(_13209_),
    .A2(_13311_),
    .B1(_13314_),
    .Y(_13315_));
 sky130_fd_sc_hd__a21boi_0 _34311_ (.A1(_13057_),
    .A2(_13313_),
    .B1_N(_13315_),
    .Y(_13316_));
 sky130_fd_sc_hd__inv_1 _34312_ (.A(_13053_),
    .Y(_13317_));
 sky130_fd_sc_hd__inv_1 _34313_ (.A(_13313_),
    .Y(_13318_));
 sky130_fd_sc_hd__nor2_1 _34314_ (.A(_13044_),
    .B(_13318_),
    .Y(_13319_));
 sky130_fd_sc_hd__nand2_1 _34315_ (.A(_13317_),
    .B(_13319_),
    .Y(_13320_));
 sky130_fd_sc_hd__nand3_1 _34317_ (.A(_13316_),
    .B(_13320_),
    .C(\inst$top.soc.cpu.adder$307.x_sub ),
    .Y(_13322_));
 sky130_fd_sc_hd__nand2_1 _34318_ (.A(_13310_),
    .B(_13322_),
    .Y(_13323_));
 sky130_fd_sc_hd__nand2_1 _34319_ (.A(_13323_),
    .B(_03010_),
    .Y(_13324_));
 sky130_fd_sc_hd__inv_1 _34320_ (.A(_03010_),
    .Y(_13325_));
 sky130_fd_sc_hd__nand3_1 _34321_ (.A(_13310_),
    .B(_13325_),
    .C(_13322_),
    .Y(_13326_));
 sky130_fd_sc_hd__nand2_2 _34322_ (.A(_13324_),
    .B(_13326_),
    .Y(_13327_));
 sky130_fd_sc_hd__o21ai_0 _34323_ (.A1(net2846),
    .A2(_13327_),
    .B1(_20803_),
    .Y(_13328_));
 sky130_fd_sc_hd__nand2_1 _34324_ (.A(_13328_),
    .B(net2017),
    .Y(_13329_));
 sky130_fd_sc_hd__nand2_1 _34325_ (.A(net1795),
    .B(_03187_),
    .Y(_13330_));
 sky130_fd_sc_hd__nand2_1 _34326_ (.A(net1868),
    .B(_03186_),
    .Y(_13331_));
 sky130_fd_sc_hd__o211ai_1 _34327_ (.A1(_03190_),
    .A2(net1229),
    .B1(_13330_),
    .C1(_13331_),
    .Y(_13332_));
 sky130_fd_sc_hd__a21oi_1 _34328_ (.A1(_13332_),
    .A2(net2861),
    .B1(net2851),
    .Y(_13333_));
 sky130_fd_sc_hd__nand2_1 _34329_ (.A(\inst$top.soc.cpu.sink__payload$12[13] ),
    .B(\inst$top.soc.cpu.sink__payload$12[12] ),
    .Y(_13334_));
 sky130_fd_sc_hd__nor2_1 _34330_ (.A(_13334_),
    .B(_13225_),
    .Y(_13335_));
 sky130_fd_sc_hd__a21oi_1 _34331_ (.A1(_13335_),
    .A2(_20789_),
    .B1(net2001),
    .Y(_13336_));
 sky130_fd_sc_hd__o21ai_0 _34332_ (.A1(_20789_),
    .A2(_13335_),
    .B1(_13336_),
    .Y(_13337_));
 sky130_fd_sc_hd__a21boi_1 _34333_ (.A1(_13329_),
    .A2(_13333_),
    .B1_N(_13337_),
    .Y(_13338_));
 sky130_fd_sc_hd__inv_1 _34334_ (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[14] ),
    .Y(_13339_));
 sky130_fd_sc_hd__inv_1 _34335_ (.A(\inst$top.soc.cpu.sink__payload$18[123] ),
    .Y(_13340_));
 sky130_fd_sc_hd__nor2_1 _34337_ (.A(\inst$top.soc.cpu.shifter.m_result$7[14] ),
    .B(net2003),
    .Y(_13342_));
 sky130_fd_sc_hd__o21ai_0 _34338_ (.A1(net2871),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[17] ),
    .B1(net2840),
    .Y(_13343_));
 sky130_fd_sc_hd__o22ai_1 _34339_ (.A1(_13340_),
    .A2(net2840),
    .B1(_13342_),
    .B2(_13343_),
    .Y(_13344_));
 sky130_fd_sc_hd__nand2_1 _34340_ (.A(_13344_),
    .B(net2015),
    .Y(_13345_));
 sky130_fd_sc_hd__a21oi_1 _34341_ (.A1(_10440_),
    .A2(net2916),
    .B1(net2009),
    .Y(_13346_));
 sky130_fd_sc_hd__o21ai_2 _34342_ (.A1(net2916),
    .A2(\inst$top.soc.cpu.divider.quotient[14] ),
    .B1(_13346_),
    .Y(_13347_));
 sky130_fd_sc_hd__a21oi_1 _34343_ (.A1(_13345_),
    .A2(net1792),
    .B1(net2831),
    .Y(_13348_));
 sky130_fd_sc_hd__nand2_1 _34344_ (.A(_12984_),
    .B(_13348_),
    .Y(_13349_));
 sky130_fd_sc_hd__o21ai_0 _34345_ (.A1(_13339_),
    .A2(_12956_),
    .B1(_13349_),
    .Y(_13350_));
 sky130_fd_sc_hd__a21oi_1 _34346_ (.A1(net786),
    .A2(net604),
    .B1(_13350_),
    .Y(_13351_));
 sky130_fd_sc_hd__nand2_1 _34347_ (.A(net710),
    .B(_13351_),
    .Y(_13352_));
 sky130_fd_sc_hd__nand2_1 _34348_ (.A(_13352_),
    .B(net2171),
    .Y(_13353_));
 sky130_fd_sc_hd__nor2_2 _34349_ (.A(_13301_),
    .B(_13353_),
    .Y(_04189_));
 sky130_fd_sc_hd__nor2_1 _34350_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[15] ),
    .B(net709),
    .Y(_13354_));
 sky130_fd_sc_hd__nand3_1 _34351_ (.A(_13272_),
    .B(_03010_),
    .C(_03016_),
    .Y(_13355_));
 sky130_fd_sc_hd__a21oi_1 _34353_ (.A1(_03015_),
    .A2(_03010_),
    .B1(_03009_),
    .Y(_13357_));
 sky130_fd_sc_hd__nand3_1 _34354_ (.A(_13355_),
    .B(net2008),
    .C(_13357_),
    .Y(_13358_));
 sky130_fd_sc_hd__nor2_1 _34355_ (.A(_03010_),
    .B(_03016_),
    .Y(_13359_));
 sky130_fd_sc_hd__nand2_1 _34356_ (.A(_13267_),
    .B(_13359_),
    .Y(_13360_));
 sky130_fd_sc_hd__a21oi_1 _34357_ (.A1(_13325_),
    .A2(_03018_),
    .B1(_03012_),
    .Y(_13361_));
 sky130_fd_sc_hd__nand2_1 _34358_ (.A(_13360_),
    .B(_13361_),
    .Y(_13362_));
 sky130_fd_sc_hd__nand2_1 _34360_ (.A(_13362_),
    .B(\inst$top.soc.cpu.adder$307.x_sub ),
    .Y(_13364_));
 sky130_fd_sc_hd__nand2_1 _34361_ (.A(_13358_),
    .B(_13364_),
    .Y(_13365_));
 sky130_fd_sc_hd__inv_1 _34362_ (.A(_03004_),
    .Y(_13366_));
 sky130_fd_sc_hd__nand2_1 _34363_ (.A(_13365_),
    .B(_13366_),
    .Y(_13367_));
 sky130_fd_sc_hd__nand3_1 _34364_ (.A(_13358_),
    .B(_03004_),
    .C(_13364_),
    .Y(_13368_));
 sky130_fd_sc_hd__nand2_1 _34365_ (.A(_13367_),
    .B(_13368_),
    .Y(_13369_));
 sky130_fd_sc_hd__nand2_1 _34366_ (.A(_13369_),
    .B(net2215),
    .Y(_13370_));
 sky130_fd_sc_hd__nand2_1 _34367_ (.A(_13370_),
    .B(_20824_),
    .Y(_13371_));
 sky130_fd_sc_hd__nand2_1 _34369_ (.A(_13371_),
    .B(net2017),
    .Y(_13373_));
 sky130_fd_sc_hd__nand2_1 _34372_ (.A(net1796),
    .B(_03194_),
    .Y(_13376_));
 sky130_fd_sc_hd__nand2_1 _34374_ (.A(net1869),
    .B(_03193_),
    .Y(_13378_));
 sky130_fd_sc_hd__o211ai_1 _34375_ (.A1(_03197_),
    .A2(net1230),
    .B1(_13376_),
    .C1(_13378_),
    .Y(_13379_));
 sky130_fd_sc_hd__a21oi_1 _34378_ (.A1(_13379_),
    .A2(net2861),
    .B1(net2851),
    .Y(_13382_));
 sky130_fd_sc_hd__nor4_1 _34379_ (.A(_20789_),
    .B(_20771_),
    .C(_20751_),
    .D(_20726_),
    .Y(_13383_));
 sky130_fd_sc_hd__nand3_1 _34380_ (.A(_13383_),
    .B(_13117_),
    .C(_13115_),
    .Y(_13384_));
 sky130_fd_sc_hd__o21ai_0 _34381_ (.A1(\inst$top.soc.cpu.sink__payload$12[15] ),
    .A2(_13384_),
    .B1(net2851),
    .Y(_13385_));
 sky130_fd_sc_hd__a21oi_1 _34382_ (.A1(\inst$top.soc.cpu.sink__payload$12[15] ),
    .A2(_13384_),
    .B1(_13385_),
    .Y(_13386_));
 sky130_fd_sc_hd__a21oi_2 _34383_ (.A1(_13373_),
    .A2(_13382_),
    .B1(_13386_),
    .Y(_13387_));
 sky130_fd_sc_hd__inv_1 _34384_ (.A(\inst$top.soc.cpu.sink__payload$18[124] ),
    .Y(_13388_));
 sky130_fd_sc_hd__nor2_1 _34385_ (.A(\inst$top.soc.cpu.shifter.m_result$7[15] ),
    .B(net2002),
    .Y(_13389_));
 sky130_fd_sc_hd__o21ai_0 _34386_ (.A1(net2869),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[16] ),
    .B1(net2836),
    .Y(_13390_));
 sky130_fd_sc_hd__o22ai_1 _34387_ (.A1(_13388_),
    .A2(net2835),
    .B1(_13389_),
    .B2(_13390_),
    .Y(_13391_));
 sky130_fd_sc_hd__nand2_1 _34388_ (.A(_13391_),
    .B(net2014),
    .Y(_13392_));
 sky130_fd_sc_hd__a21oi_1 _34389_ (.A1(_10460_),
    .A2(net2918),
    .B1(net2009),
    .Y(_13393_));
 sky130_fd_sc_hd__o21ai_4 _34390_ (.A1(net2918),
    .A2(\inst$top.soc.cpu.divider.quotient[15] ),
    .B1(_13393_),
    .Y(_13394_));
 sky130_fd_sc_hd__a21oi_1 _34391_ (.A1(_13392_),
    .A2(_13394_),
    .B1(net2830),
    .Y(_13395_));
 sky130_fd_sc_hd__inv_1 _34392_ (.A(_13395_),
    .Y(_13396_));
 sky130_fd_sc_hd__o22ai_1 _34393_ (.A1(_13396_),
    .A2(net784),
    .B1(_05597_),
    .B2(_12956_),
    .Y(_13397_));
 sky130_fd_sc_hd__a21oi_1 _34394_ (.A1(net787),
    .A2(_13387_),
    .B1(_13397_),
    .Y(_13398_));
 sky130_fd_sc_hd__nand2_1 _34395_ (.A(net709),
    .B(_13398_),
    .Y(_13399_));
 sky130_fd_sc_hd__nand2_1 _34396_ (.A(_13399_),
    .B(net2156),
    .Y(_13400_));
 sky130_fd_sc_hd__nor2_2 _34397_ (.A(_13354_),
    .B(_13400_),
    .Y(_04190_));
 sky130_fd_sc_hd__nor2_1 _34398_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[16] ),
    .B(net709),
    .Y(_13401_));
 sky130_fd_sc_hd__inv_1 _34399_ (.A(\inst$top.soc.cpu.sink__payload$18[125] ),
    .Y(_13402_));
 sky130_fd_sc_hd__nor2_1 _34400_ (.A(net2833),
    .B(_13402_),
    .Y(_13403_));
 sky130_fd_sc_hd__inv_1 _34401_ (.A(\inst$top.soc.cpu.shifter.m_result$7[16] ),
    .Y(_13404_));
 sky130_fd_sc_hd__o21ai_0 _34402_ (.A1(net2869),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[15] ),
    .B1(net2836),
    .Y(_13405_));
 sky130_fd_sc_hd__a21oi_1 _34403_ (.A1(net2869),
    .A2(_13404_),
    .B1(_13405_),
    .Y(_13406_));
 sky130_fd_sc_hd__o21ai_0 _34404_ (.A1(_13403_),
    .A2(_13406_),
    .B1(net2013),
    .Y(_13407_));
 sky130_fd_sc_hd__a21oi_1 _34405_ (.A1(_10484_),
    .A2(net2918),
    .B1(net2009),
    .Y(_13408_));
 sky130_fd_sc_hd__o21ai_4 _34406_ (.A1(net2918),
    .A2(\inst$top.soc.cpu.divider.quotient[16] ),
    .B1(_13408_),
    .Y(_13409_));
 sky130_fd_sc_hd__a21oi_1 _34407_ (.A1(_13407_),
    .A2(_13409_),
    .B1(net2829),
    .Y(_13410_));
 sky130_fd_sc_hd__inv_1 _34408_ (.A(_13410_),
    .Y(_13411_));
 sky130_fd_sc_hd__inv_1 _34409_ (.A(_13067_),
    .Y(_13412_));
 sky130_fd_sc_hd__nand3_1 _34410_ (.A(_13061_),
    .B(_13071_),
    .C(_13074_),
    .Y(_13413_));
 sky130_fd_sc_hd__nand2_1 _34411_ (.A(_13062_),
    .B(_13413_),
    .Y(_13414_));
 sky130_fd_sc_hd__inv_1 _34412_ (.A(_13064_),
    .Y(_13415_));
 sky130_fd_sc_hd__a21oi_1 _34413_ (.A1(_13414_),
    .A2(_13059_),
    .B1(_13415_),
    .Y(_13416_));
 sky130_fd_sc_hd__o21bai_1 _34414_ (.A1(_13412_),
    .A2(_13416_),
    .B1_N(_13077_),
    .Y(_13417_));
 sky130_fd_sc_hd__nand2_1 _34415_ (.A(_13066_),
    .B(_13198_),
    .Y(_13418_));
 sky130_fd_sc_hd__inv_1 _34416_ (.A(_13303_),
    .Y(_13419_));
 sky130_fd_sc_hd__nor2_1 _34417_ (.A(_03004_),
    .B(_13325_),
    .Y(_13420_));
 sky130_fd_sc_hd__inv_1 _34418_ (.A(_13420_),
    .Y(_13421_));
 sky130_fd_sc_hd__nor2_1 _34419_ (.A(_13419_),
    .B(_13421_),
    .Y(_13422_));
 sky130_fd_sc_hd__inv_1 _34420_ (.A(_13422_),
    .Y(_13423_));
 sky130_fd_sc_hd__nor2_1 _34421_ (.A(_13418_),
    .B(_13423_),
    .Y(_13424_));
 sky130_fd_sc_hd__a21boi_0 _34422_ (.A1(_13078_),
    .A2(_13198_),
    .B1_N(_13201_),
    .Y(_13425_));
 sky130_fd_sc_hd__o21ai_0 _34423_ (.A1(_03004_),
    .A2(_01062_),
    .B1(_01185_),
    .Y(_13426_));
 sky130_fd_sc_hd__a21oi_1 _34424_ (.A1(_13306_),
    .A2(_13420_),
    .B1(_13426_),
    .Y(_13427_));
 sky130_fd_sc_hd__o21ai_0 _34425_ (.A1(_13423_),
    .A2(_13425_),
    .B1(_13427_),
    .Y(_13428_));
 sky130_fd_sc_hd__a21oi_1 _34426_ (.A1(_13417_),
    .A2(_13424_),
    .B1(_13428_),
    .Y(_13429_));
 sky130_fd_sc_hd__nand2_1 _34427_ (.A(_13429_),
    .B(net2008),
    .Y(_13430_));
 sky130_fd_sc_hd__o21ai_0 _34428_ (.A1(_13042_),
    .A2(_13053_),
    .B1(_13055_),
    .Y(_13431_));
 sky130_fd_sc_hd__nor2_1 _34429_ (.A(_03010_),
    .B(_13366_),
    .Y(_13432_));
 sky130_fd_sc_hd__inv_1 _34430_ (.A(_13432_),
    .Y(_13433_));
 sky130_fd_sc_hd__nor2_1 _34431_ (.A(_13312_),
    .B(_13433_),
    .Y(_13434_));
 sky130_fd_sc_hd__inv_1 _34432_ (.A(_13434_),
    .Y(_13435_));
 sky130_fd_sc_hd__nor3_1 _34433_ (.A(_13054_),
    .B(_13205_),
    .C(_13435_),
    .Y(_13436_));
 sky130_fd_sc_hd__nand2_1 _34434_ (.A(_13431_),
    .B(_13436_),
    .Y(_13437_));
 sky130_fd_sc_hd__nand2_1 _34435_ (.A(_13314_),
    .B(_13432_),
    .Y(_13438_));
 sky130_fd_sc_hd__a21oi_1 _34436_ (.A1(_03004_),
    .A2(_03012_),
    .B1(_03003_),
    .Y(_13439_));
 sky130_fd_sc_hd__nand2_1 _34437_ (.A(_13438_),
    .B(_13439_),
    .Y(_13440_));
 sky130_fd_sc_hd__a21oi_1 _34438_ (.A1(_13210_),
    .A2(_13434_),
    .B1(_13440_),
    .Y(_13441_));
 sky130_fd_sc_hd__nand2_1 _34439_ (.A(_13437_),
    .B(_13441_),
    .Y(_13442_));
 sky130_fd_sc_hd__nand2_1 _34440_ (.A(_13442_),
    .B(net2868),
    .Y(_13443_));
 sky130_fd_sc_hd__nand2_1 _34441_ (.A(_13430_),
    .B(_13443_),
    .Y(_13444_));
 sky130_fd_sc_hd__nand2_1 _34442_ (.A(_13444_),
    .B(_02998_),
    .Y(_13445_));
 sky130_fd_sc_hd__inv_1 _34443_ (.A(_02998_),
    .Y(_13446_));
 sky130_fd_sc_hd__nand3_1 _34444_ (.A(_13430_),
    .B(_13446_),
    .C(_13443_),
    .Y(_13447_));
 sky130_fd_sc_hd__nand2_2 _34445_ (.A(_13445_),
    .B(_13447_),
    .Y(_13448_));
 sky130_fd_sc_hd__o21ai_0 _34446_ (.A1(net2848),
    .A2(_13448_),
    .B1(net3045),
    .Y(_13449_));
 sky130_fd_sc_hd__nand2_1 _34447_ (.A(net1797),
    .B(_03201_),
    .Y(_13450_));
 sky130_fd_sc_hd__nand2_1 _34448_ (.A(net1870),
    .B(_03200_),
    .Y(_13451_));
 sky130_fd_sc_hd__o211ai_1 _34449_ (.A1(_03204_),
    .A2(net1232),
    .B1(_13450_),
    .C1(_13451_),
    .Y(_13452_));
 sky130_fd_sc_hd__nor2_1 _34450_ (.A(net2019),
    .B(_13452_),
    .Y(_13453_));
 sky130_fd_sc_hd__nor2_1 _34451_ (.A(net2855),
    .B(_13453_),
    .Y(_13454_));
 sky130_fd_sc_hd__o21ai_0 _34452_ (.A1(net2863),
    .A2(_13449_),
    .B1(_13454_),
    .Y(_13455_));
 sky130_fd_sc_hd__nor3_1 _34453_ (.A(_20807_),
    .B(_20789_),
    .C(_13334_),
    .Y(_13456_));
 sky130_fd_sc_hd__nor3_1 _34454_ (.A(_20726_),
    .B(_20705_),
    .C(_13030_),
    .Y(_13457_));
 sky130_fd_sc_hd__nand2_1 _34455_ (.A(_13456_),
    .B(_13457_),
    .Y(_13458_));
 sky130_fd_sc_hd__o21ai_0 _34456_ (.A1(_13034_),
    .A2(_13458_),
    .B1(_05598_),
    .Y(_13459_));
 sky130_fd_sc_hd__nand4_1 _34457_ (.A(_13033_),
    .B(_13456_),
    .C(\inst$top.soc.cpu.sink__payload$12[16] ),
    .D(_13457_),
    .Y(_13460_));
 sky130_fd_sc_hd__nand3_1 _34458_ (.A(_13459_),
    .B(_13460_),
    .C(net2853),
    .Y(_13461_));
 sky130_fd_sc_hd__nand2_1 _34459_ (.A(_13455_),
    .B(_13461_),
    .Y(_13462_));
 sky130_fd_sc_hd__nand2_1 _34460_ (.A(_13462_),
    .B(net787),
    .Y(_13463_));
 sky130_fd_sc_hd__o21ai_0 _34461_ (.A1(net785),
    .A2(_13411_),
    .B1(_13463_),
    .Y(_13464_));
 sky130_fd_sc_hd__a21oi_1 _34462_ (.A1(net738),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[16] ),
    .B1(_13464_),
    .Y(_13465_));
 sky130_fd_sc_hd__nand2_1 _34463_ (.A(net710),
    .B(_13465_),
    .Y(_13466_));
 sky130_fd_sc_hd__nand2_1 _34464_ (.A(_13466_),
    .B(net2177),
    .Y(_13467_));
 sky130_fd_sc_hd__nor2_2 _34465_ (.A(_13401_),
    .B(_13467_),
    .Y(_04191_));
 sky130_fd_sc_hd__nor2_1 _34466_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[17] ),
    .B(net713),
    .Y(_13468_));
 sky130_fd_sc_hd__nand3_1 _34467_ (.A(_13119_),
    .B(\inst$top.soc.cpu.sink__payload$12[16] ),
    .C(_13456_),
    .Y(_13469_));
 sky130_fd_sc_hd__a21oi_1 _34468_ (.A1(_13469_),
    .A2(\inst$top.soc.cpu.sink__payload$12[17] ),
    .B1(net2001),
    .Y(_13470_));
 sky130_fd_sc_hd__o21ai_0 _34469_ (.A1(\inst$top.soc.cpu.sink__payload$12[17] ),
    .A2(_13469_),
    .B1(_13470_),
    .Y(_13471_));
 sky130_fd_sc_hd__inv_1 _34470_ (.A(_13471_),
    .Y(_13472_));
 sky130_fd_sc_hd__inv_1 _34471_ (.A(_02993_),
    .Y(_13473_));
 sky130_fd_sc_hd__nand2_1 _34472_ (.A(_13169_),
    .B(_13173_),
    .Y(_13474_));
 sky130_fd_sc_hd__nand2_1 _34473_ (.A(_02998_),
    .B(_03004_),
    .Y(_13475_));
 sky130_fd_sc_hd__inv_1 _34474_ (.A(_13359_),
    .Y(_13476_));
 sky130_fd_sc_hd__nor2_1 _34475_ (.A(_13475_),
    .B(_13476_),
    .Y(_13477_));
 sky130_fd_sc_hd__inv_1 _34476_ (.A(_13477_),
    .Y(_13478_));
 sky130_fd_sc_hd__nor2_1 _34477_ (.A(_13262_),
    .B(_13478_),
    .Y(_13479_));
 sky130_fd_sc_hd__nand2_1 _34478_ (.A(_13474_),
    .B(_13479_),
    .Y(_13480_));
 sky130_fd_sc_hd__a21oi_1 _34479_ (.A1(_02998_),
    .A2(_03003_),
    .B1(_02997_),
    .Y(_13481_));
 sky130_fd_sc_hd__o21ai_0 _34480_ (.A1(_13475_),
    .A2(_13361_),
    .B1(_13481_),
    .Y(_13482_));
 sky130_fd_sc_hd__a21oi_1 _34481_ (.A1(_13265_),
    .A2(_13477_),
    .B1(_13482_),
    .Y(_13483_));
 sky130_fd_sc_hd__nand3_1 _34482_ (.A(_13176_),
    .B(_13479_),
    .C(_13177_),
    .Y(_13484_));
 sky130_fd_sc_hd__nand3_1 _34483_ (.A(_13480_),
    .B(_13483_),
    .C(_13484_),
    .Y(_13485_));
 sky130_fd_sc_hd__nand2_1 _34484_ (.A(_03010_),
    .B(_03016_),
    .Y(_13486_));
 sky130_fd_sc_hd__nor3_1 _34485_ (.A(_02998_),
    .B(_03004_),
    .C(_13486_),
    .Y(_13487_));
 sky130_fd_sc_hd__and3_1 _34486_ (.A(_13487_),
    .B(_13140_),
    .C(_13268_),
    .X(_13488_));
 sky130_fd_sc_hd__nand2_1 _34487_ (.A(_13142_),
    .B(_13133_),
    .Y(_13489_));
 sky130_fd_sc_hd__nand3_1 _34488_ (.A(_13150_),
    .B(_13071_),
    .C(_13154_),
    .Y(_13490_));
 sky130_fd_sc_hd__nor2_1 _34489_ (.A(_13489_),
    .B(_13490_),
    .Y(_13491_));
 sky130_fd_sc_hd__nand3_1 _34490_ (.A(_13488_),
    .B(\inst$top.soc.cpu.multiplier.x_prod[0] ),
    .C(_13491_),
    .Y(_13492_));
 sky130_fd_sc_hd__o21ai_0 _34491_ (.A1(_03076_),
    .A2(_00207_),
    .B1(_00192_),
    .Y(_13493_));
 sky130_fd_sc_hd__nand2_1 _34492_ (.A(_13493_),
    .B(_13150_),
    .Y(_13494_));
 sky130_fd_sc_hd__nand2_1 _34493_ (.A(_13494_),
    .B(_13136_),
    .Y(_13495_));
 sky130_fd_sc_hd__inv_1 _34494_ (.A(_13489_),
    .Y(_13496_));
 sky130_fd_sc_hd__nand2_1 _34495_ (.A(_13495_),
    .B(_13496_),
    .Y(_13497_));
 sky130_fd_sc_hd__nor2_1 _34496_ (.A(_13143_),
    .B(_13138_),
    .Y(_13498_));
 sky130_fd_sc_hd__nor2_1 _34497_ (.A(_13145_),
    .B(_13498_),
    .Y(_13499_));
 sky130_fd_sc_hd__nand2_1 _34498_ (.A(_13497_),
    .B(_13499_),
    .Y(_13500_));
 sky130_fd_sc_hd__nand2_1 _34499_ (.A(_13500_),
    .B(_13488_),
    .Y(_13501_));
 sky130_fd_sc_hd__inv_1 _34500_ (.A(_13268_),
    .Y(_13502_));
 sky130_fd_sc_hd__o21ai_0 _34501_ (.A1(_13502_),
    .A2(_13147_),
    .B1(_13271_),
    .Y(_13503_));
 sky130_fd_sc_hd__o21ai_0 _34502_ (.A1(_00940_),
    .A2(_13325_),
    .B1(_01062_),
    .Y(_13504_));
 sky130_fd_sc_hd__nor2_1 _34503_ (.A(_02998_),
    .B(_03004_),
    .Y(_13505_));
 sky130_fd_sc_hd__nand2_1 _34504_ (.A(_13504_),
    .B(_13505_),
    .Y(_13506_));
 sky130_fd_sc_hd__a21oi_1 _34505_ (.A1(_13446_),
    .A2(_03006_),
    .B1(_03000_),
    .Y(_13507_));
 sky130_fd_sc_hd__nand2_1 _34506_ (.A(_13506_),
    .B(_13507_),
    .Y(_13508_));
 sky130_fd_sc_hd__a21oi_1 _34507_ (.A1(_13503_),
    .A2(_13487_),
    .B1(_13508_),
    .Y(_13509_));
 sky130_fd_sc_hd__nand3_1 _34508_ (.A(_13492_),
    .B(_13501_),
    .C(_13509_),
    .Y(_13510_));
 sky130_fd_sc_hd__nand2_1 _34509_ (.A(_13510_),
    .B(net2006),
    .Y(_13511_));
 sky130_fd_sc_hd__o21ai_0 _34510_ (.A1(net2006),
    .A2(_13485_),
    .B1(_13511_),
    .Y(_13512_));
 sky130_fd_sc_hd__or2_2 _34511_ (.A(_13473_),
    .B(_13512_),
    .X(_13513_));
 sky130_fd_sc_hd__nand2_1 _34512_ (.A(_13512_),
    .B(_13473_),
    .Y(_13514_));
 sky130_fd_sc_hd__nand2_2 _34513_ (.A(_13513_),
    .B(_13514_),
    .Y(_13515_));
 sky130_fd_sc_hd__o21ai_0 _34514_ (.A1(net2844),
    .A2(_13515_),
    .B1(_05640_),
    .Y(_13516_));
 sky130_fd_sc_hd__nand2_1 _34515_ (.A(net1795),
    .B(_03208_),
    .Y(_13517_));
 sky130_fd_sc_hd__nand2_1 _34516_ (.A(net1868),
    .B(_03207_),
    .Y(_13518_));
 sky130_fd_sc_hd__o211ai_1 _34517_ (.A1(_03211_),
    .A2(net1229),
    .B1(_13517_),
    .C1(_13518_),
    .Y(_13519_));
 sky130_fd_sc_hd__nand2_1 _34518_ (.A(_13519_),
    .B(net2862),
    .Y(_13520_));
 sky130_fd_sc_hd__nand2_1 _34519_ (.A(_13520_),
    .B(net2001),
    .Y(_13521_));
 sky130_fd_sc_hd__a21oi_1 _34520_ (.A1(_13516_),
    .A2(net2017),
    .B1(_13521_),
    .Y(_13522_));
 sky130_fd_sc_hd__nor2_2 _34521_ (.A(_13472_),
    .B(_13522_),
    .Y(_13523_));
 sky130_fd_sc_hd__inv_1 _34522_ (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[17] ),
    .Y(_13524_));
 sky130_fd_sc_hd__inv_1 _34523_ (.A(\inst$top.soc.cpu.sink__payload$18[126] ),
    .Y(_13525_));
 sky130_fd_sc_hd__nor2_1 _34524_ (.A(\inst$top.soc.cpu.shifter.m_result$7[17] ),
    .B(net2003),
    .Y(_13526_));
 sky130_fd_sc_hd__o21ai_0 _34525_ (.A1(net2872),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[14] ),
    .B1(net2839),
    .Y(_13527_));
 sky130_fd_sc_hd__o22ai_1 _34526_ (.A1(_13525_),
    .A2(net2839),
    .B1(_13526_),
    .B2(_13527_),
    .Y(_13528_));
 sky130_fd_sc_hd__nand2_1 _34527_ (.A(_13528_),
    .B(net2015),
    .Y(_13529_));
 sky130_fd_sc_hd__a21oi_1 _34528_ (.A1(_10497_),
    .A2(net2918),
    .B1(net2011),
    .Y(_13530_));
 sky130_fd_sc_hd__o21ai_2 _34529_ (.A1(net2918),
    .A2(\inst$top.soc.cpu.divider.quotient[17] ),
    .B1(_13530_),
    .Y(_13531_));
 sky130_fd_sc_hd__a21oi_1 _34530_ (.A1(_13529_),
    .A2(net1791),
    .B1(net2830),
    .Y(_13532_));
 sky130_fd_sc_hd__nand2_1 _34531_ (.A(_12984_),
    .B(_13532_),
    .Y(_13533_));
 sky130_fd_sc_hd__o21ai_0 _34532_ (.A1(_13524_),
    .A2(_12956_),
    .B1(_13533_),
    .Y(_13534_));
 sky130_fd_sc_hd__a21oi_1 _34533_ (.A1(_12959_),
    .A2(_13523_),
    .B1(_13534_),
    .Y(_13535_));
 sky130_fd_sc_hd__nand2_1 _34534_ (.A(net712),
    .B(_13535_),
    .Y(_13536_));
 sky130_fd_sc_hd__nand2_1 _34536_ (.A(_13536_),
    .B(net2173),
    .Y(_13538_));
 sky130_fd_sc_hd__nor2_2 _34537_ (.A(_13468_),
    .B(_13538_),
    .Y(_04192_));
 sky130_fd_sc_hd__nand2_1 _34538_ (.A(_02993_),
    .B(_02998_),
    .Y(_13539_));
 sky130_fd_sc_hd__inv_1 _34539_ (.A(_13539_),
    .Y(_13540_));
 sky130_fd_sc_hd__nand2_1 _34540_ (.A(_13442_),
    .B(_13540_),
    .Y(_13541_));
 sky130_fd_sc_hd__a21oi_1 _34541_ (.A1(_02993_),
    .A2(_02997_),
    .B1(_02992_),
    .Y(_13542_));
 sky130_fd_sc_hd__nand2_1 _34542_ (.A(_13541_),
    .B(_13542_),
    .Y(_13543_));
 sky130_fd_sc_hd__nand2_1 _34543_ (.A(_13543_),
    .B(net2868),
    .Y(_13544_));
 sky130_fd_sc_hd__nand2_1 _34544_ (.A(_13070_),
    .B(_13079_),
    .Y(_13545_));
 sky130_fd_sc_hd__nand2_1 _34545_ (.A(_13303_),
    .B(_13198_),
    .Y(_13546_));
 sky130_fd_sc_hd__nand2_1 _34546_ (.A(_13473_),
    .B(_13446_),
    .Y(_13547_));
 sky130_fd_sc_hd__nor2_1 _34547_ (.A(_13547_),
    .B(_13421_),
    .Y(_13548_));
 sky130_fd_sc_hd__inv_1 _34548_ (.A(_13548_),
    .Y(_13549_));
 sky130_fd_sc_hd__nor2_1 _34549_ (.A(_13546_),
    .B(_13549_),
    .Y(_13550_));
 sky130_fd_sc_hd__nand2_1 _34550_ (.A(_13545_),
    .B(_13550_),
    .Y(_13551_));
 sky130_fd_sc_hd__o21ai_0 _34551_ (.A1(_13419_),
    .A2(_13201_),
    .B1(_13307_),
    .Y(_13552_));
 sky130_fd_sc_hd__nand3_1 _34552_ (.A(_13426_),
    .B(_13473_),
    .C(_13446_),
    .Y(_13553_));
 sky130_fd_sc_hd__a21oi_1 _34553_ (.A1(_13473_),
    .A2(_03000_),
    .B1(_01428_),
    .Y(_13554_));
 sky130_fd_sc_hd__nand2_1 _34554_ (.A(_13553_),
    .B(_13554_),
    .Y(_13555_));
 sky130_fd_sc_hd__a21oi_1 _34555_ (.A1(_13552_),
    .A2(_13548_),
    .B1(_13555_),
    .Y(_13556_));
 sky130_fd_sc_hd__nand3_1 _34556_ (.A(_13550_),
    .B(_13073_),
    .C(_13074_),
    .Y(_13557_));
 sky130_fd_sc_hd__nand4_1 _34557_ (.A(_13551_),
    .B(_13556_),
    .C(net2008),
    .D(_13557_),
    .Y(_13558_));
 sky130_fd_sc_hd__nand2_1 _34558_ (.A(_13544_),
    .B(_13558_),
    .Y(_13559_));
 sky130_fd_sc_hd__inv_1 _34559_ (.A(_02988_),
    .Y(_13560_));
 sky130_fd_sc_hd__nand2_1 _34560_ (.A(_13559_),
    .B(_13560_),
    .Y(_13561_));
 sky130_fd_sc_hd__nand3_1 _34561_ (.A(_13544_),
    .B(_02988_),
    .C(_13558_),
    .Y(_13562_));
 sky130_fd_sc_hd__nand2_1 _34562_ (.A(_13561_),
    .B(_13562_),
    .Y(_13563_));
 sky130_fd_sc_hd__inv_1 _34563_ (.A(_13563_),
    .Y(_13564_));
 sky130_fd_sc_hd__o21ai_0 _34564_ (.A1(net2848),
    .A2(_13564_),
    .B1(_05661_),
    .Y(_13565_));
 sky130_fd_sc_hd__nand2_1 _34565_ (.A(_13565_),
    .B(net2020),
    .Y(_13566_));
 sky130_fd_sc_hd__nand2_1 _34566_ (.A(net1796),
    .B(_03215_),
    .Y(_13567_));
 sky130_fd_sc_hd__nand2_1 _34567_ (.A(net1871),
    .B(_03214_),
    .Y(_13568_));
 sky130_fd_sc_hd__o211ai_1 _34568_ (.A1(_03218_),
    .A2(net1232),
    .B1(_13567_),
    .C1(_13568_),
    .Y(_13569_));
 sky130_fd_sc_hd__a21oi_1 _34569_ (.A1(_13569_),
    .A2(net2863),
    .B1(net2856),
    .Y(_13570_));
 sky130_fd_sc_hd__nor2_1 _34570_ (.A(_05622_),
    .B(_13460_),
    .Y(_13571_));
 sky130_fd_sc_hd__o21ai_0 _34571_ (.A1(_05644_),
    .A2(_13571_),
    .B1(net2855),
    .Y(_13572_));
 sky130_fd_sc_hd__a21oi_1 _34572_ (.A1(_05644_),
    .A2(_13571_),
    .B1(_13572_),
    .Y(_13573_));
 sky130_fd_sc_hd__a21oi_1 _34573_ (.A1(_13566_),
    .A2(_13570_),
    .B1(_13573_),
    .Y(_13574_));
 sky130_fd_sc_hd__inv_1 _34574_ (.A(_13574_),
    .Y(_13575_));
 sky130_fd_sc_hd__inv_1 _34575_ (.A(\inst$top.soc.cpu.sink__payload$18[127] ),
    .Y(_13576_));
 sky130_fd_sc_hd__nor2_1 _34576_ (.A(net2834),
    .B(_13576_),
    .Y(_13577_));
 sky130_fd_sc_hd__inv_1 _34577_ (.A(\inst$top.soc.cpu.shifter.m_result$7[18] ),
    .Y(_13578_));
 sky130_fd_sc_hd__o21ai_0 _34578_ (.A1(net2871),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[13] ),
    .B1(net2836),
    .Y(_13579_));
 sky130_fd_sc_hd__a21oi_1 _34579_ (.A1(net2871),
    .A2(_13578_),
    .B1(_13579_),
    .Y(_13580_));
 sky130_fd_sc_hd__o21ai_0 _34580_ (.A1(_13577_),
    .A2(_13580_),
    .B1(net2013),
    .Y(_13581_));
 sky130_fd_sc_hd__a21oi_1 _34581_ (.A1(_10516_),
    .A2(net2918),
    .B1(net2011),
    .Y(_13582_));
 sky130_fd_sc_hd__o21ai_1 _34582_ (.A1(net2918),
    .A2(\inst$top.soc.cpu.divider.quotient[18] ),
    .B1(_13582_),
    .Y(_13583_));
 sky130_fd_sc_hd__nand2_1 _34583_ (.A(_13581_),
    .B(net1790),
    .Y(_13584_));
 sky130_fd_sc_hd__nand2_1 _34584_ (.A(_13584_),
    .B(_12997_),
    .Y(_13585_));
 sky130_fd_sc_hd__nor2_1 _34585_ (.A(_13585_),
    .B(net783),
    .Y(_13586_));
 sky130_fd_sc_hd__a21oi_1 _34586_ (.A1(net737),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[18] ),
    .B1(_13586_),
    .Y(_13587_));
 sky130_fd_sc_hd__o21ai_0 _34587_ (.A1(net736),
    .A2(_13575_),
    .B1(_13587_),
    .Y(_13588_));
 sky130_fd_sc_hd__nand2_1 _34588_ (.A(net709),
    .B(_13588_),
    .Y(_13589_));
 sky130_fd_sc_hd__nand2_1 _34589_ (.A(net657),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[18] ),
    .Y(_13590_));
 sky130_fd_sc_hd__a21oi_4 _34590_ (.A1(_13589_),
    .A2(_13590_),
    .B1(net2993),
    .Y(_04193_));
 sky130_fd_sc_hd__inv_1 _34593_ (.A(\inst$top.soc.cpu.sink__payload$18[128] ),
    .Y(_13593_));
 sky130_fd_sc_hd__nor2_1 _34594_ (.A(net2834),
    .B(_13593_),
    .Y(_13594_));
 sky130_fd_sc_hd__inv_1 _34596_ (.A(\inst$top.soc.cpu.shifter.m_result$7[19] ),
    .Y(_13596_));
 sky130_fd_sc_hd__o21ai_0 _34597_ (.A1(net2872),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[12] ),
    .B1(net2837),
    .Y(_13597_));
 sky130_fd_sc_hd__a21oi_1 _34598_ (.A1(net2873),
    .A2(_13596_),
    .B1(_13597_),
    .Y(_13598_));
 sky130_fd_sc_hd__o21ai_0 _34600_ (.A1(_13594_),
    .A2(_13598_),
    .B1(net2016),
    .Y(_13600_));
 sky130_fd_sc_hd__a21oi_1 _34602_ (.A1(_10530_),
    .A2(net2919),
    .B1(net2010),
    .Y(_13602_));
 sky130_fd_sc_hd__o21ai_1 _34603_ (.A1(net2919),
    .A2(\inst$top.soc.cpu.divider.quotient[19] ),
    .B1(_13602_),
    .Y(_13603_));
 sky130_fd_sc_hd__a21oi_1 _34605_ (.A1(_13600_),
    .A2(net1789),
    .B1(net2829),
    .Y(_13605_));
 sky130_fd_sc_hd__inv_1 _34606_ (.A(_13605_),
    .Y(_13606_));
 sky130_fd_sc_hd__nand2_1 _34608_ (.A(net738),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[19] ),
    .Y(_13608_));
 sky130_fd_sc_hd__nand2_1 _34609_ (.A(\inst$top.soc.cpu.sink__payload$12[18] ),
    .B(\inst$top.soc.cpu.sink__payload$12[17] ),
    .Y(_13609_));
 sky130_fd_sc_hd__o21ai_0 _34610_ (.A1(_13609_),
    .A2(_13469_),
    .B1(\inst$top.soc.cpu.sink__payload$12[19] ),
    .Y(_13610_));
 sky130_fd_sc_hd__nor4_1 _34611_ (.A(_05598_),
    .B(_20807_),
    .C(_13609_),
    .D(_13384_),
    .Y(_13611_));
 sky130_fd_sc_hd__a21oi_1 _34612_ (.A1(_13611_),
    .A2(_05666_),
    .B1(net2001),
    .Y(_13612_));
 sky130_fd_sc_hd__nor2_1 _34613_ (.A(_02988_),
    .B(_02993_),
    .Y(_13613_));
 sky130_fd_sc_hd__nand2_1 _34614_ (.A(_13505_),
    .B(_13613_),
    .Y(_13614_));
 sky130_fd_sc_hd__nor2_1 _34615_ (.A(_13486_),
    .B(_13271_),
    .Y(_13615_));
 sky130_fd_sc_hd__nor2_1 _34616_ (.A(_13504_),
    .B(_13615_),
    .Y(_13616_));
 sky130_fd_sc_hd__o21bai_1 _34617_ (.A1(_02988_),
    .A2(_01427_),
    .B1_N(_01539_),
    .Y(_13617_));
 sky130_fd_sc_hd__inv_1 _34618_ (.A(_13613_),
    .Y(_13618_));
 sky130_fd_sc_hd__nor2_1 _34619_ (.A(_13618_),
    .B(_13507_),
    .Y(_13619_));
 sky130_fd_sc_hd__nor2_1 _34620_ (.A(_13617_),
    .B(_13619_),
    .Y(_13620_));
 sky130_fd_sc_hd__o21ai_0 _34621_ (.A1(_13614_),
    .A2(_13616_),
    .B1(_13620_),
    .Y(_13621_));
 sky130_fd_sc_hd__inv_1 _34622_ (.A(_13149_),
    .Y(_13622_));
 sky130_fd_sc_hd__nor3_1 _34623_ (.A(_13502_),
    .B(_13486_),
    .C(_13614_),
    .Y(_13623_));
 sky130_fd_sc_hd__nand2_1 _34624_ (.A(_13622_),
    .B(_13623_),
    .Y(_13624_));
 sky130_fd_sc_hd__nand3_1 _34625_ (.A(_13153_),
    .B(_13156_),
    .C(_13623_),
    .Y(_13625_));
 sky130_fd_sc_hd__nand3b_1 _34626_ (.A_N(_13621_),
    .B(_13624_),
    .C(_13625_),
    .Y(_13626_));
 sky130_fd_sc_hd__nand2_1 _34627_ (.A(_13626_),
    .B(net2006),
    .Y(_13627_));
 sky130_fd_sc_hd__nor2_1 _34628_ (.A(_13167_),
    .B(_13163_),
    .Y(_13628_));
 sky130_fd_sc_hd__nor2_1 _34629_ (.A(_13180_),
    .B(_13165_),
    .Y(_13629_));
 sky130_fd_sc_hd__o21ai_0 _34630_ (.A1(_13171_),
    .A2(_13628_),
    .B1(_13629_),
    .Y(_13630_));
 sky130_fd_sc_hd__a21boi_0 _34631_ (.A1(_13172_),
    .A2(_13181_),
    .B1_N(_13183_),
    .Y(_13631_));
 sky130_fd_sc_hd__nand2_1 _34632_ (.A(_13630_),
    .B(_13631_),
    .Y(_13632_));
 sky130_fd_sc_hd__nand2_1 _34633_ (.A(_02988_),
    .B(_02993_),
    .Y(_13633_));
 sky130_fd_sc_hd__nor2_1 _34634_ (.A(_13475_),
    .B(_13633_),
    .Y(_13634_));
 sky130_fd_sc_hd__inv_1 _34635_ (.A(_13634_),
    .Y(_13635_));
 sky130_fd_sc_hd__nor2_1 _34636_ (.A(_13260_),
    .B(_13476_),
    .Y(_13636_));
 sky130_fd_sc_hd__inv_1 _34637_ (.A(_13636_),
    .Y(_13637_));
 sky130_fd_sc_hd__nor2_1 _34638_ (.A(_13635_),
    .B(_13637_),
    .Y(_13638_));
 sky130_fd_sc_hd__o21a_1 _34639_ (.A1(_13476_),
    .A2(_13264_),
    .B1(_13361_),
    .X(_13639_));
 sky130_fd_sc_hd__a21oi_1 _34640_ (.A1(_02988_),
    .A2(_02992_),
    .B1(_02987_),
    .Y(_13640_));
 sky130_fd_sc_hd__o21ai_0 _34641_ (.A1(_13633_),
    .A2(_13481_),
    .B1(_13640_),
    .Y(_13641_));
 sky130_fd_sc_hd__o21bai_1 _34642_ (.A1(_13635_),
    .A2(_13639_),
    .B1_N(_13641_),
    .Y(_13642_));
 sky130_fd_sc_hd__a21oi_1 _34643_ (.A1(_13632_),
    .A2(_13638_),
    .B1(_13642_),
    .Y(_13643_));
 sky130_fd_sc_hd__inv_1 _34644_ (.A(_13629_),
    .Y(_13644_));
 sky130_fd_sc_hd__nor3_1 _34645_ (.A(_13167_),
    .B(_13160_),
    .C(_13644_),
    .Y(_13645_));
 sky130_fd_sc_hd__nand3_1 _34646_ (.A(_13257_),
    .B(_13645_),
    .C(_13638_),
    .Y(_13646_));
 sky130_fd_sc_hd__nand3_1 _34647_ (.A(_13643_),
    .B(net2867),
    .C(_13646_),
    .Y(_13647_));
 sky130_fd_sc_hd__nand2_1 _34648_ (.A(_13627_),
    .B(_13647_),
    .Y(_13648_));
 sky130_fd_sc_hd__inv_1 _34649_ (.A(_02982_),
    .Y(_13649_));
 sky130_fd_sc_hd__nand2_1 _34650_ (.A(_13648_),
    .B(_13649_),
    .Y(_13650_));
 sky130_fd_sc_hd__nand3_1 _34651_ (.A(_13627_),
    .B(_02982_),
    .C(_13647_),
    .Y(_13651_));
 sky130_fd_sc_hd__nand2_1 _34652_ (.A(_13650_),
    .B(_13651_),
    .Y(_13652_));
 sky130_fd_sc_hd__inv_1 _34653_ (.A(_13652_),
    .Y(_13653_));
 sky130_fd_sc_hd__o21ai_0 _34654_ (.A1(net2845),
    .A2(_13653_),
    .B1(_05684_),
    .Y(_13654_));
 sky130_fd_sc_hd__nand2_1 _34655_ (.A(net1795),
    .B(_03222_),
    .Y(_13655_));
 sky130_fd_sc_hd__nand2_1 _34656_ (.A(net1868),
    .B(_03221_),
    .Y(_13656_));
 sky130_fd_sc_hd__o211ai_1 _34657_ (.A1(_03225_),
    .A2(net1229),
    .B1(_13655_),
    .C1(_13656_),
    .Y(_13657_));
 sky130_fd_sc_hd__a21oi_1 _34658_ (.A1(_13657_),
    .A2(net2862),
    .B1(net2854),
    .Y(_13658_));
 sky130_fd_sc_hd__a21boi_0 _34659_ (.A1(_13654_),
    .A2(net2017),
    .B1_N(_13658_),
    .Y(_13659_));
 sky130_fd_sc_hd__a21oi_2 _34660_ (.A1(_13610_),
    .A2(_13612_),
    .B1(_13659_),
    .Y(_13660_));
 sky130_fd_sc_hd__nand2_1 _34661_ (.A(_13660_),
    .B(net786),
    .Y(_13661_));
 sky130_fd_sc_hd__o211ai_1 _34662_ (.A1(net785),
    .A2(_13606_),
    .B1(_13608_),
    .C1(_13661_),
    .Y(_13662_));
 sky130_fd_sc_hd__nor2_1 _34663_ (.A(net657),
    .B(_13662_),
    .Y(_13663_));
 sky130_fd_sc_hd__nand2_1 _34665_ (.A(net657),
    .B(_05667_),
    .Y(_13665_));
 sky130_fd_sc_hd__nand2_1 _34666_ (.A(_13665_),
    .B(net2156),
    .Y(_13666_));
 sky130_fd_sc_hd__nor2_4 _34667_ (.A(_13663_),
    .B(_13666_),
    .Y(_04194_));
 sky130_fd_sc_hd__nor2_1 _34668_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[1] ),
    .B(net701),
    .Y(_13667_));
 sky130_fd_sc_hd__inv_1 _34669_ (.A(\inst$top.soc.cpu.sink__payload$18[110] ),
    .Y(_13668_));
 sky130_fd_sc_hd__nor2_1 _34670_ (.A(\inst$top.soc.cpu.shifter.m_result$7[1] ),
    .B(net2002),
    .Y(_13669_));
 sky130_fd_sc_hd__o21ai_0 _34671_ (.A1(net2869),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[30] ),
    .B1(net2833),
    .Y(_13670_));
 sky130_fd_sc_hd__o22ai_1 _34672_ (.A1(_13668_),
    .A2(net2833),
    .B1(_13669_),
    .B2(_13670_),
    .Y(_13671_));
 sky130_fd_sc_hd__nand2_1 _34673_ (.A(_13671_),
    .B(net2014),
    .Y(_13672_));
 sky130_fd_sc_hd__a21oi_1 _34674_ (.A1(_02854_),
    .A2(net2923),
    .B1(net2011),
    .Y(_13673_));
 sky130_fd_sc_hd__o21ai_1 _34675_ (.A1(net2922),
    .A2(\inst$top.soc.cpu.divider.quotient[1] ),
    .B1(_13673_),
    .Y(_13674_));
 sky130_fd_sc_hd__a21oi_1 _34676_ (.A1(_13672_),
    .A2(net1788),
    .B1(net2829),
    .Y(_13675_));
 sky130_fd_sc_hd__inv_1 _34677_ (.A(_13675_),
    .Y(_13676_));
 sky130_fd_sc_hd__nor2_1 _34679_ (.A(_03097_),
    .B(net1231),
    .Y(_13678_));
 sky130_fd_sc_hd__a221oi_1 _34680_ (.A1(net1798),
    .A2(_03094_),
    .B1(net1871),
    .B2(_03093_),
    .C1(_13678_),
    .Y(_13679_));
 sky130_fd_sc_hd__or2_2 _34681_ (.A(_00171_),
    .B(net2005),
    .X(_13680_));
 sky130_fd_sc_hd__o21ai_1 _34682_ (.A1(net2865),
    .A2(_00166_),
    .B1(_13680_),
    .Y(_13681_));
 sky130_fd_sc_hd__inv_1 _34683_ (.A(_13681_),
    .Y(_13682_));
 sky130_fd_sc_hd__nand2_1 _34684_ (.A(_13682_),
    .B(net2214),
    .Y(_13683_));
 sky130_fd_sc_hd__a21oi_1 _34685_ (.A1(_20441_),
    .A2(_13683_),
    .B1(net2863),
    .Y(_13684_));
 sky130_fd_sc_hd__a211oi_1 _34686_ (.A1(net2863),
    .A2(_13679_),
    .B1(net2855),
    .C1(_13684_),
    .Y(_13685_));
 sky130_fd_sc_hd__inv_1 _34687_ (.A(_13685_),
    .Y(_13686_));
 sky130_fd_sc_hd__o22ai_1 _34688_ (.A1(_13676_),
    .A2(net783),
    .B1(_13686_),
    .B2(net736),
    .Y(_13687_));
 sky130_fd_sc_hd__a21oi_1 _34689_ (.A1(net737),
    .A2(net1017),
    .B1(_13687_),
    .Y(_13688_));
 sky130_fd_sc_hd__nand2_1 _34690_ (.A(net696),
    .B(_13688_),
    .Y(_13689_));
 sky130_fd_sc_hd__nand2_1 _34691_ (.A(_13689_),
    .B(net2151),
    .Y(_13690_));
 sky130_fd_sc_hd__nor2_2 _34692_ (.A(_13667_),
    .B(_13690_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand2_1 _34693_ (.A(\inst$top.soc.cpu.sink__payload$12[19] ),
    .B(\inst$top.soc.cpu.sink__payload$12[18] ),
    .Y(_13691_));
 sky130_fd_sc_hd__inv_1 _34694_ (.A(_13691_),
    .Y(_13692_));
 sky130_fd_sc_hd__nand2_1 _34695_ (.A(_13571_),
    .B(_13692_),
    .Y(_13693_));
 sky130_fd_sc_hd__nand2_1 _34696_ (.A(_13693_),
    .B(\inst$top.soc.cpu.sink__payload$12[20] ),
    .Y(_13694_));
 sky130_fd_sc_hd__nand2_1 _34697_ (.A(_13694_),
    .B(net2854),
    .Y(_13695_));
 sky130_fd_sc_hd__nor2_1 _34698_ (.A(\inst$top.soc.cpu.sink__payload$12[20] ),
    .B(_13693_),
    .Y(_13696_));
 sky130_fd_sc_hd__nand2_1 _34699_ (.A(net1795),
    .B(_03229_),
    .Y(_13697_));
 sky130_fd_sc_hd__nand2_1 _34700_ (.A(net1868),
    .B(_03228_),
    .Y(_13698_));
 sky130_fd_sc_hd__o211ai_1 _34701_ (.A1(_03232_),
    .A2(net1229),
    .B1(_13697_),
    .C1(_13698_),
    .Y(_13699_));
 sky130_fd_sc_hd__a21oi_1 _34702_ (.A1(_13699_),
    .A2(net2862),
    .B1(net2854),
    .Y(_13700_));
 sky130_fd_sc_hd__nor2_1 _34703_ (.A(_02982_),
    .B(_13560_),
    .Y(_13701_));
 sky130_fd_sc_hd__inv_1 _34704_ (.A(_13701_),
    .Y(_13702_));
 sky130_fd_sc_hd__nor2_1 _34705_ (.A(_13539_),
    .B(_13702_),
    .Y(_13703_));
 sky130_fd_sc_hd__nand2_1 _34706_ (.A(_13442_),
    .B(_13703_),
    .Y(_13704_));
 sky130_fd_sc_hd__a21oi_1 _34707_ (.A1(_13649_),
    .A2(_02987_),
    .B1(_02984_),
    .Y(_13705_));
 sky130_fd_sc_hd__o21ai_0 _34708_ (.A1(_13702_),
    .A2(_13542_),
    .B1(_13705_),
    .Y(_13706_));
 sky130_fd_sc_hd__inv_1 _34709_ (.A(_13706_),
    .Y(_13707_));
 sky130_fd_sc_hd__nand3_1 _34710_ (.A(_13704_),
    .B(net2868),
    .C(_13707_),
    .Y(_13708_));
 sky130_fd_sc_hd__nor2_1 _34711_ (.A(_02988_),
    .B(_13649_),
    .Y(_13709_));
 sky130_fd_sc_hd__inv_1 _34712_ (.A(_13709_),
    .Y(_13710_));
 sky130_fd_sc_hd__nor2_1 _34713_ (.A(_13547_),
    .B(_13710_),
    .Y(_13711_));
 sky130_fd_sc_hd__inv_1 _34714_ (.A(_13711_),
    .Y(_13712_));
 sky130_fd_sc_hd__a21oi_1 _34715_ (.A1(_01539_),
    .A2(_02982_),
    .B1(_02981_),
    .Y(_13713_));
 sky130_fd_sc_hd__o21a_1 _34716_ (.A1(_13710_),
    .A2(_13554_),
    .B1(_13713_),
    .X(_13714_));
 sky130_fd_sc_hd__o21ai_0 _34717_ (.A1(_13712_),
    .A2(_13427_),
    .B1(_13714_),
    .Y(_13715_));
 sky130_fd_sc_hd__a21oi_1 _34718_ (.A1(_13415_),
    .A2(_13067_),
    .B1(_13077_),
    .Y(_13716_));
 sky130_fd_sc_hd__o21ai_0 _34719_ (.A1(_13418_),
    .A2(_13716_),
    .B1(_13425_),
    .Y(_13717_));
 sky130_fd_sc_hd__nor2_1 _34720_ (.A(_13712_),
    .B(_13423_),
    .Y(_13718_));
 sky130_fd_sc_hd__nand2_1 _34721_ (.A(_13717_),
    .B(_13718_),
    .Y(_13719_));
 sky130_fd_sc_hd__nor3_1 _34722_ (.A(_13412_),
    .B(_13060_),
    .C(_13418_),
    .Y(_13720_));
 sky130_fd_sc_hd__nand3_1 _34723_ (.A(_13718_),
    .B(_13414_),
    .C(_13720_),
    .Y(_13721_));
 sky130_fd_sc_hd__nand3b_1 _34724_ (.A_N(_13715_),
    .B(_13719_),
    .C(_13721_),
    .Y(_13722_));
 sky130_fd_sc_hd__nand2_1 _34725_ (.A(_13722_),
    .B(net2008),
    .Y(_13723_));
 sky130_fd_sc_hd__nand2_1 _34726_ (.A(_13708_),
    .B(_13723_),
    .Y(_13724_));
 sky130_fd_sc_hd__inv_1 _34727_ (.A(_02976_),
    .Y(_13725_));
 sky130_fd_sc_hd__nand2_1 _34728_ (.A(_13724_),
    .B(_13725_),
    .Y(_13726_));
 sky130_fd_sc_hd__nand3_1 _34729_ (.A(_13708_),
    .B(_02976_),
    .C(_13723_),
    .Y(_13727_));
 sky130_fd_sc_hd__nand2_1 _34730_ (.A(_13726_),
    .B(_13727_),
    .Y(_13728_));
 sky130_fd_sc_hd__inv_1 _34731_ (.A(_13728_),
    .Y(_13729_));
 sky130_fd_sc_hd__o21ai_0 _34732_ (.A1(net2843),
    .A2(_13729_),
    .B1(_05706_),
    .Y(_13730_));
 sky130_fd_sc_hd__nand2_1 _34733_ (.A(_13730_),
    .B(net2020),
    .Y(_13731_));
 sky130_fd_sc_hd__a2bb2oi_4 _34734_ (.A1_N(_13695_),
    .A2_N(_13696_),
    .B1(_13700_),
    .B2(_13731_),
    .Y(_13732_));
 sky130_fd_sc_hd__nand2_1 _34735_ (.A(_13732_),
    .B(net786),
    .Y(_13733_));
 sky130_fd_sc_hd__nand2_1 _34736_ (.A(_12957_),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[20] ),
    .Y(_13734_));
 sky130_fd_sc_hd__inv_1 _34737_ (.A(\inst$top.soc.cpu.sink__payload$18[129] ),
    .Y(_13735_));
 sky130_fd_sc_hd__nor2_1 _34739_ (.A(\inst$top.soc.cpu.shifter.m_result$7[20] ),
    .B(net2004),
    .Y(_13737_));
 sky130_fd_sc_hd__o21ai_0 _34740_ (.A1(net2870),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[11] ),
    .B1(net2841),
    .Y(_13738_));
 sky130_fd_sc_hd__o22ai_1 _34741_ (.A1(_13735_),
    .A2(net2841),
    .B1(_13737_),
    .B2(_13738_),
    .Y(_13739_));
 sky130_fd_sc_hd__nand2_1 _34742_ (.A(_13739_),
    .B(net2014),
    .Y(_13740_));
 sky130_fd_sc_hd__a21oi_1 _34743_ (.A1(_10562_),
    .A2(net2919),
    .B1(net2010),
    .Y(_13741_));
 sky130_fd_sc_hd__o21ai_1 _34744_ (.A1(net2919),
    .A2(\inst$top.soc.cpu.divider.quotient[20] ),
    .B1(_13741_),
    .Y(_13742_));
 sky130_fd_sc_hd__a21oi_1 _34745_ (.A1(_13740_),
    .A2(net1787),
    .B1(net2830),
    .Y(_13743_));
 sky130_fd_sc_hd__nand2_1 _34746_ (.A(_12984_),
    .B(_13743_),
    .Y(_13744_));
 sky130_fd_sc_hd__nand3_1 _34747_ (.A(_13733_),
    .B(_13734_),
    .C(_13744_),
    .Y(_13745_));
 sky130_fd_sc_hd__nand2_1 _34748_ (.A(net710),
    .B(_13745_),
    .Y(_13746_));
 sky130_fd_sc_hd__nand2_1 _34749_ (.A(net658),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[20] ),
    .Y(_13747_));
 sky130_fd_sc_hd__a21oi_4 _34750_ (.A1(_13746_),
    .A2(_13747_),
    .B1(net3010),
    .Y(_04196_));
 sky130_fd_sc_hd__inv_1 _34751_ (.A(\inst$top.soc.cpu.sink__payload$18[130] ),
    .Y(_13748_));
 sky130_fd_sc_hd__nor2_1 _34752_ (.A(net2841),
    .B(_13748_),
    .Y(_13749_));
 sky130_fd_sc_hd__o21ai_0 _34753_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[21] ),
    .A2(net2002),
    .B1(net2835),
    .Y(_13750_));
 sky130_fd_sc_hd__a21oi_1 _34754_ (.A1(net2004),
    .A2(_13018_),
    .B1(_13750_),
    .Y(_13751_));
 sky130_fd_sc_hd__o21ai_0 _34755_ (.A1(_13749_),
    .A2(_13751_),
    .B1(net2014),
    .Y(_13752_));
 sky130_fd_sc_hd__a21oi_1 _34756_ (.A1(_10569_),
    .A2(net2919),
    .B1(net2010),
    .Y(_13753_));
 sky130_fd_sc_hd__o21ai_1 _34757_ (.A1(net2919),
    .A2(\inst$top.soc.cpu.divider.quotient[21] ),
    .B1(_13753_),
    .Y(_13754_));
 sky130_fd_sc_hd__a21oi_1 _34758_ (.A1(_13752_),
    .A2(net1786),
    .B1(net2830),
    .Y(_13755_));
 sky130_fd_sc_hd__inv_1 _34759_ (.A(_13755_),
    .Y(_13756_));
 sky130_fd_sc_hd__nand2_1 _34760_ (.A(net739),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[21] ),
    .Y(_13757_));
 sky130_fd_sc_hd__nand2_1 _34761_ (.A(_02976_),
    .B(_02982_),
    .Y(_13758_));
 sky130_fd_sc_hd__nor2_1 _34762_ (.A(_13758_),
    .B(_13618_),
    .Y(_13759_));
 sky130_fd_sc_hd__nand2_1 _34763_ (.A(_13510_),
    .B(_13759_),
    .Y(_13760_));
 sky130_fd_sc_hd__o21ai_0 _34764_ (.A1(_01651_),
    .A2(_13725_),
    .B1(_01753_),
    .Y(_13761_));
 sky130_fd_sc_hd__a31oi_1 _34765_ (.A1(_13617_),
    .A2(_02976_),
    .A3(_02982_),
    .B1(_13761_),
    .Y(_13762_));
 sky130_fd_sc_hd__nand2_1 _34766_ (.A(_13760_),
    .B(_13762_),
    .Y(_13763_));
 sky130_fd_sc_hd__nand2_1 _34767_ (.A(_13763_),
    .B(net2006),
    .Y(_13764_));
 sky130_fd_sc_hd__nor2_1 _34768_ (.A(_02976_),
    .B(_02982_),
    .Y(_13765_));
 sky130_fd_sc_hd__inv_1 _34769_ (.A(_13765_),
    .Y(_13766_));
 sky130_fd_sc_hd__nor3_1 _34770_ (.A(_13633_),
    .B(_13766_),
    .C(_13478_),
    .Y(_13767_));
 sky130_fd_sc_hd__nand3_1 _34771_ (.A(_13259_),
    .B(_13263_),
    .C(_13767_),
    .Y(_13768_));
 sky130_fd_sc_hd__nand2_1 _34772_ (.A(_13266_),
    .B(_13767_),
    .Y(_13769_));
 sky130_fd_sc_hd__nor2_1 _34773_ (.A(_13633_),
    .B(_13766_),
    .Y(_13770_));
 sky130_fd_sc_hd__a21oi_2 _34774_ (.A1(_13725_),
    .A2(_02984_),
    .B1(_02978_),
    .Y(_13771_));
 sky130_fd_sc_hd__o21ai_0 _34775_ (.A1(_13766_),
    .A2(_13640_),
    .B1(_13771_),
    .Y(_13772_));
 sky130_fd_sc_hd__a21o_1 _34776_ (.A1(_13482_),
    .A2(_13770_),
    .B1(_13772_),
    .X(_13773_));
 sky130_fd_sc_hd__inv_1 _34777_ (.A(_13773_),
    .Y(_13774_));
 sky130_fd_sc_hd__nand4_1 _34778_ (.A(_13768_),
    .B(_13769_),
    .C(_13774_),
    .D(net2867),
    .Y(_13775_));
 sky130_fd_sc_hd__nand2_1 _34779_ (.A(_13764_),
    .B(_13775_),
    .Y(_13776_));
 sky130_fd_sc_hd__inv_1 _34780_ (.A(_02972_),
    .Y(_13777_));
 sky130_fd_sc_hd__nand2_1 _34781_ (.A(_13776_),
    .B(_13777_),
    .Y(_13778_));
 sky130_fd_sc_hd__nand3_1 _34782_ (.A(_13764_),
    .B(_02972_),
    .C(_13775_),
    .Y(_13779_));
 sky130_fd_sc_hd__nand2_2 _34783_ (.A(_13778_),
    .B(_13779_),
    .Y(_13780_));
 sky130_fd_sc_hd__o21ai_0 _34784_ (.A1(net2848),
    .A2(_13780_),
    .B1(_05725_),
    .Y(_13781_));
 sky130_fd_sc_hd__nand2_1 _34785_ (.A(_13781_),
    .B(net2018),
    .Y(_13782_));
 sky130_fd_sc_hd__nand2_1 _34786_ (.A(net1797),
    .B(_03236_),
    .Y(_13783_));
 sky130_fd_sc_hd__nand2_1 _34787_ (.A(net1870),
    .B(_03235_),
    .Y(_13784_));
 sky130_fd_sc_hd__o211ai_1 _34788_ (.A1(_03239_),
    .A2(net1231),
    .B1(_13783_),
    .C1(_13784_),
    .Y(_13785_));
 sky130_fd_sc_hd__a21oi_1 _34789_ (.A1(_13785_),
    .A2(net2863),
    .B1(net2855),
    .Y(_13786_));
 sky130_fd_sc_hd__nor4_1 _34790_ (.A(_05598_),
    .B(_20807_),
    .C(_20789_),
    .D(_20771_),
    .Y(_13787_));
 sky130_fd_sc_hd__nand2_1 _34791_ (.A(\inst$top.soc.cpu.sink__payload$12[20] ),
    .B(\inst$top.soc.cpu.sink__payload$12[19] ),
    .Y(_13788_));
 sky130_fd_sc_hd__nor2_1 _34792_ (.A(_13609_),
    .B(_13788_),
    .Y(_13789_));
 sky130_fd_sc_hd__nand3_1 _34793_ (.A(_13291_),
    .B(_13787_),
    .C(_13789_),
    .Y(_13790_));
 sky130_fd_sc_hd__o21ai_0 _34794_ (.A1(\inst$top.soc.cpu.sink__payload$12[21] ),
    .A2(_13790_),
    .B1(net2855),
    .Y(_13791_));
 sky130_fd_sc_hd__a21oi_1 _34795_ (.A1(\inst$top.soc.cpu.sink__payload$12[21] ),
    .A2(_13790_),
    .B1(_13791_),
    .Y(_13792_));
 sky130_fd_sc_hd__a21oi_2 _34796_ (.A1(_13782_),
    .A2(_13786_),
    .B1(_13792_),
    .Y(_13793_));
 sky130_fd_sc_hd__nand2_1 _34797_ (.A(_13793_),
    .B(net786),
    .Y(_13794_));
 sky130_fd_sc_hd__o211ai_1 _34798_ (.A1(net785),
    .A2(_13756_),
    .B1(_13757_),
    .C1(_13794_),
    .Y(_13795_));
 sky130_fd_sc_hd__nand2_1 _34799_ (.A(net713),
    .B(_13795_),
    .Y(_13796_));
 sky130_fd_sc_hd__nand2_1 _34800_ (.A(net659),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[21] ),
    .Y(_13797_));
 sky130_fd_sc_hd__a21oi_4 _34801_ (.A1(_13796_),
    .A2(_13797_),
    .B1(net3003),
    .Y(_04197_));
 sky130_fd_sc_hd__nand2_1 _34803_ (.A(net659),
    .B(_05729_),
    .Y(_13799_));
 sky130_fd_sc_hd__nand2_1 _34805_ (.A(_13799_),
    .B(net2173),
    .Y(_13801_));
 sky130_fd_sc_hd__inv_1 _34806_ (.A(\inst$top.soc.cpu.sink__payload$18[131] ),
    .Y(_13802_));
 sky130_fd_sc_hd__nor2_1 _34807_ (.A(net2838),
    .B(_13802_),
    .Y(_13803_));
 sky130_fd_sc_hd__inv_1 _34808_ (.A(\inst$top.soc.cpu.shifter.m_result$7[22] ),
    .Y(_13804_));
 sky130_fd_sc_hd__o21ai_0 _34809_ (.A1(net2872),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[9] ),
    .B1(net2838),
    .Y(_13805_));
 sky130_fd_sc_hd__a21oi_1 _34810_ (.A1(net2873),
    .A2(_13804_),
    .B1(_13805_),
    .Y(_13806_));
 sky130_fd_sc_hd__o21ai_0 _34811_ (.A1(_13803_),
    .A2(_13806_),
    .B1(net2015),
    .Y(_13807_));
 sky130_fd_sc_hd__a21oi_1 _34812_ (.A1(_10601_),
    .A2(net2921),
    .B1(net2012),
    .Y(_13808_));
 sky130_fd_sc_hd__o21ai_4 _34813_ (.A1(net2921),
    .A2(\inst$top.soc.cpu.divider.quotient[22] ),
    .B1(_13808_),
    .Y(_13809_));
 sky130_fd_sc_hd__a21oi_1 _34814_ (.A1(_13807_),
    .A2(_13809_),
    .B1(net2831),
    .Y(_13810_));
 sky130_fd_sc_hd__inv_1 _34815_ (.A(_13810_),
    .Y(_13811_));
 sky130_fd_sc_hd__nand2_1 _34816_ (.A(net739),
    .B(net948),
    .Y(_13812_));
 sky130_fd_sc_hd__inv_1 _34817_ (.A(_02966_),
    .Y(_13813_));
 sky130_fd_sc_hd__nor2_1 _34818_ (.A(_13539_),
    .B(_13433_),
    .Y(_13814_));
 sky130_fd_sc_hd__inv_1 _34819_ (.A(_13814_),
    .Y(_13815_));
 sky130_fd_sc_hd__nor2_1 _34820_ (.A(_02976_),
    .B(_13777_),
    .Y(_13816_));
 sky130_fd_sc_hd__inv_1 _34821_ (.A(_13816_),
    .Y(_13817_));
 sky130_fd_sc_hd__nor2_1 _34822_ (.A(_13702_),
    .B(_13817_),
    .Y(_13818_));
 sky130_fd_sc_hd__inv_1 _34823_ (.A(_13818_),
    .Y(_13819_));
 sky130_fd_sc_hd__nor2_1 _34824_ (.A(_13815_),
    .B(_13819_),
    .Y(_13820_));
 sky130_fd_sc_hd__inv_1 _34825_ (.A(_13820_),
    .Y(_13821_));
 sky130_fd_sc_hd__o21ai_0 _34826_ (.A1(_13539_),
    .A2(_13439_),
    .B1(_13542_),
    .Y(_13822_));
 sky130_fd_sc_hd__a21oi_1 _34827_ (.A1(_02972_),
    .A2(_02978_),
    .B1(_02971_),
    .Y(_13823_));
 sky130_fd_sc_hd__o21ai_0 _34828_ (.A1(_13817_),
    .A2(_13705_),
    .B1(_13823_),
    .Y(_13824_));
 sky130_fd_sc_hd__a21oi_1 _34829_ (.A1(_13822_),
    .A2(_13818_),
    .B1(_13824_),
    .Y(_13825_));
 sky130_fd_sc_hd__nand3_1 _34830_ (.A(_13317_),
    .B(_13319_),
    .C(_13820_),
    .Y(_13826_));
 sky130_fd_sc_hd__o211ai_1 _34831_ (.A1(_13821_),
    .A2(_13316_),
    .B1(_13825_),
    .C1(_13826_),
    .Y(_13827_));
 sky130_fd_sc_hd__nor2_1 _34832_ (.A(_13546_),
    .B(_13079_),
    .Y(_13828_));
 sky130_fd_sc_hd__nand2_1 _34833_ (.A(_13777_),
    .B(_02976_),
    .Y(_13829_));
 sky130_fd_sc_hd__nor3_1 _34834_ (.A(_13710_),
    .B(_13829_),
    .C(_13549_),
    .Y(_13830_));
 sky130_fd_sc_hd__o21ai_0 _34835_ (.A1(_13552_),
    .A2(_13828_),
    .B1(_13830_),
    .Y(_13831_));
 sky130_fd_sc_hd__nor2_1 _34836_ (.A(_13829_),
    .B(_13710_),
    .Y(_13832_));
 sky130_fd_sc_hd__a21oi_1 _34837_ (.A1(_13777_),
    .A2(_02555_),
    .B1(_01850_),
    .Y(_13833_));
 sky130_fd_sc_hd__o21ai_0 _34838_ (.A1(_13829_),
    .A2(_13713_),
    .B1(_13833_),
    .Y(_13834_));
 sky130_fd_sc_hd__a21oi_1 _34839_ (.A1(_13555_),
    .A2(_13832_),
    .B1(_13834_),
    .Y(_13835_));
 sky130_fd_sc_hd__inv_1 _34840_ (.A(_13416_),
    .Y(_13836_));
 sky130_fd_sc_hd__nor2_1 _34841_ (.A(_13068_),
    .B(_13546_),
    .Y(_13837_));
 sky130_fd_sc_hd__nand3_1 _34842_ (.A(_13836_),
    .B(_13830_),
    .C(_13837_),
    .Y(_13838_));
 sky130_fd_sc_hd__nand3_1 _34843_ (.A(_13831_),
    .B(_13835_),
    .C(_13838_),
    .Y(_13839_));
 sky130_fd_sc_hd__nand2_1 _34844_ (.A(_13839_),
    .B(net2008),
    .Y(_13840_));
 sky130_fd_sc_hd__o21ai_0 _34845_ (.A1(net2008),
    .A2(_13827_),
    .B1(_13840_),
    .Y(_13841_));
 sky130_fd_sc_hd__or2_2 _34846_ (.A(_13813_),
    .B(_13841_),
    .X(_13842_));
 sky130_fd_sc_hd__nand2_1 _34847_ (.A(_13841_),
    .B(_13813_),
    .Y(_13843_));
 sky130_fd_sc_hd__nand2_1 _34848_ (.A(_13842_),
    .B(_13843_),
    .Y(_13844_));
 sky130_fd_sc_hd__nand2_1 _34849_ (.A(_13844_),
    .B(net2214),
    .Y(_13845_));
 sky130_fd_sc_hd__nand2_1 _34850_ (.A(_13845_),
    .B(_05745_),
    .Y(_13846_));
 sky130_fd_sc_hd__nand2_1 _34851_ (.A(_13846_),
    .B(net2019),
    .Y(_13847_));
 sky130_fd_sc_hd__nand2_1 _34852_ (.A(net1798),
    .B(_03243_),
    .Y(_13848_));
 sky130_fd_sc_hd__nand2_1 _34853_ (.A(net1871),
    .B(_03242_),
    .Y(_13849_));
 sky130_fd_sc_hd__o211ai_1 _34854_ (.A1(_03246_),
    .A2(net1232),
    .B1(_13848_),
    .C1(_13849_),
    .Y(_13850_));
 sky130_fd_sc_hd__a21oi_1 _34856_ (.A1(_13850_),
    .A2(net2864),
    .B1(net2856),
    .Y(_13852_));
 sky130_fd_sc_hd__nand2_1 _34857_ (.A(\inst$top.soc.cpu.sink__payload$12[21] ),
    .B(\inst$top.soc.cpu.sink__payload$12[20] ),
    .Y(_13853_));
 sky130_fd_sc_hd__nor2_1 _34858_ (.A(_13853_),
    .B(_13693_),
    .Y(_13854_));
 sky130_fd_sc_hd__o21ai_0 _34859_ (.A1(_13853_),
    .A2(_13693_),
    .B1(\inst$top.soc.cpu.sink__payload$12[22] ),
    .Y(_13855_));
 sky130_fd_sc_hd__nand2_1 _34860_ (.A(_13855_),
    .B(net2854),
    .Y(_13856_));
 sky130_fd_sc_hd__a21oi_1 _34861_ (.A1(_12304_),
    .A2(_13854_),
    .B1(_13856_),
    .Y(_13857_));
 sky130_fd_sc_hd__a21oi_1 _34862_ (.A1(_13847_),
    .A2(_13852_),
    .B1(_13857_),
    .Y(_13858_));
 sky130_fd_sc_hd__nand2_1 _34863_ (.A(net603),
    .B(net786),
    .Y(_13859_));
 sky130_fd_sc_hd__o211ai_1 _34864_ (.A1(net785),
    .A2(_13811_),
    .B1(_13812_),
    .C1(_13859_),
    .Y(_13860_));
 sky130_fd_sc_hd__nor2_1 _34865_ (.A(net659),
    .B(_13860_),
    .Y(_13861_));
 sky130_fd_sc_hd__nor2_4 _34866_ (.A(_13801_),
    .B(_13861_),
    .Y(_04198_));
 sky130_fd_sc_hd__nand2_1 _34867_ (.A(\inst$top.soc.cpu.sink__payload$12[22] ),
    .B(\inst$top.soc.cpu.sink__payload$12[21] ),
    .Y(_13862_));
 sky130_fd_sc_hd__nor2_1 _34868_ (.A(_13788_),
    .B(_13862_),
    .Y(_13863_));
 sky130_fd_sc_hd__nand2_1 _34869_ (.A(_13611_),
    .B(_13863_),
    .Y(_13864_));
 sky130_fd_sc_hd__a21oi_1 _34870_ (.A1(_13864_),
    .A2(\inst$top.soc.cpu.sink__payload$12[23] ),
    .B1(net2001),
    .Y(_13865_));
 sky130_fd_sc_hd__nand3_1 _34871_ (.A(_13611_),
    .B(_05749_),
    .C(_13863_),
    .Y(_13866_));
 sky130_fd_sc_hd__nor2_1 _34872_ (.A(_02972_),
    .B(_13813_),
    .Y(_13867_));
 sky130_fd_sc_hd__inv_1 _34873_ (.A(_13867_),
    .Y(_13868_));
 sky130_fd_sc_hd__nor2_1 _34874_ (.A(_13758_),
    .B(_13868_),
    .Y(_13869_));
 sky130_fd_sc_hd__nand2_1 _34875_ (.A(_13626_),
    .B(_13869_),
    .Y(_13870_));
 sky130_fd_sc_hd__nand2_1 _34876_ (.A(_01850_),
    .B(_02966_),
    .Y(_13871_));
 sky130_fd_sc_hd__nand2_1 _34877_ (.A(_13871_),
    .B(_01957_),
    .Y(_13872_));
 sky130_fd_sc_hd__a21oi_1 _34878_ (.A1(_13761_),
    .A2(_13867_),
    .B1(_13872_),
    .Y(_13873_));
 sky130_fd_sc_hd__nand3_1 _34879_ (.A(_13870_),
    .B(net2006),
    .C(_13873_),
    .Y(_13874_));
 sky130_fd_sc_hd__nand2_1 _34880_ (.A(_13643_),
    .B(_13646_),
    .Y(_13875_));
 sky130_fd_sc_hd__nand2_1 _34881_ (.A(_13813_),
    .B(_02972_),
    .Y(_13876_));
 sky130_fd_sc_hd__nor2_1 _34882_ (.A(_13876_),
    .B(_13766_),
    .Y(_13877_));
 sky130_fd_sc_hd__nand2_1 _34883_ (.A(_13875_),
    .B(_13877_),
    .Y(_13878_));
 sky130_fd_sc_hd__nand2_1 _34884_ (.A(_13813_),
    .B(_02971_),
    .Y(_13879_));
 sky130_fd_sc_hd__inv_1 _34885_ (.A(_02968_),
    .Y(_13880_));
 sky130_fd_sc_hd__nand2_1 _34886_ (.A(_13879_),
    .B(_13880_),
    .Y(_13881_));
 sky130_fd_sc_hd__nor2_1 _34887_ (.A(_13876_),
    .B(_13771_),
    .Y(_13882_));
 sky130_fd_sc_hd__nor2_1 _34888_ (.A(_13881_),
    .B(_13882_),
    .Y(_13883_));
 sky130_fd_sc_hd__nand2_1 _34889_ (.A(_13878_),
    .B(_13883_),
    .Y(_13884_));
 sky130_fd_sc_hd__nand2_1 _34890_ (.A(_13884_),
    .B(net2865),
    .Y(_13885_));
 sky130_fd_sc_hd__nand2_1 _34891_ (.A(_13874_),
    .B(_13885_),
    .Y(_13886_));
 sky130_fd_sc_hd__nand2_1 _34892_ (.A(_13886_),
    .B(_02961_),
    .Y(_13887_));
 sky130_fd_sc_hd__inv_1 _34893_ (.A(_02961_),
    .Y(_13888_));
 sky130_fd_sc_hd__nand3_1 _34894_ (.A(_13874_),
    .B(_13885_),
    .C(_13888_),
    .Y(_13889_));
 sky130_fd_sc_hd__nand2_1 _34895_ (.A(_13887_),
    .B(_13889_),
    .Y(_13890_));
 sky130_fd_sc_hd__nand2_1 _34896_ (.A(_13890_),
    .B(net2215),
    .Y(_13891_));
 sky130_fd_sc_hd__nand2_1 _34897_ (.A(_13891_),
    .B(_05764_),
    .Y(_13892_));
 sky130_fd_sc_hd__nand2_1 _34898_ (.A(net1795),
    .B(_03250_),
    .Y(_13893_));
 sky130_fd_sc_hd__nand2_1 _34899_ (.A(net1868),
    .B(_03249_),
    .Y(_13894_));
 sky130_fd_sc_hd__o211ai_1 _34900_ (.A1(_03253_),
    .A2(net1229),
    .B1(_13893_),
    .C1(_13894_),
    .Y(_13895_));
 sky130_fd_sc_hd__a21oi_1 _34901_ (.A1(_13895_),
    .A2(net2862),
    .B1(net2854),
    .Y(_13896_));
 sky130_fd_sc_hd__a21boi_0 _34902_ (.A1(_13892_),
    .A2(net2017),
    .B1_N(_13896_),
    .Y(_13897_));
 sky130_fd_sc_hd__a21oi_4 _34903_ (.A1(_13865_),
    .A2(_13866_),
    .B1(_13897_),
    .Y(_13898_));
 sky130_fd_sc_hd__nand2_1 _34904_ (.A(_13898_),
    .B(net786),
    .Y(_13899_));
 sky130_fd_sc_hd__nand2_1 _34905_ (.A(net739),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[23] ),
    .Y(_13900_));
 sky130_fd_sc_hd__inv_1 _34906_ (.A(\inst$top.soc.cpu.sink__payload$18[132] ),
    .Y(_13901_));
 sky130_fd_sc_hd__nor2_1 _34907_ (.A(net2833),
    .B(_13901_),
    .Y(_13902_));
 sky130_fd_sc_hd__inv_1 _34908_ (.A(\inst$top.soc.cpu.shifter.m_result$7[23] ),
    .Y(_13903_));
 sky130_fd_sc_hd__o21ai_0 _34909_ (.A1(net2872),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[8] ),
    .B1(net2837),
    .Y(_13904_));
 sky130_fd_sc_hd__a21oi_1 _34910_ (.A1(net2872),
    .A2(_13903_),
    .B1(_13904_),
    .Y(_13905_));
 sky130_fd_sc_hd__o21ai_0 _34911_ (.A1(_13902_),
    .A2(_13905_),
    .B1(net2014),
    .Y(_13906_));
 sky130_fd_sc_hd__a21oi_1 _34912_ (.A1(_10622_),
    .A2(net2921),
    .B1(net2012),
    .Y(_13907_));
 sky130_fd_sc_hd__o21ai_1 _34913_ (.A1(net2921),
    .A2(\inst$top.soc.cpu.divider.quotient[23] ),
    .B1(_13907_),
    .Y(_13908_));
 sky130_fd_sc_hd__a21oi_1 _34914_ (.A1(_13906_),
    .A2(net1785),
    .B1(net2830),
    .Y(_13909_));
 sky130_fd_sc_hd__nand2_1 _34915_ (.A(_12984_),
    .B(_13909_),
    .Y(_13910_));
 sky130_fd_sc_hd__nand3_1 _34916_ (.A(_13899_),
    .B(_13900_),
    .C(_13910_),
    .Y(_13911_));
 sky130_fd_sc_hd__nor2_1 _34917_ (.A(net658),
    .B(_13911_),
    .Y(_13912_));
 sky130_fd_sc_hd__nand2_1 _34918_ (.A(net658),
    .B(_05750_),
    .Y(_13913_));
 sky130_fd_sc_hd__nand2_1 _34919_ (.A(_13913_),
    .B(net2181),
    .Y(_13914_));
 sky130_fd_sc_hd__nor2_4 _34920_ (.A(_13912_),
    .B(_13914_),
    .Y(_04199_));
 sky130_fd_sc_hd__nor2_1 _34921_ (.A(_02961_),
    .B(_02966_),
    .Y(_13915_));
 sky130_fd_sc_hd__inv_1 _34922_ (.A(_13915_),
    .Y(_13916_));
 sky130_fd_sc_hd__nor2_1 _34923_ (.A(_13916_),
    .B(_13817_),
    .Y(_13917_));
 sky130_fd_sc_hd__nand2_1 _34924_ (.A(_13917_),
    .B(_13701_),
    .Y(_13918_));
 sky130_fd_sc_hd__a21oi_2 _34925_ (.A1(_13888_),
    .A2(_02968_),
    .B1(_02963_),
    .Y(_13919_));
 sky130_fd_sc_hd__o21ai_0 _34926_ (.A1(_13916_),
    .A2(_13823_),
    .B1(_13919_),
    .Y(_13920_));
 sky130_fd_sc_hd__a21oi_1 _34927_ (.A1(_13706_),
    .A2(_13917_),
    .B1(_13920_),
    .Y(_13921_));
 sky130_fd_sc_hd__o21ai_0 _34928_ (.A1(_13918_),
    .A2(_13541_),
    .B1(_13921_),
    .Y(_13922_));
 sky130_fd_sc_hd__nand2_1 _34929_ (.A(_13922_),
    .B(net2865),
    .Y(_13923_));
 sky130_fd_sc_hd__nand2_1 _34930_ (.A(_02961_),
    .B(_02966_),
    .Y(_13924_));
 sky130_fd_sc_hd__nor2_1 _34931_ (.A(_13924_),
    .B(_13829_),
    .Y(_13925_));
 sky130_fd_sc_hd__a21oi_1 _34932_ (.A1(_01958_),
    .A2(_02961_),
    .B1(_02053_),
    .Y(_13926_));
 sky130_fd_sc_hd__o21ai_0 _34933_ (.A1(_13924_),
    .A2(_13833_),
    .B1(_13926_),
    .Y(_13927_));
 sky130_fd_sc_hd__a21oi_2 _34934_ (.A1(_13722_),
    .A2(_13925_),
    .B1(_13927_),
    .Y(_13928_));
 sky130_fd_sc_hd__nand2_1 _34935_ (.A(_13928_),
    .B(net2007),
    .Y(_13929_));
 sky130_fd_sc_hd__nand2_1 _34936_ (.A(_13923_),
    .B(_13929_),
    .Y(_13930_));
 sky130_fd_sc_hd__inv_1 _34937_ (.A(_02957_),
    .Y(_13931_));
 sky130_fd_sc_hd__nand2_1 _34938_ (.A(_13930_),
    .B(_13931_),
    .Y(_13932_));
 sky130_fd_sc_hd__nand3_1 _34939_ (.A(_13923_),
    .B(_13929_),
    .C(_02957_),
    .Y(_13933_));
 sky130_fd_sc_hd__nand2_1 _34940_ (.A(_13932_),
    .B(_13933_),
    .Y(_13934_));
 sky130_fd_sc_hd__nand2_1 _34941_ (.A(_13934_),
    .B(net2215),
    .Y(_13935_));
 sky130_fd_sc_hd__nand2_1 _34942_ (.A(_13935_),
    .B(_05785_),
    .Y(_13936_));
 sky130_fd_sc_hd__nand2_1 _34943_ (.A(_13936_),
    .B(net2020),
    .Y(_13937_));
 sky130_fd_sc_hd__nand2_1 _34944_ (.A(net1795),
    .B(_03257_),
    .Y(_13938_));
 sky130_fd_sc_hd__nand2_1 _34945_ (.A(net1869),
    .B(_03256_),
    .Y(_13939_));
 sky130_fd_sc_hd__o211ai_1 _34946_ (.A1(_03260_),
    .A2(net1229),
    .B1(_13938_),
    .C1(_13939_),
    .Y(_13940_));
 sky130_fd_sc_hd__a21oi_1 _34947_ (.A1(_13940_),
    .A2(net2862),
    .B1(net2854),
    .Y(_13941_));
 sky130_fd_sc_hd__nand2_1 _34948_ (.A(\inst$top.soc.cpu.sink__payload$12[23] ),
    .B(\inst$top.soc.cpu.sink__payload$12[22] ),
    .Y(_13942_));
 sky130_fd_sc_hd__nor4_1 _34949_ (.A(\inst$top.soc.cpu.sink__payload$12[24] ),
    .B(_13853_),
    .C(_13942_),
    .D(_13693_),
    .Y(_13943_));
 sky130_fd_sc_hd__inv_1 _34950_ (.A(_13942_),
    .Y(_13944_));
 sky130_fd_sc_hd__a21oi_1 _34951_ (.A1(_13854_),
    .A2(_13944_),
    .B1(_05768_),
    .Y(_13945_));
 sky130_fd_sc_hd__nor3_1 _34952_ (.A(net2001),
    .B(_13943_),
    .C(_13945_),
    .Y(_13946_));
 sky130_fd_sc_hd__a21oi_4 _34953_ (.A1(_13937_),
    .A2(_13941_),
    .B1(_13946_),
    .Y(_13947_));
 sky130_fd_sc_hd__nand2_1 _34954_ (.A(_13947_),
    .B(net786),
    .Y(_13948_));
 sky130_fd_sc_hd__nand2_1 _34955_ (.A(net739),
    .B(net938),
    .Y(_13949_));
 sky130_fd_sc_hd__inv_1 _34956_ (.A(\inst$top.soc.cpu.sink__payload$18[133] ),
    .Y(_13950_));
 sky130_fd_sc_hd__nor2_1 _34957_ (.A(net2840),
    .B(_13950_),
    .Y(_13951_));
 sky130_fd_sc_hd__inv_1 _34958_ (.A(\inst$top.soc.cpu.shifter.m_result$7[24] ),
    .Y(_13952_));
 sky130_fd_sc_hd__o21ai_0 _34959_ (.A1(net2871),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[7] ),
    .B1(net2840),
    .Y(_13953_));
 sky130_fd_sc_hd__a21oi_1 _34960_ (.A1(net2871),
    .A2(_13952_),
    .B1(_13953_),
    .Y(_13954_));
 sky130_fd_sc_hd__o21ai_0 _34961_ (.A1(_13951_),
    .A2(_13954_),
    .B1(net2015),
    .Y(_13955_));
 sky130_fd_sc_hd__a21oi_1 _34962_ (.A1(_10638_),
    .A2(net2921),
    .B1(net2011),
    .Y(_13956_));
 sky130_fd_sc_hd__o21ai_1 _34963_ (.A1(net2921),
    .A2(\inst$top.soc.cpu.divider.quotient[24] ),
    .B1(_13956_),
    .Y(_13957_));
 sky130_fd_sc_hd__a21oi_1 _34964_ (.A1(_13955_),
    .A2(net1784),
    .B1(net2831),
    .Y(_13958_));
 sky130_fd_sc_hd__nand2_1 _34965_ (.A(_12984_),
    .B(_13958_),
    .Y(_13959_));
 sky130_fd_sc_hd__nand3_1 _34966_ (.A(_13948_),
    .B(_13949_),
    .C(_13959_),
    .Y(_13960_));
 sky130_fd_sc_hd__nand2_1 _34967_ (.A(net713),
    .B(_13960_),
    .Y(_13961_));
 sky130_fd_sc_hd__nand2_1 _34968_ (.A(net658),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[24] ),
    .Y(_13962_));
 sky130_fd_sc_hd__a21oi_4 _34969_ (.A1(_13961_),
    .A2(_13962_),
    .B1(net3010),
    .Y(_04200_));
 sky130_fd_sc_hd__nand2_1 _34970_ (.A(net660),
    .B(_05789_),
    .Y(_13963_));
 sky130_fd_sc_hd__nand2_1 _34971_ (.A(_13963_),
    .B(net2156),
    .Y(_13964_));
 sky130_fd_sc_hd__nand2_1 _34972_ (.A(\inst$top.soc.cpu.sink__payload$12[24] ),
    .B(\inst$top.soc.cpu.sink__payload$12[23] ),
    .Y(_13965_));
 sky130_fd_sc_hd__o31ai_1 _34973_ (.A1(_13862_),
    .A2(_13965_),
    .A3(_13790_),
    .B1(\inst$top.soc.cpu.sink__payload$12[25] ),
    .Y(_13966_));
 sky130_fd_sc_hd__o41ai_1 _34974_ (.A1(\inst$top.soc.cpu.sink__payload$12[25] ),
    .A2(_13862_),
    .A3(_13965_),
    .A4(_13790_),
    .B1(net2855),
    .Y(_13967_));
 sky130_fd_sc_hd__inv_1 _34975_ (.A(_13967_),
    .Y(_13968_));
 sky130_fd_sc_hd__nor2_1 _34976_ (.A(_02957_),
    .B(_13888_),
    .Y(_13969_));
 sky130_fd_sc_hd__nand2_1 _34977_ (.A(_13867_),
    .B(_13969_),
    .Y(_13970_));
 sky130_fd_sc_hd__inv_1 _34978_ (.A(_13970_),
    .Y(_13971_));
 sky130_fd_sc_hd__nand2_1 _34979_ (.A(_13763_),
    .B(_13971_),
    .Y(_13972_));
 sky130_fd_sc_hd__o21ai_0 _34980_ (.A1(_02957_),
    .A2(_02052_),
    .B1(_02130_),
    .Y(_13973_));
 sky130_fd_sc_hd__a21oi_1 _34981_ (.A1(_13872_),
    .A2(_13969_),
    .B1(_13973_),
    .Y(_13974_));
 sky130_fd_sc_hd__nand3_1 _34982_ (.A(_13972_),
    .B(net2007),
    .C(_13974_),
    .Y(_13975_));
 sky130_fd_sc_hd__nand3_1 _34983_ (.A(_13768_),
    .B(_13774_),
    .C(_13769_),
    .Y(_13976_));
 sky130_fd_sc_hd__nor2_1 _34984_ (.A(_02961_),
    .B(_13931_),
    .Y(_13977_));
 sky130_fd_sc_hd__inv_1 _34985_ (.A(_13977_),
    .Y(_13978_));
 sky130_fd_sc_hd__nor2_1 _34986_ (.A(_13876_),
    .B(_13978_),
    .Y(_13979_));
 sky130_fd_sc_hd__nand2_1 _34987_ (.A(_13976_),
    .B(_13979_),
    .Y(_13980_));
 sky130_fd_sc_hd__a21oi_1 _34988_ (.A1(_02957_),
    .A2(_02963_),
    .B1(_02956_),
    .Y(_13981_));
 sky130_fd_sc_hd__inv_1 _34989_ (.A(_13981_),
    .Y(_13982_));
 sky130_fd_sc_hd__a21oi_1 _34990_ (.A1(_13881_),
    .A2(_13977_),
    .B1(_13982_),
    .Y(_13983_));
 sky130_fd_sc_hd__nand2_1 _34991_ (.A(_13980_),
    .B(_13983_),
    .Y(_13984_));
 sky130_fd_sc_hd__nand2_1 _34992_ (.A(_13984_),
    .B(net2866),
    .Y(_13985_));
 sky130_fd_sc_hd__nand2_1 _34993_ (.A(_13975_),
    .B(_13985_),
    .Y(_13986_));
 sky130_fd_sc_hd__nand2_1 _34994_ (.A(_13986_),
    .B(_02952_),
    .Y(_13987_));
 sky130_fd_sc_hd__inv_1 _34995_ (.A(_02952_),
    .Y(_13988_));
 sky130_fd_sc_hd__nand3_1 _34996_ (.A(_13975_),
    .B(_13988_),
    .C(_13985_),
    .Y(_13989_));
 sky130_fd_sc_hd__nand2_1 _34997_ (.A(_13987_),
    .B(_13989_),
    .Y(_13990_));
 sky130_fd_sc_hd__o21ai_0 _34998_ (.A1(net2843),
    .A2(_13990_),
    .B1(_05804_),
    .Y(_13991_));
 sky130_fd_sc_hd__nand2_1 _34999_ (.A(_13991_),
    .B(net2019),
    .Y(_13992_));
 sky130_fd_sc_hd__nand2_1 _35000_ (.A(net1796),
    .B(_03264_),
    .Y(_13993_));
 sky130_fd_sc_hd__nand2_1 _35001_ (.A(net1869),
    .B(_03263_),
    .Y(_13994_));
 sky130_fd_sc_hd__o211ai_1 _35002_ (.A1(_03267_),
    .A2(net1230),
    .B1(_13993_),
    .C1(_13994_),
    .Y(_13995_));
 sky130_fd_sc_hd__a21oi_1 _35003_ (.A1(_13995_),
    .A2(net2864),
    .B1(net2856),
    .Y(_13996_));
 sky130_fd_sc_hd__a22oi_1 _35004_ (.A1(_13966_),
    .A2(_13968_),
    .B1(_13992_),
    .B2(_13996_),
    .Y(_13997_));
 sky130_fd_sc_hd__nand2_1 _35005_ (.A(_13997_),
    .B(net787),
    .Y(_13998_));
 sky130_fd_sc_hd__nand2_1 _35006_ (.A(net738),
    .B(net933),
    .Y(_13999_));
 sky130_fd_sc_hd__inv_1 _35007_ (.A(\inst$top.soc.cpu.sink__payload$18[134] ),
    .Y(_14000_));
 sky130_fd_sc_hd__nor2_1 _35008_ (.A(net2833),
    .B(_14000_),
    .Y(_14001_));
 sky130_fd_sc_hd__inv_1 _35009_ (.A(\inst$top.soc.cpu.shifter.m_result$7[25] ),
    .Y(_14002_));
 sky130_fd_sc_hd__o21ai_0 _35010_ (.A1(net2872),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[6] ),
    .B1(net2837),
    .Y(_14003_));
 sky130_fd_sc_hd__a21oi_1 _35011_ (.A1(net2872),
    .A2(_14002_),
    .B1(_14003_),
    .Y(_14004_));
 sky130_fd_sc_hd__o21ai_0 _35012_ (.A1(_14001_),
    .A2(_14004_),
    .B1(net2016),
    .Y(_14005_));
 sky130_fd_sc_hd__a21oi_1 _35013_ (.A1(_10655_),
    .A2(net2922),
    .B1(net2012),
    .Y(_14006_));
 sky130_fd_sc_hd__o21ai_2 _35014_ (.A1(net2922),
    .A2(\inst$top.soc.cpu.divider.quotient[25] ),
    .B1(_14006_),
    .Y(_14007_));
 sky130_fd_sc_hd__a21oi_1 _35015_ (.A1(_14005_),
    .A2(_14007_),
    .B1(net2832),
    .Y(_14008_));
 sky130_fd_sc_hd__nand2_1 _35016_ (.A(_12984_),
    .B(_14008_),
    .Y(_14009_));
 sky130_fd_sc_hd__nand3_1 _35017_ (.A(_13998_),
    .B(_13999_),
    .C(_14009_),
    .Y(_14010_));
 sky130_fd_sc_hd__nor2_1 _35018_ (.A(net657),
    .B(_14010_),
    .Y(_14011_));
 sky130_fd_sc_hd__nor2_4 _35019_ (.A(_13964_),
    .B(_14011_),
    .Y(_04201_));
 sky130_fd_sc_hd__inv_1 _35020_ (.A(\inst$top.soc.cpu.sink__payload$18[135] ),
    .Y(_14012_));
 sky130_fd_sc_hd__nor2_1 _35021_ (.A(net2834),
    .B(_14012_),
    .Y(_14013_));
 sky130_fd_sc_hd__inv_1 _35022_ (.A(\inst$top.soc.cpu.shifter.m_result$7[26] ),
    .Y(_14014_));
 sky130_fd_sc_hd__o21ai_0 _35023_ (.A1(net2870),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[5] ),
    .B1(net2836),
    .Y(_14015_));
 sky130_fd_sc_hd__a21oi_1 _35024_ (.A1(net2870),
    .A2(_14014_),
    .B1(_14015_),
    .Y(_14016_));
 sky130_fd_sc_hd__o21ai_0 _35025_ (.A1(_14013_),
    .A2(_14016_),
    .B1(net2013),
    .Y(_14017_));
 sky130_fd_sc_hd__a21oi_1 _35026_ (.A1(_10668_),
    .A2(net2922),
    .B1(net2012),
    .Y(_14018_));
 sky130_fd_sc_hd__o21ai_2 _35027_ (.A1(net2922),
    .A2(\inst$top.soc.cpu.divider.quotient[26] ),
    .B1(_14018_),
    .Y(_14019_));
 sky130_fd_sc_hd__a21oi_1 _35028_ (.A1(_14017_),
    .A2(_14019_),
    .B1(net2829),
    .Y(_14020_));
 sky130_fd_sc_hd__inv_1 _35029_ (.A(_14020_),
    .Y(_14021_));
 sky130_fd_sc_hd__nand2_1 _35030_ (.A(net737),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[26] ),
    .Y(_14022_));
 sky130_fd_sc_hd__nor2_1 _35031_ (.A(_13318_),
    .B(_13815_),
    .Y(_14023_));
 sky130_fd_sc_hd__nand2_1 _35032_ (.A(_02952_),
    .B(_02957_),
    .Y(_14024_));
 sky130_fd_sc_hd__nor3_1 _35033_ (.A(_13916_),
    .B(_14024_),
    .C(_13819_),
    .Y(_14025_));
 sky130_fd_sc_hd__nand3_1 _35034_ (.A(_13058_),
    .B(_14023_),
    .C(_14025_),
    .Y(_14026_));
 sky130_fd_sc_hd__nor2_1 _35035_ (.A(_14024_),
    .B(_13916_),
    .Y(_14027_));
 sky130_fd_sc_hd__a21oi_1 _35036_ (.A1(_02952_),
    .A2(_02956_),
    .B1(_02951_),
    .Y(_14028_));
 sky130_fd_sc_hd__o21ai_0 _35037_ (.A1(_14024_),
    .A2(_13919_),
    .B1(_14028_),
    .Y(_14029_));
 sky130_fd_sc_hd__a21oi_1 _35038_ (.A1(_13824_),
    .A2(_14027_),
    .B1(_14029_),
    .Y(_14030_));
 sky130_fd_sc_hd__nor2_1 _35039_ (.A(_13815_),
    .B(_13315_),
    .Y(_14031_));
 sky130_fd_sc_hd__o21ai_0 _35040_ (.A1(_13822_),
    .A2(_14031_),
    .B1(_14025_),
    .Y(_14032_));
 sky130_fd_sc_hd__nand3_1 _35041_ (.A(_14026_),
    .B(_14030_),
    .C(_14032_),
    .Y(_14033_));
 sky130_fd_sc_hd__nand2_1 _35042_ (.A(_14033_),
    .B(net2867),
    .Y(_14034_));
 sky130_fd_sc_hd__nor2_1 _35043_ (.A(_02952_),
    .B(_02957_),
    .Y(_14035_));
 sky130_fd_sc_hd__inv_1 _35044_ (.A(_14035_),
    .Y(_14036_));
 sky130_fd_sc_hd__nor2_1 _35045_ (.A(_13924_),
    .B(_14036_),
    .Y(_14037_));
 sky130_fd_sc_hd__nand2_1 _35046_ (.A(_13839_),
    .B(_14037_),
    .Y(_14038_));
 sky130_fd_sc_hd__a21oi_1 _35047_ (.A1(_13988_),
    .A2(_02603_),
    .B1(_02616_),
    .Y(_14039_));
 sky130_fd_sc_hd__o21ai_0 _35048_ (.A1(_14036_),
    .A2(_13926_),
    .B1(_14039_),
    .Y(_14040_));
 sky130_fd_sc_hd__nor2_1 _35049_ (.A(\inst$top.soc.cpu.adder$307.x_sub ),
    .B(_14040_),
    .Y(_14041_));
 sky130_fd_sc_hd__nand2_1 _35050_ (.A(_14038_),
    .B(_14041_),
    .Y(_14042_));
 sky130_fd_sc_hd__nand2_1 _35051_ (.A(_14034_),
    .B(_14042_),
    .Y(_14043_));
 sky130_fd_sc_hd__nand2_1 _35052_ (.A(_14043_),
    .B(_02947_),
    .Y(_14044_));
 sky130_fd_sc_hd__nand3b_1 _35053_ (.A_N(_02947_),
    .B(_14034_),
    .C(_14042_),
    .Y(_14045_));
 sky130_fd_sc_hd__nand2_1 _35054_ (.A(_14044_),
    .B(_14045_),
    .Y(_14046_));
 sky130_fd_sc_hd__o21ai_0 _35055_ (.A1(net2849),
    .A2(_14046_),
    .B1(_05822_),
    .Y(_14047_));
 sky130_fd_sc_hd__nand2_1 _35056_ (.A(_14047_),
    .B(net2019),
    .Y(_14048_));
 sky130_fd_sc_hd__nand2_1 _35057_ (.A(net1798),
    .B(_03271_),
    .Y(_14049_));
 sky130_fd_sc_hd__nand2_1 _35058_ (.A(net1871),
    .B(_03270_),
    .Y(_14050_));
 sky130_fd_sc_hd__o211ai_1 _35059_ (.A1(_03274_),
    .A2(net1232),
    .B1(_14049_),
    .C1(_14050_),
    .Y(_14051_));
 sky130_fd_sc_hd__a21oi_1 _35060_ (.A1(_14051_),
    .A2(net2863),
    .B1(net2855),
    .Y(_14052_));
 sky130_fd_sc_hd__nand4_1 _35061_ (.A(_13854_),
    .B(\inst$top.soc.cpu.sink__payload$12[25] ),
    .C(\inst$top.soc.cpu.sink__payload$12[24] ),
    .D(_13944_),
    .Y(_14053_));
 sky130_fd_sc_hd__inv_1 _35062_ (.A(_14053_),
    .Y(_14054_));
 sky130_fd_sc_hd__nand2_1 _35063_ (.A(_14054_),
    .B(\inst$top.soc.cpu.sink__payload$12[26] ),
    .Y(_14055_));
 sky130_fd_sc_hd__nand2_1 _35064_ (.A(_14053_),
    .B(_12420_),
    .Y(_14056_));
 sky130_fd_sc_hd__a21oi_1 _35065_ (.A1(_14055_),
    .A2(_14056_),
    .B1(net2001),
    .Y(_14057_));
 sky130_fd_sc_hd__a21oi_1 _35066_ (.A1(_14048_),
    .A2(_14052_),
    .B1(_14057_),
    .Y(_14058_));
 sky130_fd_sc_hd__nand2_1 _35067_ (.A(_14058_),
    .B(net787),
    .Y(_14059_));
 sky130_fd_sc_hd__o211ai_1 _35068_ (.A1(net783),
    .A2(_14021_),
    .B1(_14022_),
    .C1(_14059_),
    .Y(_14060_));
 sky130_fd_sc_hd__nand2_1 _35069_ (.A(net705),
    .B(_14060_),
    .Y(_14061_));
 sky130_fd_sc_hd__nand2_1 _35071_ (.A(net652),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[26] ),
    .Y(_14063_));
 sky130_fd_sc_hd__a21oi_4 _35072_ (.A1(_14061_),
    .A2(_14063_),
    .B1(net2993),
    .Y(_04202_));
 sky130_fd_sc_hd__nand2_1 _35073_ (.A(net660),
    .B(_19948_),
    .Y(_14064_));
 sky130_fd_sc_hd__nand2_1 _35074_ (.A(_14064_),
    .B(net2175),
    .Y(_14065_));
 sky130_fd_sc_hd__inv_1 _35075_ (.A(\inst$top.soc.cpu.sink__payload$18[136] ),
    .Y(_14066_));
 sky130_fd_sc_hd__nor2_1 _35076_ (.A(net2834),
    .B(_14066_),
    .Y(_14067_));
 sky130_fd_sc_hd__inv_1 _35077_ (.A(\inst$top.soc.cpu.shifter.m_result$7[27] ),
    .Y(_14068_));
 sky130_fd_sc_hd__o21ai_0 _35078_ (.A1(net2869),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[4] ),
    .B1(net2836),
    .Y(_14069_));
 sky130_fd_sc_hd__a21oi_1 _35079_ (.A1(net2869),
    .A2(_14068_),
    .B1(_14069_),
    .Y(_14070_));
 sky130_fd_sc_hd__o21ai_0 _35080_ (.A1(_14067_),
    .A2(_14070_),
    .B1(net2013),
    .Y(_14071_));
 sky130_fd_sc_hd__a21oi_1 _35081_ (.A1(_10699_),
    .A2(net2924),
    .B1(net2012),
    .Y(_14072_));
 sky130_fd_sc_hd__o21ai_2 _35082_ (.A1(net2921),
    .A2(\inst$top.soc.cpu.divider.quotient[27] ),
    .B1(_14072_),
    .Y(_14073_));
 sky130_fd_sc_hd__a21oi_1 _35083_ (.A1(_14071_),
    .A2(_14073_),
    .B1(net2829),
    .Y(_14074_));
 sky130_fd_sc_hd__inv_1 _35084_ (.A(_14074_),
    .Y(_14075_));
 sky130_fd_sc_hd__nand2_1 _35085_ (.A(net738),
    .B(net924),
    .Y(_14076_));
 sky130_fd_sc_hd__inv_1 _35086_ (.A(_02943_),
    .Y(_14077_));
 sky130_fd_sc_hd__inv_1 _35087_ (.A(_13877_),
    .Y(_14078_));
 sky130_fd_sc_hd__nand2_1 _35088_ (.A(_02947_),
    .B(_02952_),
    .Y(_14079_));
 sky130_fd_sc_hd__nor2_1 _35089_ (.A(_14079_),
    .B(_13978_),
    .Y(_14080_));
 sky130_fd_sc_hd__inv_1 _35090_ (.A(_14080_),
    .Y(_14081_));
 sky130_fd_sc_hd__nor2_1 _35091_ (.A(_14078_),
    .B(_14081_),
    .Y(_14082_));
 sky130_fd_sc_hd__nand3_1 _35092_ (.A(_13184_),
    .B(_13638_),
    .C(_14082_),
    .Y(_14083_));
 sky130_fd_sc_hd__nand2_1 _35093_ (.A(_02947_),
    .B(_02951_),
    .Y(_14084_));
 sky130_fd_sc_hd__inv_1 _35094_ (.A(_02946_),
    .Y(_14085_));
 sky130_fd_sc_hd__nand2_1 _35095_ (.A(_14084_),
    .B(_14085_),
    .Y(_14086_));
 sky130_fd_sc_hd__a31oi_1 _35096_ (.A1(_13982_),
    .A2(_02947_),
    .A3(_02952_),
    .B1(_14086_),
    .Y(_14087_));
 sky130_fd_sc_hd__o21ai_0 _35097_ (.A1(_14081_),
    .A2(_13883_),
    .B1(_14087_),
    .Y(_14088_));
 sky130_fd_sc_hd__a21oi_1 _35098_ (.A1(_13642_),
    .A2(_14082_),
    .B1(_14088_),
    .Y(_14089_));
 sky130_fd_sc_hd__nand2_1 _35099_ (.A(_14083_),
    .B(_14089_),
    .Y(_14090_));
 sky130_fd_sc_hd__a21oi_1 _35100_ (.A1(_14090_),
    .A2(_14077_),
    .B1(net2005),
    .Y(_14091_));
 sky130_fd_sc_hd__o21ai_0 _35101_ (.A1(_14077_),
    .A2(_14090_),
    .B1(_14091_),
    .Y(_14092_));
 sky130_fd_sc_hd__inv_1 _35102_ (.A(_02918_),
    .Y(_14093_));
 sky130_fd_sc_hd__nor2_1 _35103_ (.A(_02947_),
    .B(_02952_),
    .Y(_14094_));
 sky130_fd_sc_hd__nand2_1 _35104_ (.A(_13969_),
    .B(_14094_),
    .Y(_14095_));
 sky130_fd_sc_hd__nor3_1 _35105_ (.A(_13758_),
    .B(_13868_),
    .C(_14095_),
    .Y(_14096_));
 sky130_fd_sc_hd__nand3_1 _35106_ (.A(_13158_),
    .B(_13623_),
    .C(_14096_),
    .Y(_14097_));
 sky130_fd_sc_hd__inv_1 _35107_ (.A(_02257_),
    .Y(_14098_));
 sky130_fd_sc_hd__o21ai_0 _35108_ (.A1(_02947_),
    .A2(_02196_),
    .B1(_14098_),
    .Y(_14099_));
 sky130_fd_sc_hd__a21oi_1 _35109_ (.A1(_13973_),
    .A2(_14094_),
    .B1(_14099_),
    .Y(_14100_));
 sky130_fd_sc_hd__o21ai_0 _35110_ (.A1(_14095_),
    .A2(_13873_),
    .B1(_14100_),
    .Y(_14101_));
 sky130_fd_sc_hd__a21oi_1 _35111_ (.A1(_13621_),
    .A2(_14096_),
    .B1(_14101_),
    .Y(_14102_));
 sky130_fd_sc_hd__nand2_1 _35112_ (.A(_14097_),
    .B(_14102_),
    .Y(_14103_));
 sky130_fd_sc_hd__o21ai_0 _35113_ (.A1(_14093_),
    .A2(_14103_),
    .B1(net2007),
    .Y(_14104_));
 sky130_fd_sc_hd__a21o_1 _35114_ (.A1(_14093_),
    .A2(_14103_),
    .B1(_14104_),
    .X(_14105_));
 sky130_fd_sc_hd__nand3_1 _35115_ (.A(_14092_),
    .B(net2215),
    .C(_14105_),
    .Y(_14106_));
 sky130_fd_sc_hd__nand2_1 _35116_ (.A(_14106_),
    .B(_05835_),
    .Y(_14107_));
 sky130_fd_sc_hd__nand2_1 _35117_ (.A(_14107_),
    .B(net2020),
    .Y(_14108_));
 sky130_fd_sc_hd__nand2_1 _35118_ (.A(net1796),
    .B(_03278_),
    .Y(_14109_));
 sky130_fd_sc_hd__nand2_1 _35119_ (.A(net1869),
    .B(_03277_),
    .Y(_14110_));
 sky130_fd_sc_hd__o211ai_1 _35120_ (.A1(_03281_),
    .A2(net1230),
    .B1(_14109_),
    .C1(_14110_),
    .Y(_14111_));
 sky130_fd_sc_hd__a21oi_1 _35121_ (.A1(_14111_),
    .A2(net2863),
    .B1(net2856),
    .Y(_14112_));
 sky130_fd_sc_hd__nor3_1 _35122_ (.A(_12420_),
    .B(_12384_),
    .C(_13965_),
    .Y(_14113_));
 sky130_fd_sc_hd__inv_1 _35123_ (.A(_14113_),
    .Y(_14114_));
 sky130_fd_sc_hd__nor2_1 _35124_ (.A(_14114_),
    .B(_13864_),
    .Y(_14115_));
 sky130_fd_sc_hd__o21ai_0 _35125_ (.A1(_19947_),
    .A2(_14115_),
    .B1(net2854),
    .Y(_14116_));
 sky130_fd_sc_hd__a41oi_1 _35126_ (.A1(_19947_),
    .A2(_13611_),
    .A3(_13863_),
    .A4(_14113_),
    .B1(_14116_),
    .Y(_14117_));
 sky130_fd_sc_hd__a21oi_2 _35127_ (.A1(_14108_),
    .A2(_14112_),
    .B1(_14117_),
    .Y(_14118_));
 sky130_fd_sc_hd__nand2_1 _35128_ (.A(_14118_),
    .B(net787),
    .Y(_14119_));
 sky130_fd_sc_hd__o211ai_1 _35129_ (.A1(net783),
    .A2(_14075_),
    .B1(_14076_),
    .C1(_14119_),
    .Y(_14120_));
 sky130_fd_sc_hd__nor2_1 _35130_ (.A(net656),
    .B(_14120_),
    .Y(_14121_));
 sky130_fd_sc_hd__nor2_4 _35131_ (.A(_14065_),
    .B(_14121_),
    .Y(_04203_));
 sky130_fd_sc_hd__nor2_1 _35132_ (.A(_02947_),
    .B(_14093_),
    .Y(_14122_));
 sky130_fd_sc_hd__inv_1 _35133_ (.A(_14122_),
    .Y(_14123_));
 sky130_fd_sc_hd__nor2_1 _35134_ (.A(_14036_),
    .B(_14123_),
    .Y(_14124_));
 sky130_fd_sc_hd__nand2_1 _35135_ (.A(_13927_),
    .B(_14124_),
    .Y(_14125_));
 sky130_fd_sc_hd__o21ai_0 _35136_ (.A1(_14098_),
    .A2(_14093_),
    .B1(_02324_),
    .Y(_14126_));
 sky130_fd_sc_hd__nor2_1 _35137_ (.A(_14123_),
    .B(_14039_),
    .Y(_14127_));
 sky130_fd_sc_hd__nor2_1 _35138_ (.A(_14126_),
    .B(_14127_),
    .Y(_14128_));
 sky130_fd_sc_hd__nand2_1 _35139_ (.A(_14125_),
    .B(_14128_),
    .Y(_14129_));
 sky130_fd_sc_hd__a31oi_1 _35140_ (.A1(_13715_),
    .A2(_13925_),
    .A3(_14124_),
    .B1(_14129_),
    .Y(_14130_));
 sky130_fd_sc_hd__and3_1 _35141_ (.A(_13718_),
    .B(_13925_),
    .C(_14124_),
    .X(_14131_));
 sky130_fd_sc_hd__nand2_1 _35142_ (.A(_13202_),
    .B(_14131_),
    .Y(_14132_));
 sky130_fd_sc_hd__nand2_1 _35143_ (.A(_14130_),
    .B(_14132_),
    .Y(_14133_));
 sky130_fd_sc_hd__xor2_1 _35144_ (.A(_02938_),
    .B(_14133_),
    .X(_14134_));
 sky130_fd_sc_hd__nand2_1 _35145_ (.A(_14134_),
    .B(net2005),
    .Y(_14135_));
 sky130_fd_sc_hd__inv_1 _35146_ (.A(_02938_),
    .Y(_14136_));
 sky130_fd_sc_hd__nand2_1 _35147_ (.A(_02947_),
    .B(_02943_),
    .Y(_14137_));
 sky130_fd_sc_hd__nor4_1 _35148_ (.A(_14024_),
    .B(_14137_),
    .C(_13916_),
    .D(_13817_),
    .Y(_14138_));
 sky130_fd_sc_hd__nand4_1 _35149_ (.A(_13213_),
    .B(_13434_),
    .C(_13703_),
    .D(_14138_),
    .Y(_14139_));
 sky130_fd_sc_hd__nor2_1 _35150_ (.A(_14024_),
    .B(_14137_),
    .Y(_14140_));
 sky130_fd_sc_hd__a21oi_1 _35151_ (.A1(_02946_),
    .A2(_02943_),
    .B1(_02942_),
    .Y(_14141_));
 sky130_fd_sc_hd__o21ai_0 _35152_ (.A1(_14137_),
    .A2(_14028_),
    .B1(_14141_),
    .Y(_14142_));
 sky130_fd_sc_hd__a21oi_1 _35153_ (.A1(_13920_),
    .A2(_14140_),
    .B1(_14142_),
    .Y(_14143_));
 sky130_fd_sc_hd__nand2_1 _35154_ (.A(_13440_),
    .B(_13703_),
    .Y(_14144_));
 sky130_fd_sc_hd__nand2_1 _35155_ (.A(_14144_),
    .B(_13707_),
    .Y(_14145_));
 sky130_fd_sc_hd__nand2_1 _35156_ (.A(_14145_),
    .B(_14138_),
    .Y(_14146_));
 sky130_fd_sc_hd__nand3_1 _35157_ (.A(_14139_),
    .B(_14143_),
    .C(_14146_),
    .Y(_14147_));
 sky130_fd_sc_hd__xor2_1 _35158_ (.A(_14136_),
    .B(_14147_),
    .X(_14148_));
 sky130_fd_sc_hd__nand2_1 _35159_ (.A(_14148_),
    .B(net2868),
    .Y(_14149_));
 sky130_fd_sc_hd__nand2_1 _35160_ (.A(_14135_),
    .B(_14149_),
    .Y(_14150_));
 sky130_fd_sc_hd__nand2_1 _35161_ (.A(_14150_),
    .B(net2214),
    .Y(_14151_));
 sky130_fd_sc_hd__nand2_1 _35162_ (.A(_14151_),
    .B(_05847_),
    .Y(_14152_));
 sky130_fd_sc_hd__nand2_1 _35163_ (.A(_14152_),
    .B(net2019),
    .Y(_14153_));
 sky130_fd_sc_hd__nand2_1 _35164_ (.A(net1798),
    .B(_03285_),
    .Y(_14154_));
 sky130_fd_sc_hd__nand2_1 _35165_ (.A(net1871),
    .B(_03284_),
    .Y(_14155_));
 sky130_fd_sc_hd__o211ai_1 _35166_ (.A1(_03288_),
    .A2(net1232),
    .B1(_14154_),
    .C1(_14155_),
    .Y(_14156_));
 sky130_fd_sc_hd__a21oi_1 _35167_ (.A1(_14156_),
    .A2(net2863),
    .B1(net2856),
    .Y(_14157_));
 sky130_fd_sc_hd__nor4_1 _35168_ (.A(\inst$top.soc.cpu.sink__payload$12[28] ),
    .B(_19947_),
    .C(_12420_),
    .D(_14053_),
    .Y(_14158_));
 sky130_fd_sc_hd__a31oi_1 _35169_ (.A1(_14054_),
    .A2(\inst$top.soc.cpu.sink__payload$12[27] ),
    .A3(\inst$top.soc.cpu.sink__payload$12[26] ),
    .B1(_12481_),
    .Y(_14159_));
 sky130_fd_sc_hd__nor3_1 _35170_ (.A(net2001),
    .B(_14158_),
    .C(_14159_),
    .Y(_14160_));
 sky130_fd_sc_hd__a21oi_4 _35171_ (.A1(_14153_),
    .A2(_14157_),
    .B1(_14160_),
    .Y(_14161_));
 sky130_fd_sc_hd__nand2_1 _35172_ (.A(_14161_),
    .B(net786),
    .Y(_14162_));
 sky130_fd_sc_hd__nand2_1 _35173_ (.A(net739),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[28] ),
    .Y(_14163_));
 sky130_fd_sc_hd__inv_1 _35174_ (.A(\inst$top.soc.cpu.sink__payload$18[137] ),
    .Y(_14164_));
 sky130_fd_sc_hd__nor2_1 _35175_ (.A(net2838),
    .B(_14164_),
    .Y(_14165_));
 sky130_fd_sc_hd__inv_1 _35176_ (.A(\inst$top.soc.cpu.shifter.m_result$7[28] ),
    .Y(_14166_));
 sky130_fd_sc_hd__o21ai_0 _35177_ (.A1(net2872),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[3] ),
    .B1(net2837),
    .Y(_14167_));
 sky130_fd_sc_hd__a21oi_1 _35178_ (.A1(net2872),
    .A2(_14166_),
    .B1(_14167_),
    .Y(_14168_));
 sky130_fd_sc_hd__o21ai_0 _35179_ (.A1(_14165_),
    .A2(_14168_),
    .B1(net2015),
    .Y(_14169_));
 sky130_fd_sc_hd__nand2_1 _35180_ (.A(net2923),
    .B(\inst$top.soc.cpu.divider.remainder[28] ),
    .Y(_14170_));
 sky130_fd_sc_hd__o21ai_0 _35181_ (.A1(net2922),
    .A2(_10224_),
    .B1(_14170_),
    .Y(_14171_));
 sky130_fd_sc_hd__nand2_1 _35182_ (.A(_14171_),
    .B(\inst$top.soc.cpu.d.sink__payload$6.divide ),
    .Y(_14172_));
 sky130_fd_sc_hd__a21oi_1 _35183_ (.A1(_14169_),
    .A2(_14172_),
    .B1(net2831),
    .Y(_14173_));
 sky130_fd_sc_hd__nand2_1 _35184_ (.A(_12984_),
    .B(_14173_),
    .Y(_14174_));
 sky130_fd_sc_hd__nand3_1 _35185_ (.A(_14162_),
    .B(_14163_),
    .C(_14174_),
    .Y(_14175_));
 sky130_fd_sc_hd__nand2_1 _35186_ (.A(net712),
    .B(_14175_),
    .Y(_14176_));
 sky130_fd_sc_hd__nand2_1 _35187_ (.A(net659),
    .B(\inst$top.soc.cpu.gprf.x_bypass1_data[28] ),
    .Y(_14177_));
 sky130_fd_sc_hd__a21oi_4 _35190_ (.A1(_14176_),
    .A2(_14177_),
    .B1(net3003),
    .Y(_04204_));
 sky130_fd_sc_hd__nand2_1 _35191_ (.A(net658),
    .B(_19921_),
    .Y(_14180_));
 sky130_fd_sc_hd__nand2_1 _35192_ (.A(_14180_),
    .B(net2181),
    .Y(_14181_));
 sky130_fd_sc_hd__inv_1 _35193_ (.A(_02933_),
    .Y(_14182_));
 sky130_fd_sc_hd__nor2_1 _35194_ (.A(_02938_),
    .B(_14077_),
    .Y(_14183_));
 sky130_fd_sc_hd__inv_1 _35195_ (.A(_14183_),
    .Y(_14184_));
 sky130_fd_sc_hd__nor2_1 _35196_ (.A(_14079_),
    .B(_14184_),
    .Y(_14185_));
 sky130_fd_sc_hd__nand3_1 _35197_ (.A(_13976_),
    .B(_13979_),
    .C(_14185_),
    .Y(_14186_));
 sky130_fd_sc_hd__inv_1 _35198_ (.A(_14185_),
    .Y(_14187_));
 sky130_fd_sc_hd__a21oi_1 _35199_ (.A1(_14136_),
    .A2(_02942_),
    .B1(_02940_),
    .Y(_14188_));
 sky130_fd_sc_hd__o21ai_0 _35200_ (.A1(_14187_),
    .A2(_13983_),
    .B1(_14188_),
    .Y(_14189_));
 sky130_fd_sc_hd__a21oi_1 _35201_ (.A1(_14086_),
    .A2(_14183_),
    .B1(_14189_),
    .Y(_14190_));
 sky130_fd_sc_hd__nand2_1 _35202_ (.A(_14186_),
    .B(_14190_),
    .Y(_14191_));
 sky130_fd_sc_hd__xor2_1 _35203_ (.A(_14182_),
    .B(_14191_),
    .X(_14192_));
 sky130_fd_sc_hd__nand2_1 _35204_ (.A(_14192_),
    .B(net2866),
    .Y(_14193_));
 sky130_fd_sc_hd__nand2_1 _35205_ (.A(_02938_),
    .B(_02918_),
    .Y(_14194_));
 sky130_fd_sc_hd__inv_1 _35206_ (.A(_14194_),
    .Y(_14195_));
 sky130_fd_sc_hd__nand2_1 _35207_ (.A(_14195_),
    .B(_14094_),
    .Y(_14196_));
 sky130_fd_sc_hd__nor2_1 _35208_ (.A(_14196_),
    .B(_13970_),
    .Y(_14197_));
 sky130_fd_sc_hd__nand4_1 _35209_ (.A(_13272_),
    .B(_13487_),
    .C(_13759_),
    .D(_14197_),
    .Y(_14198_));
 sky130_fd_sc_hd__nand2_1 _35210_ (.A(_13508_),
    .B(_13759_),
    .Y(_14199_));
 sky130_fd_sc_hd__nand2_1 _35211_ (.A(_13762_),
    .B(_14199_),
    .Y(_14200_));
 sky130_fd_sc_hd__a21oi_1 _35212_ (.A1(_02641_),
    .A2(_02938_),
    .B1(_02383_),
    .Y(_14201_));
 sky130_fd_sc_hd__inv_1 _35213_ (.A(_14201_),
    .Y(_14202_));
 sky130_fd_sc_hd__a21oi_1 _35214_ (.A1(_14099_),
    .A2(_14195_),
    .B1(_14202_),
    .Y(_14203_));
 sky130_fd_sc_hd__o21ai_0 _35215_ (.A1(_14196_),
    .A2(_13974_),
    .B1(_14203_),
    .Y(_14204_));
 sky130_fd_sc_hd__a21oi_1 _35216_ (.A1(_14200_),
    .A2(_14197_),
    .B1(_14204_),
    .Y(_14205_));
 sky130_fd_sc_hd__nand2_1 _35217_ (.A(_14198_),
    .B(_14205_),
    .Y(_14206_));
 sky130_fd_sc_hd__nand2_1 _35218_ (.A(_14206_),
    .B(_14182_),
    .Y(_14207_));
 sky130_fd_sc_hd__nand3_1 _35219_ (.A(_14198_),
    .B(_14205_),
    .C(_02933_),
    .Y(_14208_));
 sky130_fd_sc_hd__nand2_1 _35220_ (.A(_14207_),
    .B(_14208_),
    .Y(_14209_));
 sky130_fd_sc_hd__nand2_1 _35221_ (.A(_14209_),
    .B(net2005),
    .Y(_14210_));
 sky130_fd_sc_hd__nand2_1 _35222_ (.A(_14193_),
    .B(_14210_),
    .Y(_14211_));
 sky130_fd_sc_hd__nand2_1 _35223_ (.A(_14211_),
    .B(net2215),
    .Y(_14212_));
 sky130_fd_sc_hd__nand2_1 _35224_ (.A(_14212_),
    .B(_05859_),
    .Y(_14213_));
 sky130_fd_sc_hd__nand2_1 _35225_ (.A(_14213_),
    .B(net2020),
    .Y(_14214_));
 sky130_fd_sc_hd__nand2_1 _35226_ (.A(net1796),
    .B(_03292_),
    .Y(_14215_));
 sky130_fd_sc_hd__nand2_1 _35227_ (.A(net1868),
    .B(_03291_),
    .Y(_14216_));
 sky130_fd_sc_hd__o211ai_1 _35228_ (.A1(_03295_),
    .A2(net1230),
    .B1(_14215_),
    .C1(_14216_),
    .Y(_14217_));
 sky130_fd_sc_hd__a21oi_1 _35229_ (.A1(_14217_),
    .A2(net2862),
    .B1(net2854),
    .Y(_14218_));
 sky130_fd_sc_hd__nand2_1 _35230_ (.A(\inst$top.soc.cpu.sink__payload$12[28] ),
    .B(\inst$top.soc.cpu.sink__payload$12[27] ),
    .Y(_14219_));
 sky130_fd_sc_hd__or4_1 _35231_ (.A(_13790_),
    .B(_13862_),
    .C(_14114_),
    .D(_14219_),
    .X(_14220_));
 sky130_fd_sc_hd__nor4_1 _35232_ (.A(_13862_),
    .B(_14114_),
    .C(_14219_),
    .D(_13790_),
    .Y(_14221_));
 sky130_fd_sc_hd__nand2_1 _35233_ (.A(_14221_),
    .B(_19920_),
    .Y(_14222_));
 sky130_fd_sc_hd__nand2_1 _35234_ (.A(_14222_),
    .B(net2854),
    .Y(_14223_));
 sky130_fd_sc_hd__a21oi_1 _35235_ (.A1(\inst$top.soc.cpu.sink__payload$12[29] ),
    .A2(_14220_),
    .B1(_14223_),
    .Y(_14224_));
 sky130_fd_sc_hd__a21oi_2 _35236_ (.A1(_14214_),
    .A2(_14218_),
    .B1(_14224_),
    .Y(_14225_));
 sky130_fd_sc_hd__nand2_1 _35237_ (.A(_14225_),
    .B(net786),
    .Y(_14226_));
 sky130_fd_sc_hd__nand2_1 _35238_ (.A(net739),
    .B(net915),
    .Y(_14227_));
 sky130_fd_sc_hd__inv_1 _35239_ (.A(\inst$top.soc.cpu.sink__payload$18[138] ),
    .Y(_14228_));
 sky130_fd_sc_hd__nor2_1 _35240_ (.A(net2833),
    .B(_14228_),
    .Y(_14229_));
 sky130_fd_sc_hd__inv_1 _35241_ (.A(\inst$top.soc.cpu.shifter.m_result$7[29] ),
    .Y(_14230_));
 sky130_fd_sc_hd__o21ai_0 _35242_ (.A1(net2869),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[2] ),
    .B1(net2835),
    .Y(_14231_));
 sky130_fd_sc_hd__a21oi_1 _35243_ (.A1(net2870),
    .A2(_14230_),
    .B1(_14231_),
    .Y(_14232_));
 sky130_fd_sc_hd__o21ai_0 _35244_ (.A1(_14229_),
    .A2(_14232_),
    .B1(net2014),
    .Y(_14233_));
 sky130_fd_sc_hd__a21oi_1 _35245_ (.A1(_10745_),
    .A2(net2923),
    .B1(net2011),
    .Y(_14234_));
 sky130_fd_sc_hd__o21ai_1 _35246_ (.A1(net2921),
    .A2(\inst$top.soc.cpu.divider.quotient[29] ),
    .B1(_14234_),
    .Y(_14235_));
 sky130_fd_sc_hd__a21oi_1 _35247_ (.A1(_14233_),
    .A2(net1783),
    .B1(net2830),
    .Y(_14236_));
 sky130_fd_sc_hd__nand2_1 _35248_ (.A(_12984_),
    .B(_14236_),
    .Y(_14237_));
 sky130_fd_sc_hd__nand3_1 _35249_ (.A(_14226_),
    .B(_14227_),
    .C(_14237_),
    .Y(_14238_));
 sky130_fd_sc_hd__nor2_1 _35250_ (.A(net658),
    .B(_14238_),
    .Y(_14239_));
 sky130_fd_sc_hd__nor2_4 _35251_ (.A(_14181_),
    .B(_14239_),
    .Y(_04205_));
 sky130_fd_sc_hd__nor2_1 _35252_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[2] ),
    .B(net701),
    .Y(_14240_));
 sky130_fd_sc_hd__inv_1 _35253_ (.A(\inst$top.soc.cpu.sink__payload$18[111] ),
    .Y(_14241_));
 sky130_fd_sc_hd__nor2_1 _35254_ (.A(net2833),
    .B(_14241_),
    .Y(_14242_));
 sky130_fd_sc_hd__o21ai_0 _35255_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[2] ),
    .A2(net2002),
    .B1(net2835),
    .Y(_14243_));
 sky130_fd_sc_hd__a21oi_1 _35256_ (.A1(net2002),
    .A2(_14230_),
    .B1(_14243_),
    .Y(_14244_));
 sky130_fd_sc_hd__o21ai_0 _35257_ (.A1(_14242_),
    .A2(_14244_),
    .B1(net2016),
    .Y(_14245_));
 sky130_fd_sc_hd__a21oi_1 _35258_ (.A1(_10328_),
    .A2(net2924),
    .B1(net2011),
    .Y(_14246_));
 sky130_fd_sc_hd__o21ai_1 _35259_ (.A1(net2921),
    .A2(\inst$top.soc.cpu.divider.quotient[2] ),
    .B1(_14246_),
    .Y(_14247_));
 sky130_fd_sc_hd__a21oi_1 _35260_ (.A1(_14245_),
    .A2(net1782),
    .B1(net2832),
    .Y(_14248_));
 sky130_fd_sc_hd__inv_1 _35261_ (.A(_14248_),
    .Y(_14249_));
 sky130_fd_sc_hd__nand2_1 _35262_ (.A(net2865),
    .B(_00170_),
    .Y(_14250_));
 sky130_fd_sc_hd__o21ai_0 _35263_ (.A1(net2865),
    .A2(_00165_),
    .B1(_14250_),
    .Y(_14251_));
 sky130_fd_sc_hd__xor2_2 _35264_ (.A(_13071_),
    .B(_14251_),
    .X(_14252_));
 sky130_fd_sc_hd__nand2_1 _35265_ (.A(net869),
    .B(net2214),
    .Y(_14253_));
 sky130_fd_sc_hd__nand2_1 _35266_ (.A(_20483_),
    .B(_14253_),
    .Y(_14254_));
 sky130_fd_sc_hd__nand2_1 _35267_ (.A(_14254_),
    .B(net2018),
    .Y(_14255_));
 sky130_fd_sc_hd__nand2_1 _35268_ (.A(net1797),
    .B(_03101_),
    .Y(_14256_));
 sky130_fd_sc_hd__nand2_1 _35269_ (.A(net1870),
    .B(_03100_),
    .Y(_14257_));
 sky130_fd_sc_hd__o211ai_1 _35270_ (.A1(_03104_),
    .A2(net1231),
    .B1(_14256_),
    .C1(_14257_),
    .Y(_14258_));
 sky130_fd_sc_hd__a21oi_1 _35271_ (.A1(_14258_),
    .A2(net2861),
    .B1(net2852),
    .Y(_14259_));
 sky130_fd_sc_hd__a22oi_1 _35272_ (.A1(\inst$top.soc.cpu.sink__payload$12[2] ),
    .A2(net2852),
    .B1(_14255_),
    .B2(_14259_),
    .Y(_14260_));
 sky130_fd_sc_hd__inv_1 _35273_ (.A(_14260_),
    .Y(_14261_));
 sky130_fd_sc_hd__o22ai_1 _35274_ (.A1(_14249_),
    .A2(net783),
    .B1(_14261_),
    .B2(net736),
    .Y(_14262_));
 sky130_fd_sc_hd__a21oi_1 _35275_ (.A1(net737),
    .A2(net1063),
    .B1(_14262_),
    .Y(_14263_));
 sky130_fd_sc_hd__nand2_1 _35276_ (.A(net701),
    .B(_14263_),
    .Y(_14264_));
 sky130_fd_sc_hd__nand2_1 _35277_ (.A(_14264_),
    .B(net2154),
    .Y(_14265_));
 sky130_fd_sc_hd__nor2_2 _35278_ (.A(_14240_),
    .B(_14265_),
    .Y(_04206_));
 sky130_fd_sc_hd__nand2_1 _35279_ (.A(net657),
    .B(_19905_),
    .Y(_14266_));
 sky130_fd_sc_hd__nand2_1 _35280_ (.A(_14266_),
    .B(net2156),
    .Y(_14267_));
 sky130_fd_sc_hd__inv_1 _35281_ (.A(\inst$top.soc.cpu.sink__payload$18[139] ),
    .Y(_14268_));
 sky130_fd_sc_hd__nor2_1 _35282_ (.A(net2834),
    .B(_14268_),
    .Y(_14269_));
 sky130_fd_sc_hd__inv_1 _35283_ (.A(\inst$top.soc.cpu.shifter.m_result$7[30] ),
    .Y(_14270_));
 sky130_fd_sc_hd__o21ai_0 _35284_ (.A1(net2869),
    .A2(\inst$top.soc.cpu.shifter.m_result$7[1] ),
    .B1(net2835),
    .Y(_14271_));
 sky130_fd_sc_hd__a21oi_1 _35285_ (.A1(net2869),
    .A2(_14270_),
    .B1(_14271_),
    .Y(_14272_));
 sky130_fd_sc_hd__o21ai_0 _35286_ (.A1(_14269_),
    .A2(_14272_),
    .B1(net2013),
    .Y(_14273_));
 sky130_fd_sc_hd__a21oi_1 _35287_ (.A1(_10772_),
    .A2(net2923),
    .B1(net2012),
    .Y(_14274_));
 sky130_fd_sc_hd__o21ai_2 _35288_ (.A1(net2922),
    .A2(\inst$top.soc.cpu.divider.quotient[30] ),
    .B1(_14274_),
    .Y(_14275_));
 sky130_fd_sc_hd__nand2_1 _35289_ (.A(_14273_),
    .B(_14275_),
    .Y(_14276_));
 sky130_fd_sc_hd__nand2_1 _35290_ (.A(_14276_),
    .B(_12997_),
    .Y(_14277_));
 sky130_fd_sc_hd__nor2_1 _35291_ (.A(_14277_),
    .B(net783),
    .Y(_14278_));
 sky130_fd_sc_hd__a21oi_1 _35292_ (.A1(net737),
    .A2(net910),
    .B1(_14278_),
    .Y(_14279_));
 sky130_fd_sc_hd__nand3_1 _35293_ (.A(net665),
    .B(net755),
    .C(_14279_),
    .Y(_14280_));
 sky130_fd_sc_hd__nand2_1 _35294_ (.A(_02933_),
    .B(_02938_),
    .Y(_14281_));
 sky130_fd_sc_hd__nor2_1 _35295_ (.A(_14281_),
    .B(_14123_),
    .Y(_14282_));
 sky130_fd_sc_hd__nand4_1 _35296_ (.A(_13308_),
    .B(_13830_),
    .C(_14037_),
    .D(_14282_),
    .Y(_14283_));
 sky130_fd_sc_hd__nand3_1 _35297_ (.A(_14126_),
    .B(_02933_),
    .C(_02938_),
    .Y(_14284_));
 sky130_fd_sc_hd__a21oi_1 _35298_ (.A1(_02383_),
    .A2(_02933_),
    .B1(_02438_),
    .Y(_14285_));
 sky130_fd_sc_hd__nand2_1 _35299_ (.A(_14284_),
    .B(_14285_),
    .Y(_14286_));
 sky130_fd_sc_hd__nand2_1 _35300_ (.A(_14282_),
    .B(_14037_),
    .Y(_14287_));
 sky130_fd_sc_hd__nor2_1 _35301_ (.A(_14287_),
    .B(_13835_),
    .Y(_14288_));
 sky130_fd_sc_hd__a211oi_1 _35302_ (.A1(_14040_),
    .A2(_14282_),
    .B1(_14286_),
    .C1(_14288_),
    .Y(_14289_));
 sky130_fd_sc_hd__nand2_1 _35303_ (.A(_14283_),
    .B(_14289_),
    .Y(_14290_));
 sky130_fd_sc_hd__xor2_1 _35304_ (.A(_02928_),
    .B(_14290_),
    .X(_14291_));
 sky130_fd_sc_hd__nand2_1 _35305_ (.A(_14291_),
    .B(net2005),
    .Y(_14292_));
 sky130_fd_sc_hd__nand2_1 _35306_ (.A(_14182_),
    .B(_14136_),
    .Y(_14293_));
 sky130_fd_sc_hd__nor2_1 _35307_ (.A(_14137_),
    .B(_14293_),
    .Y(_14294_));
 sky130_fd_sc_hd__a21oi_1 _35308_ (.A1(_14182_),
    .A2(_02940_),
    .B1(_02935_),
    .Y(_14295_));
 sky130_fd_sc_hd__o21ai_0 _35309_ (.A1(_14293_),
    .A2(_14141_),
    .B1(_14295_),
    .Y(_14296_));
 sky130_fd_sc_hd__a21oi_1 _35310_ (.A1(_14033_),
    .A2(_14294_),
    .B1(_14296_),
    .Y(_14297_));
 sky130_fd_sc_hd__xor2_1 _35311_ (.A(_02928_),
    .B(_14297_),
    .X(_14298_));
 sky130_fd_sc_hd__nand2_1 _35312_ (.A(_14298_),
    .B(net2866),
    .Y(_14299_));
 sky130_fd_sc_hd__nand2_1 _35313_ (.A(_14292_),
    .B(_14299_),
    .Y(_14300_));
 sky130_fd_sc_hd__nand2_1 _35314_ (.A(_14300_),
    .B(net2215),
    .Y(_14301_));
 sky130_fd_sc_hd__nand2_1 _35315_ (.A(_14301_),
    .B(_05874_),
    .Y(_14302_));
 sky130_fd_sc_hd__nand2_1 _35316_ (.A(_14302_),
    .B(net2017),
    .Y(_14303_));
 sky130_fd_sc_hd__nand2_1 _35317_ (.A(net1795),
    .B(_03299_),
    .Y(_14304_));
 sky130_fd_sc_hd__nand2_1 _35318_ (.A(net1868),
    .B(_03298_),
    .Y(_14305_));
 sky130_fd_sc_hd__o211ai_1 _35319_ (.A1(_03302_),
    .A2(net1229),
    .B1(_14304_),
    .C1(_14305_),
    .Y(_14306_));
 sky130_fd_sc_hd__a21oi_1 _35320_ (.A1(_14306_),
    .A2(net2862),
    .B1(net2856),
    .Y(_14307_));
 sky130_fd_sc_hd__nand2_1 _35321_ (.A(_14303_),
    .B(_14307_),
    .Y(_14308_));
 sky130_fd_sc_hd__nor4_1 _35322_ (.A(_19920_),
    .B(_12420_),
    .C(_14219_),
    .D(_14053_),
    .Y(_14309_));
 sky130_fd_sc_hd__or2_2 _35323_ (.A(_19900_),
    .B(_14309_),
    .X(_14310_));
 sky130_fd_sc_hd__nand2_1 _35324_ (.A(_14309_),
    .B(_19900_),
    .Y(_14311_));
 sky130_fd_sc_hd__nand3_1 _35325_ (.A(_14310_),
    .B(net2853),
    .C(_14311_),
    .Y(_14312_));
 sky130_fd_sc_hd__nand2_1 _35326_ (.A(_14308_),
    .B(_14312_),
    .Y(_14313_));
 sky130_fd_sc_hd__nor2_1 _35327_ (.A(net736),
    .B(_14313_),
    .Y(_14314_));
 sky130_fd_sc_hd__nor2_1 _35328_ (.A(_14280_),
    .B(_14314_),
    .Y(_14315_));
 sky130_fd_sc_hd__nor2_4 _35329_ (.A(_14267_),
    .B(_14315_),
    .Y(_04207_));
 sky130_fd_sc_hd__nand4_1 _35330_ (.A(\inst$top.soc.cpu.sink__payload$12[30] ),
    .B(\inst$top.soc.cpu.sink__payload$12[29] ),
    .C(\inst$top.soc.cpu.sink__payload$12[28] ),
    .D(\inst$top.soc.cpu.sink__payload$12[27] ),
    .Y(_14316_));
 sky130_fd_sc_hd__nor4_1 _35331_ (.A(\inst$top.soc.cpu.sink__payload$12[31] ),
    .B(_14114_),
    .C(_14316_),
    .D(_13864_),
    .Y(_14317_));
 sky130_fd_sc_hd__nor3_1 _35332_ (.A(_14114_),
    .B(_14316_),
    .C(_13864_),
    .Y(_14318_));
 sky130_fd_sc_hd__o21ai_0 _35333_ (.A1(_19869_),
    .A2(_14318_),
    .B1(net2851),
    .Y(_14319_));
 sky130_fd_sc_hd__nand2_1 _35334_ (.A(_05889_),
    .B(net2017),
    .Y(_14320_));
 sky130_fd_sc_hd__nor3_1 _35335_ (.A(_02928_),
    .B(_02933_),
    .C(_14184_),
    .Y(_14321_));
 sky130_fd_sc_hd__inv_1 _35336_ (.A(_14321_),
    .Y(_14322_));
 sky130_fd_sc_hd__nand2_1 _35337_ (.A(_14321_),
    .B(_14080_),
    .Y(_14323_));
 sky130_fd_sc_hd__a21boi_0 _35338_ (.A1(_13641_),
    .A2(_13877_),
    .B1_N(_13883_),
    .Y(_14324_));
 sky130_fd_sc_hd__o21bai_1 _35339_ (.A1(_02933_),
    .A2(_14188_),
    .B1_N(_02935_),
    .Y(_14325_));
 sky130_fd_sc_hd__inv_1 _35340_ (.A(_02928_),
    .Y(_14326_));
 sky130_fd_sc_hd__a21oi_1 _35341_ (.A1(_14325_),
    .A2(_14326_),
    .B1(_02930_),
    .Y(_14327_));
 sky130_fd_sc_hd__o221a_2 _35342_ (.A1(_14087_),
    .A2(_14322_),
    .B1(_14323_),
    .B2(_14324_),
    .C1(_14327_),
    .X(_14328_));
 sky130_fd_sc_hd__nor3_1 _35343_ (.A(_13635_),
    .B(_14078_),
    .C(_14323_),
    .Y(_14329_));
 sky130_fd_sc_hd__nand2_1 _35344_ (.A(_13362_),
    .B(_14329_),
    .Y(_14330_));
 sky130_fd_sc_hd__nand2_1 _35345_ (.A(_14328_),
    .B(_14330_),
    .Y(_14331_));
 sky130_fd_sc_hd__nand2_1 _35346_ (.A(_14331_),
    .B(_02922_),
    .Y(_14332_));
 sky130_fd_sc_hd__nand3_1 _35347_ (.A(_14328_),
    .B(_09916_),
    .C(_14330_),
    .Y(_14333_));
 sky130_fd_sc_hd__nand3_1 _35348_ (.A(_14332_),
    .B(_14333_),
    .C(net2866),
    .Y(_14334_));
 sky130_fd_sc_hd__nor3_1 _35349_ (.A(_14326_),
    .B(_14182_),
    .C(_14194_),
    .Y(_14335_));
 sky130_fd_sc_hd__nand2_1 _35350_ (.A(_14103_),
    .B(_14335_),
    .Y(_14336_));
 sky130_fd_sc_hd__nand3_1 _35351_ (.A(_14202_),
    .B(_02928_),
    .C(_02933_),
    .Y(_14337_));
 sky130_fd_sc_hd__a21oi_1 _35352_ (.A1(_02438_),
    .A2(_02928_),
    .B1(_02678_),
    .Y(_14338_));
 sky130_fd_sc_hd__nand3_1 _35353_ (.A(_14336_),
    .B(_14337_),
    .C(_14338_),
    .Y(_14339_));
 sky130_fd_sc_hd__xor2_1 _35354_ (.A(_09916_),
    .B(_14339_),
    .X(_14340_));
 sky130_fd_sc_hd__nand2_1 _35355_ (.A(_14340_),
    .B(net2005),
    .Y(_14341_));
 sky130_fd_sc_hd__nand2_1 _35356_ (.A(_14334_),
    .B(_14341_),
    .Y(_14342_));
 sky130_fd_sc_hd__nor2_1 _35357_ (.A(net2843),
    .B(_14342_),
    .Y(_14343_));
 sky130_fd_sc_hd__nand2_1 _35358_ (.A(net1795),
    .B(_03306_),
    .Y(_14344_));
 sky130_fd_sc_hd__nand2_1 _35359_ (.A(net1868),
    .B(_03305_),
    .Y(_14345_));
 sky130_fd_sc_hd__o211ai_1 _35360_ (.A1(_03309_),
    .A2(net1229),
    .B1(_14344_),
    .C1(_14345_),
    .Y(_14346_));
 sky130_fd_sc_hd__a21oi_1 _35361_ (.A1(_14346_),
    .A2(net2862),
    .B1(net2856),
    .Y(_14347_));
 sky130_fd_sc_hd__o21ai_0 _35362_ (.A1(_14320_),
    .A2(_14343_),
    .B1(_14347_),
    .Y(_14348_));
 sky130_fd_sc_hd__o21ai_1 _35363_ (.A1(_14317_),
    .A2(_14319_),
    .B1(_14348_),
    .Y(_14349_));
 sky130_fd_sc_hd__nor2_1 _35364_ (.A(net736),
    .B(_14349_),
    .Y(_14350_));
 sky130_fd_sc_hd__inv_1 _35365_ (.A(\inst$top.soc.cpu.sink__payload$18[140] ),
    .Y(_14351_));
 sky130_fd_sc_hd__nor2_1 _35366_ (.A(net2834),
    .B(_14351_),
    .Y(_14352_));
 sky130_fd_sc_hd__o21ai_0 _35367_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[0] ),
    .A2(net2871),
    .B1(net2840),
    .Y(_14353_));
 sky130_fd_sc_hd__a21oi_1 _35368_ (.A1(_12990_),
    .A2(net2871),
    .B1(_14353_),
    .Y(_14354_));
 sky130_fd_sc_hd__o21ai_0 _35369_ (.A1(_14352_),
    .A2(_14354_),
    .B1(net2013),
    .Y(_14355_));
 sky130_fd_sc_hd__a21oi_1 _35370_ (.A1(_09930_),
    .A2(net2922),
    .B1(net2012),
    .Y(_14356_));
 sky130_fd_sc_hd__o21ai_1 _35371_ (.A1(net2923),
    .A2(\inst$top.soc.cpu.divider.quotient[31] ),
    .B1(_14356_),
    .Y(_14357_));
 sky130_fd_sc_hd__nand2_1 _35372_ (.A(_14355_),
    .B(net1781),
    .Y(_14358_));
 sky130_fd_sc_hd__nand2_1 _35373_ (.A(_14358_),
    .B(_12997_),
    .Y(_14359_));
 sky130_fd_sc_hd__nor2_1 _35374_ (.A(_14359_),
    .B(net783),
    .Y(_14360_));
 sky130_fd_sc_hd__a21oi_1 _35375_ (.A1(net737),
    .A2(net905),
    .B1(_14360_),
    .Y(_14361_));
 sky130_fd_sc_hd__nand3_1 _35376_ (.A(net665),
    .B(net755),
    .C(_14361_),
    .Y(_14362_));
 sky130_fd_sc_hd__nor2_1 _35377_ (.A(_14350_),
    .B(_14362_),
    .Y(_14363_));
 sky130_fd_sc_hd__nand2_1 _35378_ (.A(net654),
    .B(_19875_),
    .Y(_14364_));
 sky130_fd_sc_hd__nand2_1 _35379_ (.A(_14364_),
    .B(net2154),
    .Y(_14365_));
 sky130_fd_sc_hd__nor2_2 _35380_ (.A(_14363_),
    .B(_14365_),
    .Y(_04208_));
 sky130_fd_sc_hd__nor2_1 _35382_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[3] ),
    .B(net701),
    .Y(_14367_));
 sky130_fd_sc_hd__nand2_1 _35383_ (.A(_13156_),
    .B(net2005),
    .Y(_14368_));
 sky130_fd_sc_hd__o21ai_0 _35384_ (.A1(net2005),
    .A2(_13257_),
    .B1(_14368_),
    .Y(_14369_));
 sky130_fd_sc_hd__xor2_2 _35385_ (.A(_13061_),
    .B(_14369_),
    .X(_14370_));
 sky130_fd_sc_hd__nand2_1 _35386_ (.A(net830),
    .B(net2214),
    .Y(_14371_));
 sky130_fd_sc_hd__nand3_1 _35387_ (.A(_20524_),
    .B(_14371_),
    .C(net2018),
    .Y(_14372_));
 sky130_fd_sc_hd__nor2_1 _35388_ (.A(_03111_),
    .B(net1231),
    .Y(_14373_));
 sky130_fd_sc_hd__a221oi_1 _35389_ (.A1(net1797),
    .A2(_03108_),
    .B1(net1870),
    .B2(_03107_),
    .C1(_14373_),
    .Y(_14374_));
 sky130_fd_sc_hd__a21oi_1 _35390_ (.A1(_14374_),
    .A2(net2861),
    .B1(net2852),
    .Y(_14375_));
 sky130_fd_sc_hd__a22o_1 _35391_ (.A1(net2852),
    .A2(_03113_),
    .B1(_14372_),
    .B2(_14375_),
    .X(_14376_));
 sky130_fd_sc_hd__inv_1 _35392_ (.A(\inst$top.soc.cpu.sink__payload$18[112] ),
    .Y(_14377_));
 sky130_fd_sc_hd__nor2_1 _35393_ (.A(net2833),
    .B(_14377_),
    .Y(_14378_));
 sky130_fd_sc_hd__o21ai_0 _35394_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[3] ),
    .A2(net2003),
    .B1(net2837),
    .Y(_14379_));
 sky130_fd_sc_hd__a21oi_1 _35395_ (.A1(net2004),
    .A2(_14166_),
    .B1(_14379_),
    .Y(_14380_));
 sky130_fd_sc_hd__o21ai_0 _35396_ (.A1(_14378_),
    .A2(_14380_),
    .B1(net2013),
    .Y(_14381_));
 sky130_fd_sc_hd__a21oi_1 _35397_ (.A1(_10329_),
    .A2(net2924),
    .B1(net2011),
    .Y(_14382_));
 sky130_fd_sc_hd__o21ai_1 _35398_ (.A1(net2921),
    .A2(\inst$top.soc.cpu.divider.quotient[3] ),
    .B1(_14382_),
    .Y(_14383_));
 sky130_fd_sc_hd__a21oi_1 _35399_ (.A1(_14381_),
    .A2(net1780),
    .B1(net2829),
    .Y(_14384_));
 sky130_fd_sc_hd__inv_1 _35400_ (.A(_14384_),
    .Y(_14385_));
 sky130_fd_sc_hd__o22ai_1 _35401_ (.A1(_14385_),
    .A2(net784),
    .B1(_20537_),
    .B2(_12956_),
    .Y(_14386_));
 sky130_fd_sc_hd__a21oi_1 _35402_ (.A1(net787),
    .A2(_14376_),
    .B1(_14386_),
    .Y(_14387_));
 sky130_fd_sc_hd__nand2_1 _35403_ (.A(net701),
    .B(_14387_),
    .Y(_14388_));
 sky130_fd_sc_hd__nand2_1 _35404_ (.A(_14388_),
    .B(net2154),
    .Y(_14389_));
 sky130_fd_sc_hd__nor2_2 _35405_ (.A(_14367_),
    .B(_14389_),
    .Y(_04209_));
 sky130_fd_sc_hd__nor2_1 _35406_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[4] ),
    .B(net701),
    .Y(_14390_));
 sky130_fd_sc_hd__inv_1 _35407_ (.A(\inst$top.soc.cpu.sink__payload$18[113] ),
    .Y(_14391_));
 sky130_fd_sc_hd__nor2_1 _35408_ (.A(net2833),
    .B(_14391_),
    .Y(_14392_));
 sky130_fd_sc_hd__o21ai_0 _35409_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[4] ),
    .A2(net2002),
    .B1(net2835),
    .Y(_14393_));
 sky130_fd_sc_hd__a21oi_1 _35410_ (.A1(net2002),
    .A2(_14068_),
    .B1(_14393_),
    .Y(_14394_));
 sky130_fd_sc_hd__o21ai_0 _35411_ (.A1(_14392_),
    .A2(_14394_),
    .B1(net2013),
    .Y(_14395_));
 sky130_fd_sc_hd__a21oi_1 _35412_ (.A1(_10369_),
    .A2(net2920),
    .B1(net2011),
    .Y(_14396_));
 sky130_fd_sc_hd__o21ai_1 _35413_ (.A1(net2919),
    .A2(\inst$top.soc.cpu.divider.quotient[4] ),
    .B1(_14396_),
    .Y(_14397_));
 sky130_fd_sc_hd__a21oi_1 _35414_ (.A1(_14395_),
    .A2(net1779),
    .B1(net2832),
    .Y(_14398_));
 sky130_fd_sc_hd__inv_1 _35415_ (.A(_14398_),
    .Y(_14399_));
 sky130_fd_sc_hd__nand2_1 _35416_ (.A(_13047_),
    .B(net2865),
    .Y(_14400_));
 sky130_fd_sc_hd__o21ai_0 _35417_ (.A1(net2865),
    .A2(_13414_),
    .B1(_14400_),
    .Y(_14401_));
 sky130_fd_sc_hd__xor2_2 _35418_ (.A(_03065_),
    .B(_14401_),
    .X(_14402_));
 sky130_fd_sc_hd__nand2_1 _35419_ (.A(net812),
    .B(net2214),
    .Y(_14403_));
 sky130_fd_sc_hd__nand2_1 _35420_ (.A(_20554_),
    .B(_14403_),
    .Y(_14404_));
 sky130_fd_sc_hd__nand2_1 _35421_ (.A(_14404_),
    .B(net2018),
    .Y(_14405_));
 sky130_fd_sc_hd__nand2_1 _35422_ (.A(net1797),
    .B(_03117_),
    .Y(_14406_));
 sky130_fd_sc_hd__nand2_1 _35423_ (.A(net1870),
    .B(_03116_),
    .Y(_14407_));
 sky130_fd_sc_hd__o211ai_1 _35424_ (.A1(_03120_),
    .A2(net1231),
    .B1(_14406_),
    .C1(_14407_),
    .Y(_14408_));
 sky130_fd_sc_hd__a21oi_1 _35425_ (.A1(_14408_),
    .A2(net2861),
    .B1(net2853),
    .Y(_14409_));
 sky130_fd_sc_hd__or2_2 _35426_ (.A(\inst$top.soc.cpu.sink__payload$12[4] ),
    .B(_03112_),
    .X(_14410_));
 sky130_fd_sc_hd__a21oi_1 _35427_ (.A1(_14410_),
    .A2(_13031_),
    .B1(_13129_),
    .Y(_14411_));
 sky130_fd_sc_hd__a21oi_1 _35428_ (.A1(_14405_),
    .A2(_14409_),
    .B1(_14411_),
    .Y(_14412_));
 sky130_fd_sc_hd__inv_1 _35429_ (.A(_14412_),
    .Y(_14413_));
 sky130_fd_sc_hd__o22ai_1 _35430_ (.A1(_14399_),
    .A2(net783),
    .B1(_14413_),
    .B2(net736),
    .Y(_14414_));
 sky130_fd_sc_hd__a21oi_1 _35431_ (.A1(net737),
    .A2(net1013),
    .B1(_14414_),
    .Y(_14415_));
 sky130_fd_sc_hd__nand2_1 _35432_ (.A(net701),
    .B(_14415_),
    .Y(_14416_));
 sky130_fd_sc_hd__nand2_1 _35433_ (.A(_14416_),
    .B(net2151),
    .Y(_14417_));
 sky130_fd_sc_hd__nor2_2 _35434_ (.A(_14390_),
    .B(_14417_),
    .Y(_04210_));
 sky130_fd_sc_hd__nor2_1 _35435_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[5] ),
    .B(net704),
    .Y(_14418_));
 sky130_fd_sc_hd__inv_1 _35436_ (.A(\inst$top.soc.cpu.sink__payload$18[114] ),
    .Y(_14419_));
 sky130_fd_sc_hd__nor2_1 _35437_ (.A(net2835),
    .B(_14419_),
    .Y(_14420_));
 sky130_fd_sc_hd__o21ai_0 _35438_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[5] ),
    .A2(net2002),
    .B1(net2835),
    .Y(_14421_));
 sky130_fd_sc_hd__a21oi_1 _35439_ (.A1(net2002),
    .A2(_14014_),
    .B1(_14421_),
    .Y(_14422_));
 sky130_fd_sc_hd__o21ai_0 _35440_ (.A1(_14420_),
    .A2(_14422_),
    .B1(net2014),
    .Y(_14423_));
 sky130_fd_sc_hd__a21oi_1 _35441_ (.A1(_10832_),
    .A2(net2920),
    .B1(net2010),
    .Y(_14424_));
 sky130_fd_sc_hd__o21ai_2 _35442_ (.A1(net2919),
    .A2(\inst$top.soc.cpu.divider.quotient[5] ),
    .B1(_14424_),
    .Y(_14425_));
 sky130_fd_sc_hd__a21oi_1 _35443_ (.A1(_14423_),
    .A2(_14425_),
    .B1(net2830),
    .Y(_14426_));
 sky130_fd_sc_hd__inv_1 _35444_ (.A(_14426_),
    .Y(_14427_));
 sky130_fd_sc_hd__nand2_1 _35445_ (.A(_13259_),
    .B(net2865),
    .Y(_14428_));
 sky130_fd_sc_hd__nor2_1 _35446_ (.A(_00162_),
    .B(_13490_),
    .Y(_14429_));
 sky130_fd_sc_hd__nor2_1 _35447_ (.A(_14429_),
    .B(_13495_),
    .Y(_14430_));
 sky130_fd_sc_hd__nand2_1 _35448_ (.A(_14430_),
    .B(net2005),
    .Y(_14431_));
 sky130_fd_sc_hd__nand2_1 _35449_ (.A(_14428_),
    .B(_14431_),
    .Y(_14432_));
 sky130_fd_sc_hd__xor2_1 _35450_ (.A(_03060_),
    .B(_14432_),
    .X(_14433_));
 sky130_fd_sc_hd__inv_1 _35451_ (.A(_14433_),
    .Y(_14434_));
 sky130_fd_sc_hd__o21ai_0 _35452_ (.A1(net2847),
    .A2(_14434_),
    .B1(_20581_),
    .Y(_14435_));
 sky130_fd_sc_hd__nand2_1 _35453_ (.A(_14435_),
    .B(net2018),
    .Y(_14436_));
 sky130_fd_sc_hd__nand2_1 _35454_ (.A(net1797),
    .B(_03124_),
    .Y(_14437_));
 sky130_fd_sc_hd__nand2_1 _35455_ (.A(net1870),
    .B(_03123_),
    .Y(_14438_));
 sky130_fd_sc_hd__o211ai_1 _35456_ (.A1(_03127_),
    .A2(net1231),
    .B1(_14437_),
    .C1(_14438_),
    .Y(_14439_));
 sky130_fd_sc_hd__a21oi_1 _35457_ (.A1(_14439_),
    .A2(net2861),
    .B1(net2852),
    .Y(_14440_));
 sky130_fd_sc_hd__xor2_1 _35458_ (.A(_20566_),
    .B(_13116_),
    .X(_14441_));
 sky130_fd_sc_hd__nor2_1 _35459_ (.A(net2001),
    .B(_14441_),
    .Y(_14442_));
 sky130_fd_sc_hd__a21oi_1 _35460_ (.A1(_14436_),
    .A2(_14440_),
    .B1(_14442_),
    .Y(_14443_));
 sky130_fd_sc_hd__inv_1 _35461_ (.A(_14443_),
    .Y(_14444_));
 sky130_fd_sc_hd__o22ai_1 _35462_ (.A1(_14427_),
    .A2(net784),
    .B1(_14444_),
    .B2(net736),
    .Y(_14445_));
 sky130_fd_sc_hd__a21oi_1 _35463_ (.A1(net737),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[5] ),
    .B1(_14445_),
    .Y(_14446_));
 sky130_fd_sc_hd__nand2_1 _35464_ (.A(net704),
    .B(_14446_),
    .Y(_14447_));
 sky130_fd_sc_hd__nand2_1 _35465_ (.A(_14447_),
    .B(net2152),
    .Y(_14448_));
 sky130_fd_sc_hd__nor2_2 _35466_ (.A(_14418_),
    .B(_14448_),
    .Y(_04211_));
 sky130_fd_sc_hd__nor2_1 _35467_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[6] ),
    .B(net714),
    .Y(_14449_));
 sky130_fd_sc_hd__inv_1 _35468_ (.A(\inst$top.soc.cpu.sink__payload$18[115] ),
    .Y(_14450_));
 sky130_fd_sc_hd__nor2_1 _35469_ (.A(net2839),
    .B(_14450_),
    .Y(_14451_));
 sky130_fd_sc_hd__o21ai_0 _35470_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[6] ),
    .A2(net2003),
    .B1(net2837),
    .Y(_14452_));
 sky130_fd_sc_hd__a21oi_1 _35471_ (.A1(net2004),
    .A2(_14002_),
    .B1(_14452_),
    .Y(_14453_));
 sky130_fd_sc_hd__o21ai_0 _35472_ (.A1(_14451_),
    .A2(_14453_),
    .B1(net2015),
    .Y(_14454_));
 sky130_fd_sc_hd__a21oi_1 _35473_ (.A1(_10322_),
    .A2(net2920),
    .B1(net2010),
    .Y(_14455_));
 sky130_fd_sc_hd__o21ai_2 _35474_ (.A1(net2919),
    .A2(\inst$top.soc.cpu.divider.quotient[6] ),
    .B1(_14455_),
    .Y(_14456_));
 sky130_fd_sc_hd__a21oi_1 _35475_ (.A1(_14454_),
    .A2(net1778),
    .B1(net2831),
    .Y(_14457_));
 sky130_fd_sc_hd__inv_1 _35476_ (.A(_14457_),
    .Y(_14458_));
 sky130_fd_sc_hd__nand2_1 _35477_ (.A(net1797),
    .B(_03131_),
    .Y(_14459_));
 sky130_fd_sc_hd__nand2_1 _35478_ (.A(net1870),
    .B(_03130_),
    .Y(_14460_));
 sky130_fd_sc_hd__o211ai_1 _35479_ (.A1(_03134_),
    .A2(net1232),
    .B1(_14459_),
    .C1(_14460_),
    .Y(_14461_));
 sky130_fd_sc_hd__nand2_1 _35480_ (.A(_13416_),
    .B(net2008),
    .Y(_14462_));
 sky130_fd_sc_hd__o21ai_0 _35481_ (.A1(net2006),
    .A2(_13053_),
    .B1(_14462_),
    .Y(_14463_));
 sky130_fd_sc_hd__xor2_2 _35482_ (.A(_03054_),
    .B(_14463_),
    .X(_14464_));
 sky130_fd_sc_hd__nand2_1 _35483_ (.A(net735),
    .B(net2214),
    .Y(_14465_));
 sky130_fd_sc_hd__nand3_1 _35484_ (.A(_14465_),
    .B(net2018),
    .C(_20610_),
    .Y(_14466_));
 sky130_fd_sc_hd__o21ai_0 _35485_ (.A1(net2018),
    .A2(_14461_),
    .B1(_14466_),
    .Y(_14467_));
 sky130_fd_sc_hd__nand3_1 _35486_ (.A(\inst$top.soc.cpu.sink__payload$12[5] ),
    .B(\inst$top.soc.cpu.sink__payload$12[4] ),
    .C(_03112_),
    .Y(_14468_));
 sky130_fd_sc_hd__xor2_1 _35487_ (.A(\inst$top.soc.cpu.sink__payload$12[6] ),
    .B(_14468_),
    .X(_14469_));
 sky130_fd_sc_hd__mux2i_1 _35488_ (.A0(_14467_),
    .A1(_14469_),
    .S(net2852),
    .Y(_14470_));
 sky130_fd_sc_hd__inv_1 _35489_ (.A(_14470_),
    .Y(_14471_));
 sky130_fd_sc_hd__o22ai_1 _35490_ (.A1(_14458_),
    .A2(net785),
    .B1(_14471_),
    .B2(_12960_),
    .Y(_14472_));
 sky130_fd_sc_hd__a21oi_1 _35491_ (.A1(net739),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[6] ),
    .B1(_14472_),
    .Y(_14473_));
 sky130_fd_sc_hd__nand2_1 _35492_ (.A(net714),
    .B(_14473_),
    .Y(_14474_));
 sky130_fd_sc_hd__nand2_1 _35493_ (.A(_14474_),
    .B(net2175),
    .Y(_14475_));
 sky130_fd_sc_hd__nor2_2 _35494_ (.A(_14449_),
    .B(_14475_),
    .Y(_04212_));
 sky130_fd_sc_hd__nor2_1 _35495_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[7] ),
    .B(net701),
    .Y(_14476_));
 sky130_fd_sc_hd__nor2_1 _35497_ (.A(\inst$top.soc.cpu.sink__payload$12[7] ),
    .B(_13117_),
    .Y(_14478_));
 sky130_fd_sc_hd__o21ai_0 _35498_ (.A1(_20623_),
    .A2(_13288_),
    .B1(net2851),
    .Y(_14479_));
 sky130_fd_sc_hd__inv_1 _35499_ (.A(_03049_),
    .Y(_14480_));
 sky130_fd_sc_hd__a31oi_1 _35500_ (.A1(_13156_),
    .A2(_13133_),
    .A3(_13150_),
    .B1(_13139_),
    .Y(_14481_));
 sky130_fd_sc_hd__nand2_1 _35501_ (.A(_13259_),
    .B(_13168_),
    .Y(_14482_));
 sky130_fd_sc_hd__nand3_1 _35502_ (.A(_14482_),
    .B(net2867),
    .C(_13170_),
    .Y(_14483_));
 sky130_fd_sc_hd__o21ai_0 _35503_ (.A1(net2867),
    .A2(_14481_),
    .B1(_14483_),
    .Y(_14484_));
 sky130_fd_sc_hd__xor2_4 _35504_ (.A(_14480_),
    .B(_14484_),
    .X(_14485_));
 sky130_fd_sc_hd__nand2_1 _35505_ (.A(_14485_),
    .B(net2215),
    .Y(_14486_));
 sky130_fd_sc_hd__nand3_1 _35506_ (.A(_20646_),
    .B(net2017),
    .C(_14486_),
    .Y(_14487_));
 sky130_fd_sc_hd__nor2_1 _35507_ (.A(_03141_),
    .B(net1229),
    .Y(_14488_));
 sky130_fd_sc_hd__a221oi_1 _35508_ (.A1(net1795),
    .A2(_03138_),
    .B1(net1868),
    .B2(_03137_),
    .C1(_14488_),
    .Y(_14489_));
 sky130_fd_sc_hd__a21oi_1 _35509_ (.A1(_14489_),
    .A2(net2862),
    .B1(net2854),
    .Y(_14490_));
 sky130_fd_sc_hd__nand2_1 _35510_ (.A(_14487_),
    .B(_14490_),
    .Y(_14491_));
 sky130_fd_sc_hd__o21ai_1 _35511_ (.A1(_14478_),
    .A2(_14479_),
    .B1(_14491_),
    .Y(_14492_));
 sky130_fd_sc_hd__inv_1 _35512_ (.A(\inst$top.soc.cpu.sink__payload$18[116] ),
    .Y(_14493_));
 sky130_fd_sc_hd__nor2_1 _35513_ (.A(net2834),
    .B(_14493_),
    .Y(_14494_));
 sky130_fd_sc_hd__o21ai_0 _35514_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[7] ),
    .A2(net2003),
    .B1(net2840),
    .Y(_14495_));
 sky130_fd_sc_hd__a21oi_1 _35515_ (.A1(net2003),
    .A2(_13952_),
    .B1(_14495_),
    .Y(_14496_));
 sky130_fd_sc_hd__o21ai_0 _35516_ (.A1(_14494_),
    .A2(_14496_),
    .B1(net2013),
    .Y(_14497_));
 sky130_fd_sc_hd__a21oi_1 _35517_ (.A1(_10323_),
    .A2(net2916),
    .B1(net2009),
    .Y(_14498_));
 sky130_fd_sc_hd__o21ai_1 _35518_ (.A1(net2919),
    .A2(\inst$top.soc.cpu.divider.quotient[7] ),
    .B1(_14498_),
    .Y(_14499_));
 sky130_fd_sc_hd__a21oi_1 _35519_ (.A1(_14497_),
    .A2(net1777),
    .B1(net2829),
    .Y(_14500_));
 sky130_fd_sc_hd__inv_1 _35520_ (.A(_14500_),
    .Y(_14501_));
 sky130_fd_sc_hd__o22ai_1 _35521_ (.A1(_14501_),
    .A2(net783),
    .B1(_20663_),
    .B2(_12956_),
    .Y(_14502_));
 sky130_fd_sc_hd__a21oi_1 _35522_ (.A1(net787),
    .A2(net620),
    .B1(_14502_),
    .Y(_14503_));
 sky130_fd_sc_hd__nand2_1 _35523_ (.A(net709),
    .B(_14503_),
    .Y(_14504_));
 sky130_fd_sc_hd__nand2_1 _35525_ (.A(_14504_),
    .B(net2151),
    .Y(_14506_));
 sky130_fd_sc_hd__nor2_2 _35526_ (.A(_14476_),
    .B(_14506_),
    .Y(_04213_));
 sky130_fd_sc_hd__nor2_1 _35527_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[8] ),
    .B(net712),
    .Y(_14507_));
 sky130_fd_sc_hd__inv_1 _35528_ (.A(\inst$top.soc.cpu.sink__payload$18[117] ),
    .Y(_14508_));
 sky130_fd_sc_hd__nor2_1 _35529_ (.A(net2839),
    .B(_14508_),
    .Y(_14509_));
 sky130_fd_sc_hd__o21ai_0 _35530_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[8] ),
    .A2(net2003),
    .B1(net2837),
    .Y(_14510_));
 sky130_fd_sc_hd__a21oi_1 _35531_ (.A1(net2004),
    .A2(_13903_),
    .B1(_14510_),
    .Y(_14511_));
 sky130_fd_sc_hd__o21ai_0 _35532_ (.A1(_14509_),
    .A2(_14511_),
    .B1(net2015),
    .Y(_14512_));
 sky130_fd_sc_hd__a21oi_1 _35533_ (.A1(_10324_),
    .A2(net2917),
    .B1(net2009),
    .Y(_14513_));
 sky130_fd_sc_hd__o21ai_2 _35534_ (.A1(net2917),
    .A2(\inst$top.soc.cpu.divider.quotient[8] ),
    .B1(_14513_),
    .Y(_14514_));
 sky130_fd_sc_hd__a21oi_1 _35535_ (.A1(_14512_),
    .A2(net1776),
    .B1(net2831),
    .Y(_14515_));
 sky130_fd_sc_hd__inv_1 _35536_ (.A(_14515_),
    .Y(_14516_));
 sky130_fd_sc_hd__nand2_1 _35537_ (.A(_13431_),
    .B(\inst$top.soc.cpu.adder$307.x_sub ),
    .Y(_14517_));
 sky130_fd_sc_hd__o21ai_0 _35538_ (.A1(net2868),
    .A2(_13417_),
    .B1(_14517_),
    .Y(_14518_));
 sky130_fd_sc_hd__xnor2_2 _35539_ (.A(_03044_),
    .B(_14518_),
    .Y(_14519_));
 sky130_fd_sc_hd__o21ai_0 _35540_ (.A1(net2847),
    .A2(net734),
    .B1(_20679_),
    .Y(_14520_));
 sky130_fd_sc_hd__nand2_1 _35541_ (.A(_14520_),
    .B(net2018),
    .Y(_14521_));
 sky130_fd_sc_hd__nand2_1 _35542_ (.A(net1797),
    .B(_03145_),
    .Y(_14522_));
 sky130_fd_sc_hd__nand2_1 _35543_ (.A(net1870),
    .B(_03144_),
    .Y(_14523_));
 sky130_fd_sc_hd__o211ai_1 _35544_ (.A1(_03148_),
    .A2(net1231),
    .B1(_14522_),
    .C1(_14523_),
    .Y(_14524_));
 sky130_fd_sc_hd__a21oi_1 _35545_ (.A1(_14524_),
    .A2(net2861),
    .B1(net2852),
    .Y(_14525_));
 sky130_fd_sc_hd__nand2_1 _35546_ (.A(_13034_),
    .B(_20664_),
    .Y(_14526_));
 sky130_fd_sc_hd__nand2_1 _35547_ (.A(_13033_),
    .B(\inst$top.soc.cpu.sink__payload$12[8] ),
    .Y(_14527_));
 sky130_fd_sc_hd__a21oi_1 _35548_ (.A1(_14526_),
    .A2(_14527_),
    .B1(net2001),
    .Y(_14528_));
 sky130_fd_sc_hd__a21oi_1 _35549_ (.A1(_14521_),
    .A2(_14525_),
    .B1(_14528_),
    .Y(_14529_));
 sky130_fd_sc_hd__inv_1 _35550_ (.A(_14529_),
    .Y(_14530_));
 sky130_fd_sc_hd__o22ai_1 _35551_ (.A1(_14516_),
    .A2(net785),
    .B1(_12960_),
    .B2(_14530_),
    .Y(_14531_));
 sky130_fd_sc_hd__a21oi_1 _35552_ (.A1(net739),
    .A2(net1008),
    .B1(_14531_),
    .Y(_14532_));
 sky130_fd_sc_hd__nand2_1 _35553_ (.A(net712),
    .B(_14532_),
    .Y(_14533_));
 sky130_fd_sc_hd__nand2_1 _35554_ (.A(_14533_),
    .B(net2173),
    .Y(_14534_));
 sky130_fd_sc_hd__nor2_2 _35555_ (.A(_14507_),
    .B(_14534_),
    .Y(_04214_));
 sky130_fd_sc_hd__nor2_1 _35556_ (.A(\inst$top.soc.cpu.gprf.x_bypass1_data[9] ),
    .B(net710),
    .Y(_14535_));
 sky130_fd_sc_hd__inv_1 _35557_ (.A(\inst$top.soc.cpu.sink__payload$18[118] ),
    .Y(_14536_));
 sky130_fd_sc_hd__nor2_1 _35558_ (.A(net2838),
    .B(_14536_),
    .Y(_14537_));
 sky130_fd_sc_hd__o21ai_0 _35559_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[9] ),
    .A2(net2003),
    .B1(net2837),
    .Y(_14538_));
 sky130_fd_sc_hd__a21oi_1 _35560_ (.A1(net2003),
    .A2(_13804_),
    .B1(_14538_),
    .Y(_14539_));
 sky130_fd_sc_hd__o21ai_0 _35561_ (.A1(_14537_),
    .A2(_14539_),
    .B1(net2014),
    .Y(_14540_));
 sky130_fd_sc_hd__a21oi_1 _35562_ (.A1(_10325_),
    .A2(net2916),
    .B1(net2009),
    .Y(_14541_));
 sky130_fd_sc_hd__o21ai_2 _35563_ (.A1(net2917),
    .A2(\inst$top.soc.cpu.divider.quotient[9] ),
    .B1(_14541_),
    .Y(_14542_));
 sky130_fd_sc_hd__a21oi_1 _35564_ (.A1(_14540_),
    .A2(net1775),
    .B1(net2831),
    .Y(_14543_));
 sky130_fd_sc_hd__inv_1 _35565_ (.A(_14543_),
    .Y(_14544_));
 sky130_fd_sc_hd__inv_1 _35566_ (.A(_03039_),
    .Y(_14545_));
 sky130_fd_sc_hd__a21oi_1 _35567_ (.A1(\inst$top.soc.cpu.multiplier.x_prod[0] ),
    .A2(_13491_),
    .B1(_13500_),
    .Y(_14546_));
 sky130_fd_sc_hd__nand2_1 _35568_ (.A(_14546_),
    .B(net2006),
    .Y(_14547_));
 sky130_fd_sc_hd__nand2_1 _35569_ (.A(_13179_),
    .B(net2867),
    .Y(_14548_));
 sky130_fd_sc_hd__nand2_1 _35570_ (.A(_14547_),
    .B(_14548_),
    .Y(_14549_));
 sky130_fd_sc_hd__xor2_2 _35571_ (.A(_14545_),
    .B(_14549_),
    .X(_14550_));
 sky130_fd_sc_hd__o21ai_0 _35572_ (.A1(net2846),
    .A2(net662),
    .B1(_20699_),
    .Y(_14551_));
 sky130_fd_sc_hd__nand2_1 _35573_ (.A(_14551_),
    .B(net2017),
    .Y(_14552_));
 sky130_fd_sc_hd__nand2_1 _35574_ (.A(net1796),
    .B(_03152_),
    .Y(_14553_));
 sky130_fd_sc_hd__nand2_1 _35575_ (.A(net1869),
    .B(_03151_),
    .Y(_14554_));
 sky130_fd_sc_hd__o211ai_1 _35576_ (.A1(_03155_),
    .A2(net1230),
    .B1(_14553_),
    .C1(_14554_),
    .Y(_14555_));
 sky130_fd_sc_hd__a21oi_1 _35577_ (.A1(_14555_),
    .A2(net2861),
    .B1(net2851),
    .Y(_14556_));
 sky130_fd_sc_hd__inv_1 _35578_ (.A(_13289_),
    .Y(_14557_));
 sky130_fd_sc_hd__o21ai_0 _35579_ (.A1(\inst$top.soc.cpu.sink__payload$12[9] ),
    .A2(_14557_),
    .B1(net2851),
    .Y(_14558_));
 sky130_fd_sc_hd__a21oi_1 _35580_ (.A1(\inst$top.soc.cpu.sink__payload$12[9] ),
    .A2(_14557_),
    .B1(_14558_),
    .Y(_14559_));
 sky130_fd_sc_hd__a21oi_1 _35581_ (.A1(_14552_),
    .A2(_14556_),
    .B1(_14559_),
    .Y(_14560_));
 sky130_fd_sc_hd__inv_1 _35582_ (.A(_14560_),
    .Y(_14561_));
 sky130_fd_sc_hd__o22ai_1 _35583_ (.A1(_14544_),
    .A2(net785),
    .B1(net736),
    .B2(_14561_),
    .Y(_14562_));
 sky130_fd_sc_hd__a21oi_1 _35584_ (.A1(net739),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[9] ),
    .B1(_14562_),
    .Y(_14563_));
 sky130_fd_sc_hd__nand2_1 _35585_ (.A(net710),
    .B(_14563_),
    .Y(_14564_));
 sky130_fd_sc_hd__nand2_1 _35586_ (.A(_14564_),
    .B(net2172),
    .Y(_14565_));
 sky130_fd_sc_hd__nor2_2 _35587_ (.A(_14535_),
    .B(_14565_),
    .Y(_04215_));
 sky130_fd_sc_hd__nor2_1 _35588_ (.A(net2886),
    .B(net696),
    .Y(_14566_));
 sky130_fd_sc_hd__a21oi_1 _35589_ (.A1(_20232_),
    .A2(_20330_),
    .B1(_12955_),
    .Y(_14567_));
 sky130_fd_sc_hd__nand3_1 _35590_ (.A(_14567_),
    .B(_20334_),
    .C(_20342_),
    .Y(_14568_));
 sky130_fd_sc_hd__o21ai_1 _35592_ (.A1(_14568_),
    .A2(net652),
    .B1(net2151),
    .Y(_14570_));
 sky130_fd_sc_hd__nor2_4 _35593_ (.A(_14566_),
    .B(_14570_),
    .Y(_04216_));
 sky130_fd_sc_hd__nor2_1 _35594_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[0] ),
    .B(net704),
    .Y(_14571_));
 sky130_fd_sc_hd__nor2_1 _35595_ (.A(\inst$top.soc.cpu.sink__payload$24[34] ),
    .B(net2452),
    .Y(_14572_));
 sky130_fd_sc_hd__nor2_1 _35596_ (.A(net2607),
    .B(_19833_),
    .Y(_14573_));
 sky130_fd_sc_hd__nor2_1 _35597_ (.A(net2597),
    .B(_19834_),
    .Y(_14574_));
 sky130_fd_sc_hd__nor2_1 _35598_ (.A(\inst$top.soc.cpu.sink__payload$24[35] ),
    .B(_06038_),
    .Y(_14575_));
 sky130_fd_sc_hd__nor4_1 _35599_ (.A(_14572_),
    .B(_14573_),
    .C(_14574_),
    .D(_14575_),
    .Y(_14576_));
 sky130_fd_sc_hd__nor2_1 _35600_ (.A(net2652),
    .B(_19836_),
    .Y(_14577_));
 sky130_fd_sc_hd__nor2_1 _35601_ (.A(\inst$top.soc.cpu.sink__payload$24[32] ),
    .B(net2463),
    .Y(_14578_));
 sky130_fd_sc_hd__xor2_1 _35602_ (.A(net2618),
    .B(\inst$top.soc.cpu.sink__payload$24[33] ),
    .X(_14579_));
 sky130_fd_sc_hd__nor3_1 _35603_ (.A(_14577_),
    .B(_14578_),
    .C(_14579_),
    .Y(_14580_));
 sky130_fd_sc_hd__xnor2_1 _35604_ (.A(\inst$top.soc.cpu.sink__payload$24[36] ),
    .B(net2590),
    .Y(_14581_));
 sky130_fd_sc_hd__nand4_1 _35605_ (.A(_14576_),
    .B(_19830_),
    .C(_14580_),
    .D(_14581_),
    .Y(_14582_));
 sky130_fd_sc_hd__nand2_1 _35606_ (.A(_20260_),
    .B(_20240_),
    .Y(_14583_));
 sky130_fd_sc_hd__nor3_1 _35607_ (.A(_20277_),
    .B(_14582_),
    .C(_14583_),
    .Y(_14584_));
 sky130_fd_sc_hd__nor2_2 _35609_ (.A(_20239_),
    .B(_20260_),
    .Y(_14586_));
 sky130_fd_sc_hd__inv_2 _35610_ (.A(net781),
    .Y(_14587_));
 sky130_fd_sc_hd__nand3_1 _35611_ (.A(_20260_),
    .B(_20240_),
    .C(_20277_),
    .Y(_14588_));
 sky130_fd_sc_hd__inv_1 _35612_ (.A(net780),
    .Y(_14589_));
 sky130_fd_sc_hd__nand2_1 _35613_ (.A(net730),
    .B(_13006_),
    .Y(_14590_));
 sky130_fd_sc_hd__o21ai_0 _35614_ (.A1(net731),
    .A2(_12982_),
    .B1(_14590_),
    .Y(_14591_));
 sky130_fd_sc_hd__a21oi_1 _35615_ (.A1(net732),
    .A2(net1064),
    .B1(_14591_),
    .Y(_14592_));
 sky130_fd_sc_hd__nand2_1 _35616_ (.A(net704),
    .B(_14592_),
    .Y(_14593_));
 sky130_fd_sc_hd__nand2_1 _35617_ (.A(_14593_),
    .B(net2152),
    .Y(_14594_));
 sky130_fd_sc_hd__nor2_2 _35618_ (.A(_14571_),
    .B(_14594_),
    .Y(_04217_));
 sky130_fd_sc_hd__nor2_1 _35619_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[10] ),
    .B(net709),
    .Y(_14595_));
 sky130_fd_sc_hd__nand2_1 _35622_ (.A(net730),
    .B(_13026_),
    .Y(_14598_));
 sky130_fd_sc_hd__nand4_1 _35623_ (.A(_14576_),
    .B(_19830_),
    .C(_14580_),
    .D(_14581_),
    .Y(_14599_));
 sky130_fd_sc_hd__nor3_2 _35624_ (.A(_20277_),
    .B(_14599_),
    .C(_14583_),
    .Y(_14600_));
 sky130_fd_sc_hd__nand2_1 _35625_ (.A(net729),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[10] ),
    .Y(_14601_));
 sky130_fd_sc_hd__o211ai_1 _35626_ (.A1(net731),
    .A2(_13095_),
    .B1(_14598_),
    .C1(_14601_),
    .Y(_14602_));
 sky130_fd_sc_hd__o21ai_1 _35628_ (.A1(_14602_),
    .A2(net657),
    .B1(net2156),
    .Y(_14604_));
 sky130_fd_sc_hd__nor2_4 _35629_ (.A(_14595_),
    .B(_14604_),
    .Y(_04218_));
 sky130_fd_sc_hd__nor2_1 _35632_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[11] ),
    .B(net710),
    .Y(_14607_));
 sky130_fd_sc_hd__nand2_1 _35634_ (.A(_13190_),
    .B(net781),
    .Y(_14609_));
 sky130_fd_sc_hd__o21ai_0 _35635_ (.A1(net779),
    .A2(_13113_),
    .B1(_14609_),
    .Y(_14610_));
 sky130_fd_sc_hd__a21oi_1 _35636_ (.A1(net732),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[11] ),
    .B1(_14610_),
    .Y(_14611_));
 sky130_fd_sc_hd__nand2_1 _35637_ (.A(net702),
    .B(_14611_),
    .Y(_14612_));
 sky130_fd_sc_hd__nand2_1 _35638_ (.A(_14612_),
    .B(net2155),
    .Y(_14613_));
 sky130_fd_sc_hd__nor2_4 _35639_ (.A(_14607_),
    .B(_14613_),
    .Y(_04219_));
 sky130_fd_sc_hd__nor2_1 _35640_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[12] ),
    .B(net712),
    .Y(_14614_));
 sky130_fd_sc_hd__nand2_1 _35641_ (.A(_13228_),
    .B(net781),
    .Y(_14615_));
 sky130_fd_sc_hd__nand2_1 _35642_ (.A(_14589_),
    .B(_13238_),
    .Y(_14616_));
 sky130_fd_sc_hd__nand2_1 _35643_ (.A(_14615_),
    .B(_14616_),
    .Y(_14617_));
 sky130_fd_sc_hd__a21oi_1 _35644_ (.A1(net733),
    .A2(net988),
    .B1(_14617_),
    .Y(_14618_));
 sky130_fd_sc_hd__nand2_1 _35645_ (.A(net712),
    .B(_14618_),
    .Y(_14619_));
 sky130_fd_sc_hd__nand2_1 _35646_ (.A(_14619_),
    .B(net2173),
    .Y(_14620_));
 sky130_fd_sc_hd__nor2_4 _35647_ (.A(_14614_),
    .B(_14620_),
    .Y(_04220_));
 sky130_fd_sc_hd__nor2_1 _35648_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[13] ),
    .B(net704),
    .Y(_14621_));
 sky130_fd_sc_hd__nand2_1 _35649_ (.A(net602),
    .B(net781),
    .Y(_14622_));
 sky130_fd_sc_hd__o21ai_0 _35650_ (.A1(net780),
    .A2(_13255_),
    .B1(_14622_),
    .Y(_14623_));
 sky130_fd_sc_hd__a21oi_1 _35651_ (.A1(net732),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[13] ),
    .B1(_14623_),
    .Y(_14624_));
 sky130_fd_sc_hd__nand2_1 _35652_ (.A(net709),
    .B(_14624_),
    .Y(_14625_));
 sky130_fd_sc_hd__nand2_1 _35653_ (.A(_14625_),
    .B(net2152),
    .Y(_14626_));
 sky130_fd_sc_hd__nor2_4 _35654_ (.A(_14621_),
    .B(_14626_),
    .Y(_04221_));
 sky130_fd_sc_hd__nor2_1 _35655_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[14] ),
    .B(net707),
    .Y(_14627_));
 sky130_fd_sc_hd__inv_1 _35656_ (.A(net604),
    .Y(_14628_));
 sky130_fd_sc_hd__nor2_1 _35657_ (.A(_14587_),
    .B(_14628_),
    .Y(_14629_));
 sky130_fd_sc_hd__nor2_1 _35658_ (.A(_20277_),
    .B(_14583_),
    .Y(_14630_));
 sky130_fd_sc_hd__o22ai_1 _35659_ (.A1(net2590),
    .A2(_19826_),
    .B1(_19834_),
    .B2(net2597),
    .Y(_14631_));
 sky130_fd_sc_hd__a2111oi_0 _35660_ (.A1(_19826_),
    .A2(net2590),
    .B1(_14573_),
    .C1(_14575_),
    .D1(_14578_),
    .Y(_14632_));
 sky130_fd_sc_hd__nor2_1 _35661_ (.A(_19829_),
    .B(_14579_),
    .Y(_14633_));
 sky130_fd_sc_hd__nand2_1 _35662_ (.A(_14632_),
    .B(_14633_),
    .Y(_14634_));
 sky130_fd_sc_hd__nor4_1 _35663_ (.A(_14572_),
    .B(_14577_),
    .C(_14631_),
    .D(_14634_),
    .Y(_14635_));
 sky130_fd_sc_hd__nand2_1 _35664_ (.A(_14630_),
    .B(_14635_),
    .Y(_14636_));
 sky130_fd_sc_hd__nand2_1 _35665_ (.A(net730),
    .B(_13348_),
    .Y(_14637_));
 sky130_fd_sc_hd__o21ai_0 _35666_ (.A1(_13339_),
    .A2(_14636_),
    .B1(_14637_),
    .Y(_14638_));
 sky130_fd_sc_hd__nor2_1 _35667_ (.A(_14629_),
    .B(_14638_),
    .Y(_14639_));
 sky130_fd_sc_hd__nand2_1 _35668_ (.A(net706),
    .B(_14639_),
    .Y(_14640_));
 sky130_fd_sc_hd__nand2_1 _35669_ (.A(_14640_),
    .B(net2152),
    .Y(_14641_));
 sky130_fd_sc_hd__nor2_4 _35670_ (.A(_14627_),
    .B(_14641_),
    .Y(_04222_));
 sky130_fd_sc_hd__nor2_1 _35671_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[15] ),
    .B(net705),
    .Y(_14642_));
 sky130_fd_sc_hd__nand2_1 _35673_ (.A(net729),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[15] ),
    .Y(_14644_));
 sky130_fd_sc_hd__nand2_1 _35674_ (.A(net730),
    .B(_13395_),
    .Y(_14645_));
 sky130_fd_sc_hd__nand2_1 _35675_ (.A(_14644_),
    .B(_14645_),
    .Y(_14646_));
 sky130_fd_sc_hd__a21oi_1 _35676_ (.A1(net781),
    .A2(_13387_),
    .B1(_14646_),
    .Y(_14647_));
 sky130_fd_sc_hd__nand2_1 _35677_ (.A(net705),
    .B(_14647_),
    .Y(_14648_));
 sky130_fd_sc_hd__nand2_1 _35678_ (.A(_14648_),
    .B(net2152),
    .Y(_14649_));
 sky130_fd_sc_hd__nor2_4 _35679_ (.A(_14642_),
    .B(_14649_),
    .Y(_04223_));
 sky130_fd_sc_hd__nor2_1 _35680_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[16] ),
    .B(net711),
    .Y(_14650_));
 sky130_fd_sc_hd__nand2_1 _35681_ (.A(_13462_),
    .B(net782),
    .Y(_14651_));
 sky130_fd_sc_hd__o21ai_0 _35682_ (.A1(net780),
    .A2(_13411_),
    .B1(_14651_),
    .Y(_14652_));
 sky130_fd_sc_hd__a21oi_1 _35683_ (.A1(net733),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[16] ),
    .B1(_14652_),
    .Y(_14653_));
 sky130_fd_sc_hd__nand2_1 _35684_ (.A(net710),
    .B(_14653_),
    .Y(_14654_));
 sky130_fd_sc_hd__nand2_1 _35685_ (.A(_14654_),
    .B(net2157),
    .Y(_14655_));
 sky130_fd_sc_hd__nor2_4 _35686_ (.A(_14650_),
    .B(_14655_),
    .Y(_04224_));
 sky130_fd_sc_hd__nor2_1 _35687_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[17] ),
    .B(net713),
    .Y(_14656_));
 sky130_fd_sc_hd__nand2_1 _35689_ (.A(net730),
    .B(_13532_),
    .Y(_14658_));
 sky130_fd_sc_hd__o21ai_0 _35690_ (.A1(_13524_),
    .A2(_14636_),
    .B1(_14658_),
    .Y(_14659_));
 sky130_fd_sc_hd__inv_1 _35691_ (.A(_13523_),
    .Y(_14660_));
 sky130_fd_sc_hd__nor2_1 _35692_ (.A(_14587_),
    .B(_14660_),
    .Y(_14661_));
 sky130_fd_sc_hd__nor2_1 _35693_ (.A(_14659_),
    .B(_14661_),
    .Y(_14662_));
 sky130_fd_sc_hd__nand2_1 _35694_ (.A(net713),
    .B(_14662_),
    .Y(_14663_));
 sky130_fd_sc_hd__nand2_1 _35696_ (.A(_14663_),
    .B(net2173),
    .Y(_14665_));
 sky130_fd_sc_hd__nor2_4 _35697_ (.A(_14656_),
    .B(_14665_),
    .Y(_04225_));
 sky130_fd_sc_hd__nor2_1 _35699_ (.A(_13585_),
    .B(net779),
    .Y(_14667_));
 sky130_fd_sc_hd__a21oi_1 _35700_ (.A1(net729),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[18] ),
    .B1(_14667_),
    .Y(_14668_));
 sky130_fd_sc_hd__o21ai_0 _35701_ (.A1(net731),
    .A2(_13575_),
    .B1(_14668_),
    .Y(_14669_));
 sky130_fd_sc_hd__nand2_1 _35702_ (.A(net704),
    .B(_14669_),
    .Y(_14670_));
 sky130_fd_sc_hd__nand2_1 _35703_ (.A(net656),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[18] ),
    .Y(_14671_));
 sky130_fd_sc_hd__a21oi_4 _35704_ (.A1(_14670_),
    .A2(_14671_),
    .B1(net2994),
    .Y(_04226_));
 sky130_fd_sc_hd__nand2_1 _35707_ (.A(net729),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[19] ),
    .Y(_14674_));
 sky130_fd_sc_hd__nand2_1 _35708_ (.A(_13660_),
    .B(net782),
    .Y(_14675_));
 sky130_fd_sc_hd__o211ai_1 _35709_ (.A1(_14588_),
    .A2(_13606_),
    .B1(_14674_),
    .C1(_14675_),
    .Y(_14676_));
 sky130_fd_sc_hd__nor2_1 _35710_ (.A(net657),
    .B(_14676_),
    .Y(_14677_));
 sky130_fd_sc_hd__nand2_1 _35711_ (.A(net657),
    .B(_20005_),
    .Y(_14678_));
 sky130_fd_sc_hd__nand2_1 _35712_ (.A(_14678_),
    .B(net2172),
    .Y(_14679_));
 sky130_fd_sc_hd__nor2_4 _35713_ (.A(_14677_),
    .B(_14679_),
    .Y(_04227_));
 sky130_fd_sc_hd__nor2_1 _35714_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[1] ),
    .B(net705),
    .Y(_14680_));
 sky130_fd_sc_hd__o22ai_1 _35715_ (.A1(_13676_),
    .A2(net779),
    .B1(_13686_),
    .B2(net731),
    .Y(_14681_));
 sky130_fd_sc_hd__a21oi_1 _35716_ (.A1(net732),
    .A2(net1017),
    .B1(_14681_),
    .Y(_14682_));
 sky130_fd_sc_hd__nand2_1 _35717_ (.A(net705),
    .B(_14682_),
    .Y(_14683_));
 sky130_fd_sc_hd__nand2_1 _35718_ (.A(_14683_),
    .B(net2153),
    .Y(_14684_));
 sky130_fd_sc_hd__nor2_4 _35719_ (.A(_14680_),
    .B(_14684_),
    .Y(_04228_));
 sky130_fd_sc_hd__nand2_1 _35720_ (.A(_13732_),
    .B(net782),
    .Y(_14685_));
 sky130_fd_sc_hd__nand2_1 _35721_ (.A(_14589_),
    .B(_13743_),
    .Y(_14686_));
 sky130_fd_sc_hd__nand2_1 _35722_ (.A(_14600_),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[20] ),
    .Y(_14687_));
 sky130_fd_sc_hd__nand3_1 _35723_ (.A(_14685_),
    .B(_14686_),
    .C(_14687_),
    .Y(_14688_));
 sky130_fd_sc_hd__nand2_1 _35724_ (.A(net714),
    .B(_14688_),
    .Y(_14689_));
 sky130_fd_sc_hd__nand2_1 _35725_ (.A(net659),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[20] ),
    .Y(_14690_));
 sky130_fd_sc_hd__a21oi_4 _35726_ (.A1(_14689_),
    .A2(_14690_),
    .B1(net3003),
    .Y(_04229_));
 sky130_fd_sc_hd__nand2_1 _35727_ (.A(_13793_),
    .B(net782),
    .Y(_14691_));
 sky130_fd_sc_hd__nand2_1 _35728_ (.A(_14600_),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[21] ),
    .Y(_14692_));
 sky130_fd_sc_hd__o211ai_1 _35729_ (.A1(_14588_),
    .A2(_13756_),
    .B1(_14691_),
    .C1(_14692_),
    .Y(_14693_));
 sky130_fd_sc_hd__nand2_1 _35730_ (.A(net712),
    .B(_14693_),
    .Y(_14694_));
 sky130_fd_sc_hd__nand2_1 _35731_ (.A(net659),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[21] ),
    .Y(_14695_));
 sky130_fd_sc_hd__a21oi_4 _35732_ (.A1(_14694_),
    .A2(_14695_),
    .B1(net3003),
    .Y(_04230_));
 sky130_fd_sc_hd__nand2_1 _35733_ (.A(net659),
    .B(_19986_),
    .Y(_14696_));
 sky130_fd_sc_hd__nand2_1 _35734_ (.A(_14696_),
    .B(net2176),
    .Y(_14697_));
 sky130_fd_sc_hd__nand2_1 _35735_ (.A(_14600_),
    .B(net948),
    .Y(_14698_));
 sky130_fd_sc_hd__nand2_1 _35736_ (.A(net603),
    .B(net782),
    .Y(_14699_));
 sky130_fd_sc_hd__o211ai_1 _35737_ (.A1(net780),
    .A2(_13811_),
    .B1(_14698_),
    .C1(_14699_),
    .Y(_14700_));
 sky130_fd_sc_hd__nor2_1 _35738_ (.A(net658),
    .B(_14700_),
    .Y(_14701_));
 sky130_fd_sc_hd__nor2_4 _35739_ (.A(_14697_),
    .B(_14701_),
    .Y(_04231_));
 sky130_fd_sc_hd__nand2_1 _35740_ (.A(_13898_),
    .B(net782),
    .Y(_14702_));
 sky130_fd_sc_hd__nand2_1 _35741_ (.A(net730),
    .B(_13909_),
    .Y(_14703_));
 sky130_fd_sc_hd__nand2_1 _35742_ (.A(_14600_),
    .B(net943),
    .Y(_14704_));
 sky130_fd_sc_hd__nand3_1 _35743_ (.A(_14702_),
    .B(_14703_),
    .C(_14704_),
    .Y(_14705_));
 sky130_fd_sc_hd__nor2_1 _35744_ (.A(net657),
    .B(_14705_),
    .Y(_14706_));
 sky130_fd_sc_hd__nand2_1 _35745_ (.A(net657),
    .B(_19979_),
    .Y(_14707_));
 sky130_fd_sc_hd__nand2_1 _35746_ (.A(_14707_),
    .B(net2172),
    .Y(_14708_));
 sky130_fd_sc_hd__nor2_4 _35747_ (.A(_14706_),
    .B(_14708_),
    .Y(_04232_));
 sky130_fd_sc_hd__nand2_1 _35748_ (.A(_13947_),
    .B(net782),
    .Y(_14709_));
 sky130_fd_sc_hd__nand2_1 _35749_ (.A(net730),
    .B(_13958_),
    .Y(_14710_));
 sky130_fd_sc_hd__nand2_1 _35750_ (.A(net729),
    .B(net938),
    .Y(_14711_));
 sky130_fd_sc_hd__nand3_1 _35751_ (.A(_14709_),
    .B(_14710_),
    .C(_14711_),
    .Y(_14712_));
 sky130_fd_sc_hd__nand2_1 _35752_ (.A(net713),
    .B(_14712_),
    .Y(_14713_));
 sky130_fd_sc_hd__nand2_1 _35753_ (.A(net659),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[24] ),
    .Y(_14714_));
 sky130_fd_sc_hd__a21oi_4 _35754_ (.A1(_14713_),
    .A2(_14714_),
    .B1(net3003),
    .Y(_04233_));
 sky130_fd_sc_hd__inv_1 _35755_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[25] ),
    .Y(_14715_));
 sky130_fd_sc_hd__nand2_1 _35756_ (.A(net650),
    .B(_14715_),
    .Y(_14716_));
 sky130_fd_sc_hd__nand2_1 _35757_ (.A(_14716_),
    .B(net2150),
    .Y(_14717_));
 sky130_fd_sc_hd__nand2_1 _35758_ (.A(_13997_),
    .B(net781),
    .Y(_14718_));
 sky130_fd_sc_hd__nand2_1 _35759_ (.A(net730),
    .B(_14008_),
    .Y(_14719_));
 sky130_fd_sc_hd__nand2_1 _35760_ (.A(net729),
    .B(net933),
    .Y(_14720_));
 sky130_fd_sc_hd__nand3_1 _35761_ (.A(_14718_),
    .B(_14719_),
    .C(_14720_),
    .Y(_14721_));
 sky130_fd_sc_hd__nor2_1 _35762_ (.A(net650),
    .B(_14721_),
    .Y(_14722_));
 sky130_fd_sc_hd__nor2_4 _35763_ (.A(_14717_),
    .B(_14722_),
    .Y(_04234_));
 sky130_fd_sc_hd__nand2_1 _35764_ (.A(_14058_),
    .B(net781),
    .Y(_14723_));
 sky130_fd_sc_hd__nand2_1 _35765_ (.A(net729),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[26] ),
    .Y(_14724_));
 sky130_fd_sc_hd__o211ai_1 _35766_ (.A1(net779),
    .A2(_14021_),
    .B1(_14723_),
    .C1(_14724_),
    .Y(_14725_));
 sky130_fd_sc_hd__nand2_1 _35767_ (.A(net698),
    .B(_14725_),
    .Y(_14726_));
 sky130_fd_sc_hd__nand2_1 _35768_ (.A(net652),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[26] ),
    .Y(_14727_));
 sky130_fd_sc_hd__a21oi_4 _35769_ (.A1(_14726_),
    .A2(_14727_),
    .B1(net2993),
    .Y(_04235_));
 sky130_fd_sc_hd__inv_1 _35770_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[27] ),
    .Y(_14728_));
 sky130_fd_sc_hd__nand2_1 _35771_ (.A(net656),
    .B(_14728_),
    .Y(_14729_));
 sky130_fd_sc_hd__nand2_1 _35772_ (.A(_14729_),
    .B(net2152),
    .Y(_14730_));
 sky130_fd_sc_hd__nand2_1 _35773_ (.A(net729),
    .B(net924),
    .Y(_14731_));
 sky130_fd_sc_hd__nand2_1 _35774_ (.A(_14118_),
    .B(net781),
    .Y(_14732_));
 sky130_fd_sc_hd__o211ai_1 _35775_ (.A1(net780),
    .A2(_14075_),
    .B1(_14731_),
    .C1(_14732_),
    .Y(_14733_));
 sky130_fd_sc_hd__nor2_1 _35776_ (.A(net656),
    .B(_14733_),
    .Y(_14734_));
 sky130_fd_sc_hd__nor2_4 _35777_ (.A(_14730_),
    .B(_14734_),
    .Y(_04236_));
 sky130_fd_sc_hd__nand2_1 _35778_ (.A(_14161_),
    .B(net782),
    .Y(_14735_));
 sky130_fd_sc_hd__nand2_1 _35779_ (.A(net730),
    .B(_14173_),
    .Y(_14736_));
 sky130_fd_sc_hd__nand2_1 _35780_ (.A(net729),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[28] ),
    .Y(_14737_));
 sky130_fd_sc_hd__nand3_1 _35781_ (.A(_14735_),
    .B(_14736_),
    .C(_14737_),
    .Y(_14738_));
 sky130_fd_sc_hd__nand2_1 _35782_ (.A(net711),
    .B(_14738_),
    .Y(_14739_));
 sky130_fd_sc_hd__nand2_1 _35783_ (.A(net660),
    .B(\inst$top.soc.cpu.gprf.x_bypass2_data[28] ),
    .Y(_14740_));
 sky130_fd_sc_hd__a21oi_4 _35784_ (.A1(_14739_),
    .A2(_14740_),
    .B1(net3003),
    .Y(_04237_));
 sky130_fd_sc_hd__nand2_1 _35785_ (.A(net658),
    .B(_19926_),
    .Y(_14741_));
 sky130_fd_sc_hd__nand2_1 _35786_ (.A(_14741_),
    .B(net2176),
    .Y(_14742_));
 sky130_fd_sc_hd__nand2_1 _35787_ (.A(_14225_),
    .B(net782),
    .Y(_14743_));
 sky130_fd_sc_hd__nand2_1 _35788_ (.A(net733),
    .B(net915),
    .Y(_14744_));
 sky130_fd_sc_hd__nand2_1 _35789_ (.A(net730),
    .B(_14236_),
    .Y(_14745_));
 sky130_fd_sc_hd__nand3_1 _35790_ (.A(_14743_),
    .B(_14744_),
    .C(_14745_),
    .Y(_14746_));
 sky130_fd_sc_hd__nor2_1 _35791_ (.A(net658),
    .B(_14746_),
    .Y(_14747_));
 sky130_fd_sc_hd__nor2_4 _35792_ (.A(_14742_),
    .B(_14747_),
    .Y(_04238_));
 sky130_fd_sc_hd__nor2_1 _35793_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[2] ),
    .B(net696),
    .Y(_14748_));
 sky130_fd_sc_hd__o22ai_1 _35794_ (.A1(_14249_),
    .A2(net779),
    .B1(_14261_),
    .B2(net731),
    .Y(_14749_));
 sky130_fd_sc_hd__a21oi_1 _35795_ (.A1(net732),
    .A2(net1063),
    .B1(_14749_),
    .Y(_14750_));
 sky130_fd_sc_hd__nand2_1 _35796_ (.A(net698),
    .B(_14750_),
    .Y(_14751_));
 sky130_fd_sc_hd__nand2_1 _35797_ (.A(_14751_),
    .B(net2150),
    .Y(_14752_));
 sky130_fd_sc_hd__nor2_4 _35798_ (.A(_14748_),
    .B(_14752_),
    .Y(_04239_));
 sky130_fd_sc_hd__nand2_1 _35799_ (.A(net656),
    .B(_19914_),
    .Y(_14753_));
 sky130_fd_sc_hd__nand2_1 _35800_ (.A(_14753_),
    .B(net2152),
    .Y(_14754_));
 sky130_fd_sc_hd__nor2_1 _35801_ (.A(_14277_),
    .B(net779),
    .Y(_14755_));
 sky130_fd_sc_hd__a31oi_1 _35802_ (.A1(_14630_),
    .A2(_14635_),
    .A3(net910),
    .B1(_14755_),
    .Y(_14756_));
 sky130_fd_sc_hd__nand3_1 _35803_ (.A(net665),
    .B(_14756_),
    .C(net755),
    .Y(_14757_));
 sky130_fd_sc_hd__nor2_1 _35804_ (.A(net731),
    .B(_14313_),
    .Y(_14758_));
 sky130_fd_sc_hd__nor2_1 _35805_ (.A(_14757_),
    .B(_14758_),
    .Y(_14759_));
 sky130_fd_sc_hd__nor2_4 _35806_ (.A(_14754_),
    .B(_14759_),
    .Y(_04240_));
 sky130_fd_sc_hd__inv_1 _35807_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[31] ),
    .Y(_14760_));
 sky130_fd_sc_hd__nand2_1 _35808_ (.A(net654),
    .B(_14760_),
    .Y(_14761_));
 sky130_fd_sc_hd__nand2_1 _35809_ (.A(_14761_),
    .B(net2154),
    .Y(_14762_));
 sky130_fd_sc_hd__nor2_1 _35810_ (.A(net731),
    .B(_14349_),
    .Y(_14763_));
 sky130_fd_sc_hd__nor2_1 _35811_ (.A(_14359_),
    .B(net780),
    .Y(_14764_));
 sky130_fd_sc_hd__a31oi_1 _35812_ (.A1(_14630_),
    .A2(_14635_),
    .A3(net905),
    .B1(_14764_),
    .Y(_14765_));
 sky130_fd_sc_hd__nand3_1 _35813_ (.A(net665),
    .B(_14765_),
    .C(net755),
    .Y(_14766_));
 sky130_fd_sc_hd__nor2_1 _35814_ (.A(_14763_),
    .B(_14766_),
    .Y(_14767_));
 sky130_fd_sc_hd__nor2_4 _35815_ (.A(_14762_),
    .B(_14767_),
    .Y(_04241_));
 sky130_fd_sc_hd__nor2_1 _35816_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[3] ),
    .B(net696),
    .Y(_14768_));
 sky130_fd_sc_hd__nand2_1 _35817_ (.A(_14376_),
    .B(net781),
    .Y(_14769_));
 sky130_fd_sc_hd__o21ai_0 _35818_ (.A1(_14385_),
    .A2(net779),
    .B1(_14769_),
    .Y(_14770_));
 sky130_fd_sc_hd__a21oi_1 _35819_ (.A1(net732),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[3] ),
    .B1(_14770_),
    .Y(_14771_));
 sky130_fd_sc_hd__nand2_1 _35820_ (.A(net698),
    .B(_14771_),
    .Y(_14772_));
 sky130_fd_sc_hd__nand2_1 _35821_ (.A(_14772_),
    .B(net2150),
    .Y(_14773_));
 sky130_fd_sc_hd__nor2_4 _35822_ (.A(_14768_),
    .B(_14773_),
    .Y(_04242_));
 sky130_fd_sc_hd__nor2_1 _35824_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[4] ),
    .B(net705),
    .Y(_14775_));
 sky130_fd_sc_hd__o22ai_1 _35825_ (.A1(_14399_),
    .A2(net779),
    .B1(_14413_),
    .B2(net731),
    .Y(_14776_));
 sky130_fd_sc_hd__a21oi_1 _35826_ (.A1(net732),
    .A2(net1013),
    .B1(_14776_),
    .Y(_14777_));
 sky130_fd_sc_hd__nand2_1 _35827_ (.A(net696),
    .B(_14777_),
    .Y(_14778_));
 sky130_fd_sc_hd__nand2_1 _35828_ (.A(_14778_),
    .B(net2151),
    .Y(_14779_));
 sky130_fd_sc_hd__nor2_4 _35829_ (.A(_14775_),
    .B(_14779_),
    .Y(_04243_));
 sky130_fd_sc_hd__nor2_1 _35830_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[5] ),
    .B(net704),
    .Y(_14780_));
 sky130_fd_sc_hd__o22ai_1 _35831_ (.A1(_14427_),
    .A2(net779),
    .B1(_14444_),
    .B2(net731),
    .Y(_14781_));
 sky130_fd_sc_hd__a21oi_1 _35832_ (.A1(net732),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[5] ),
    .B1(_14781_),
    .Y(_14782_));
 sky130_fd_sc_hd__nand2_1 _35833_ (.A(net704),
    .B(_14782_),
    .Y(_14783_));
 sky130_fd_sc_hd__nand2_1 _35834_ (.A(_14783_),
    .B(net2152),
    .Y(_14784_));
 sky130_fd_sc_hd__nor2_4 _35835_ (.A(_14780_),
    .B(_14784_),
    .Y(_04244_));
 sky130_fd_sc_hd__nor2_1 _35836_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[6] ),
    .B(net707),
    .Y(_14785_));
 sky130_fd_sc_hd__o22ai_1 _35837_ (.A1(_14458_),
    .A2(net780),
    .B1(_14471_),
    .B2(net731),
    .Y(_14786_));
 sky130_fd_sc_hd__a21oi_1 _35838_ (.A1(net732),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[6] ),
    .B1(_14786_),
    .Y(_14787_));
 sky130_fd_sc_hd__nand2_1 _35839_ (.A(net707),
    .B(_14787_),
    .Y(_14788_));
 sky130_fd_sc_hd__nand2_1 _35840_ (.A(_14788_),
    .B(net2171),
    .Y(_14789_));
 sky130_fd_sc_hd__nor2_4 _35841_ (.A(_14785_),
    .B(_14789_),
    .Y(_04245_));
 sky130_fd_sc_hd__nor2_1 _35842_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[7] ),
    .B(net705),
    .Y(_14790_));
 sky130_fd_sc_hd__nand2_1 _35843_ (.A(net620),
    .B(net781),
    .Y(_14791_));
 sky130_fd_sc_hd__nand2_1 _35844_ (.A(net729),
    .B(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[7] ),
    .Y(_14792_));
 sky130_fd_sc_hd__o211ai_1 _35845_ (.A1(net779),
    .A2(_14501_),
    .B1(_14791_),
    .C1(_14792_),
    .Y(_14793_));
 sky130_fd_sc_hd__o21ai_1 _35846_ (.A1(_14793_),
    .A2(net656),
    .B1(net2152),
    .Y(_14794_));
 sky130_fd_sc_hd__nor2_4 _35847_ (.A(_14790_),
    .B(_14794_),
    .Y(_04246_));
 sky130_fd_sc_hd__nor2_1 _35848_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[8] ),
    .B(net707),
    .Y(_14795_));
 sky130_fd_sc_hd__inv_1 _35849_ (.A(net1008),
    .Y(_14796_));
 sky130_fd_sc_hd__nor2_1 _35850_ (.A(_14796_),
    .B(_14636_),
    .Y(_14797_));
 sky130_fd_sc_hd__o22ai_1 _35851_ (.A1(_14516_),
    .A2(net780),
    .B1(_14587_),
    .B2(_14530_),
    .Y(_14798_));
 sky130_fd_sc_hd__nor2_1 _35852_ (.A(_14797_),
    .B(_14798_),
    .Y(_14799_));
 sky130_fd_sc_hd__nand2_1 _35853_ (.A(net711),
    .B(_14799_),
    .Y(_14800_));
 sky130_fd_sc_hd__nand2_1 _35854_ (.A(_14800_),
    .B(net2175),
    .Y(_14801_));
 sky130_fd_sc_hd__nor2_4 _35855_ (.A(_14795_),
    .B(_14801_),
    .Y(_04247_));
 sky130_fd_sc_hd__nor2_1 _35856_ (.A(\inst$top.soc.cpu.gprf.x_bypass2_data[9] ),
    .B(net707),
    .Y(_14802_));
 sky130_fd_sc_hd__o22ai_1 _35857_ (.A1(_14544_),
    .A2(net780),
    .B1(_14587_),
    .B2(_14561_),
    .Y(_14803_));
 sky130_fd_sc_hd__a21oi_1 _35858_ (.A1(net732),
    .A2(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[9] ),
    .B1(_14803_),
    .Y(_14804_));
 sky130_fd_sc_hd__nand2_1 _35859_ (.A(net711),
    .B(_14804_),
    .Y(_14805_));
 sky130_fd_sc_hd__nand2_1 _35861_ (.A(_14805_),
    .B(net2171),
    .Y(_14807_));
 sky130_fd_sc_hd__nor2_4 _35862_ (.A(_14802_),
    .B(_14807_),
    .Y(_04248_));
 sky130_fd_sc_hd__nor2_1 _35863_ (.A(net2883),
    .B(net707),
    .Y(_14808_));
 sky130_fd_sc_hd__nand2_1 _35864_ (.A(_14630_),
    .B(_14599_),
    .Y(_14809_));
 sky130_fd_sc_hd__o21ai_1 _35865_ (.A1(_14809_),
    .A2(net656),
    .B1(net2171),
    .Y(_14810_));
 sky130_fd_sc_hd__nor2_4 _35866_ (.A(_14808_),
    .B(_14810_),
    .Y(_04249_));
 sky130_fd_sc_hd__nand3_1 _35867_ (.A(_20364_),
    .B(\inst$top.soc.cpu.d.sink__payload.load ),
    .C(net2238),
    .Y(_14811_));
 sky130_fd_sc_hd__nand2_1 _35868_ (.A(_09837_),
    .B(\inst$top.soc.cpu.d.sink__payload.store ),
    .Y(_14812_));
 sky130_fd_sc_hd__nand2_1 _35869_ (.A(_14811_),
    .B(_14812_),
    .Y(_14813_));
 sky130_fd_sc_hd__clkinv_1 _35870_ (.A(net764),
    .Y(_14814_));
 sky130_fd_sc_hd__nor2_1 _35872_ (.A(net869),
    .B(net728),
    .Y(_14816_));
 sky130_fd_sc_hd__o21ai_0 _35875_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[0] ),
    .A2(net763),
    .B1(net2028),
    .Y(_14819_));
 sky130_fd_sc_hd__nor2_1 _35876_ (.A(_14816_),
    .B(_14819_),
    .Y(_04250_));
 sky130_fd_sc_hd__o21ai_0 _35879_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[10] ),
    .A2(net766),
    .B1(net2027),
    .Y(_14822_));
 sky130_fd_sc_hd__a21oi_2 _35880_ (.A1(_13217_),
    .A2(net765),
    .B1(_14822_),
    .Y(_04251_));
 sky130_fd_sc_hd__nand2_1 _35881_ (.A(_13277_),
    .B(_13278_),
    .Y(_14823_));
 sky130_fd_sc_hd__o21ai_0 _35882_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[11] ),
    .A2(net767),
    .B1(net2049),
    .Y(_14824_));
 sky130_fd_sc_hd__a21oi_2 _35883_ (.A1(_14823_),
    .A2(net767),
    .B1(_14824_),
    .Y(_04252_));
 sky130_fd_sc_hd__o21ai_0 _35884_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[12] ),
    .A2(net767),
    .B1(net2049),
    .Y(_14825_));
 sky130_fd_sc_hd__a21oi_2 _35885_ (.A1(_13327_),
    .A2(net767),
    .B1(_14825_),
    .Y(_04253_));
 sky130_fd_sc_hd__inv_1 _35886_ (.A(_13369_),
    .Y(_14826_));
 sky130_fd_sc_hd__o21ai_0 _35887_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[13] ),
    .A2(net768),
    .B1(net2049),
    .Y(_14827_));
 sky130_fd_sc_hd__a21oi_2 _35888_ (.A1(_14826_),
    .A2(net768),
    .B1(_14827_),
    .Y(_04254_));
 sky130_fd_sc_hd__o21ai_0 _35889_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[14] ),
    .A2(net766),
    .B1(net2027),
    .Y(_14828_));
 sky130_fd_sc_hd__a21oi_2 _35890_ (.A1(_13448_),
    .A2(net765),
    .B1(_14828_),
    .Y(_04255_));
 sky130_fd_sc_hd__o21ai_0 _35892_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[15] ),
    .A2(net767),
    .B1(net2027),
    .Y(_14830_));
 sky130_fd_sc_hd__a21oi_2 _35893_ (.A1(_13515_),
    .A2(net767),
    .B1(_14830_),
    .Y(_04256_));
 sky130_fd_sc_hd__o21ai_0 _35894_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[16] ),
    .A2(net765),
    .B1(net2028),
    .Y(_14831_));
 sky130_fd_sc_hd__a21oi_2 _35895_ (.A1(_13564_),
    .A2(net765),
    .B1(_14831_),
    .Y(_04257_));
 sky130_fd_sc_hd__o21ai_0 _35896_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[17] ),
    .A2(net765),
    .B1(net2027),
    .Y(_14832_));
 sky130_fd_sc_hd__a21oi_2 _35897_ (.A1(_13653_),
    .A2(net765),
    .B1(_14832_),
    .Y(_04258_));
 sky130_fd_sc_hd__o21ai_0 _35899_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[18] ),
    .A2(net765),
    .B1(net2028),
    .Y(_14834_));
 sky130_fd_sc_hd__a21oi_2 _35900_ (.A1(_13729_),
    .A2(net765),
    .B1(_14834_),
    .Y(_04259_));
 sky130_fd_sc_hd__o21ai_0 _35901_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[19] ),
    .A2(net765),
    .B1(net2027),
    .Y(_14835_));
 sky130_fd_sc_hd__a21oi_2 _35902_ (.A1(_13780_),
    .A2(net765),
    .B1(_14835_),
    .Y(_04260_));
 sky130_fd_sc_hd__nor2_1 _35903_ (.A(net830),
    .B(net728),
    .Y(_14836_));
 sky130_fd_sc_hd__o21ai_0 _35904_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[1] ),
    .A2(net763),
    .B1(net2028),
    .Y(_14837_));
 sky130_fd_sc_hd__nor2_1 _35905_ (.A(_14836_),
    .B(_14837_),
    .Y(_04261_));
 sky130_fd_sc_hd__inv_1 _35906_ (.A(_13844_),
    .Y(_14838_));
 sky130_fd_sc_hd__o21ai_0 _35908_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[20] ),
    .A2(net768),
    .B1(net2049),
    .Y(_14840_));
 sky130_fd_sc_hd__a21oi_2 _35909_ (.A1(_14838_),
    .A2(net768),
    .B1(_14840_),
    .Y(_04262_));
 sky130_fd_sc_hd__inv_1 _35910_ (.A(_13890_),
    .Y(_14841_));
 sky130_fd_sc_hd__o21ai_0 _35911_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[21] ),
    .A2(net768),
    .B1(net2050),
    .Y(_14842_));
 sky130_fd_sc_hd__a21oi_2 _35912_ (.A1(_14841_),
    .A2(net768),
    .B1(_14842_),
    .Y(_04263_));
 sky130_fd_sc_hd__inv_1 _35913_ (.A(_13934_),
    .Y(_14843_));
 sky130_fd_sc_hd__o21ai_0 _35914_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[22] ),
    .A2(net768),
    .B1(net2050),
    .Y(_14844_));
 sky130_fd_sc_hd__a21oi_2 _35915_ (.A1(_14843_),
    .A2(net768),
    .B1(_14844_),
    .Y(_04264_));
 sky130_fd_sc_hd__o21ai_0 _35916_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[23] ),
    .A2(net767),
    .B1(net2049),
    .Y(_14845_));
 sky130_fd_sc_hd__a21oi_2 _35917_ (.A1(_13990_),
    .A2(net767),
    .B1(_14845_),
    .Y(_04265_));
 sky130_fd_sc_hd__o21ai_0 _35918_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[24] ),
    .A2(net777),
    .B1(net2060),
    .Y(_14846_));
 sky130_fd_sc_hd__a21oi_2 _35919_ (.A1(_14046_),
    .A2(net777),
    .B1(_14846_),
    .Y(_04266_));
 sky130_fd_sc_hd__and2_1 _35921_ (.A(_14092_),
    .B(_14105_),
    .X(_14848_));
 sky130_fd_sc_hd__nor2_1 _35922_ (.A(_14848_),
    .B(net728),
    .Y(_14849_));
 sky130_fd_sc_hd__a211oi_2 _35923_ (.A1(net728),
    .A2(_09271_),
    .B1(net2948),
    .C1(_14849_),
    .Y(_04267_));
 sky130_fd_sc_hd__inv_1 _35924_ (.A(_14150_),
    .Y(_14850_));
 sky130_fd_sc_hd__o21ai_0 _35926_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[26] ),
    .A2(net777),
    .B1(net2059),
    .Y(_14852_));
 sky130_fd_sc_hd__a21oi_2 _35927_ (.A1(_14850_),
    .A2(net777),
    .B1(_14852_),
    .Y(_04268_));
 sky130_fd_sc_hd__inv_1 _35928_ (.A(_14211_),
    .Y(_14853_));
 sky130_fd_sc_hd__o21ai_0 _35929_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[27] ),
    .A2(net777),
    .B1(net2049),
    .Y(_14854_));
 sky130_fd_sc_hd__a21oi_2 _35930_ (.A1(_14853_),
    .A2(net777),
    .B1(_14854_),
    .Y(_04269_));
 sky130_fd_sc_hd__inv_1 _35931_ (.A(_14300_),
    .Y(_14855_));
 sky130_fd_sc_hd__o21ai_0 _35932_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[28] ),
    .A2(net777),
    .B1(net2049),
    .Y(_14856_));
 sky130_fd_sc_hd__a21oi_2 _35933_ (.A1(_14855_),
    .A2(net777),
    .B1(_14856_),
    .Y(_04270_));
 sky130_fd_sc_hd__inv_2 _35934_ (.A(_14342_),
    .Y(_14857_));
 sky130_fd_sc_hd__o21ai_0 _35936_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[29] ),
    .A2(net763),
    .B1(net2082),
    .Y(_14859_));
 sky130_fd_sc_hd__a21oi_2 _35937_ (.A1(_14857_),
    .A2(net763),
    .B1(_14859_),
    .Y(_04271_));
 sky130_fd_sc_hd__nor2_1 _35938_ (.A(net812),
    .B(net728),
    .Y(_14860_));
 sky130_fd_sc_hd__o21ai_0 _35939_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[2] ),
    .A2(net763),
    .B1(net2028),
    .Y(_14861_));
 sky130_fd_sc_hd__nor2_1 _35940_ (.A(_14860_),
    .B(_14861_),
    .Y(_04272_));
 sky130_fd_sc_hd__o21ai_0 _35941_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[3] ),
    .A2(net763),
    .B1(net2028),
    .Y(_14862_));
 sky130_fd_sc_hd__a21oi_2 _35942_ (.A1(_14434_),
    .A2(net763),
    .B1(_14862_),
    .Y(_04273_));
 sky130_fd_sc_hd__inv_1 _35943_ (.A(net735),
    .Y(_14863_));
 sky130_fd_sc_hd__o21ai_0 _35945_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[4] ),
    .A2(net763),
    .B1(net2028),
    .Y(_14865_));
 sky130_fd_sc_hd__a21oi_2 _35946_ (.A1(_14863_),
    .A2(net764),
    .B1(_14865_),
    .Y(_04274_));
 sky130_fd_sc_hd__inv_1 _35947_ (.A(_14485_),
    .Y(_14866_));
 sky130_fd_sc_hd__o21ai_0 _35948_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[5] ),
    .A2(net763),
    .B1(net2037),
    .Y(_14867_));
 sky130_fd_sc_hd__a21oi_2 _35949_ (.A1(_14866_),
    .A2(net763),
    .B1(_14867_),
    .Y(_04275_));
 sky130_fd_sc_hd__o21ai_0 _35950_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[6] ),
    .A2(net766),
    .B1(net2027),
    .Y(_14868_));
 sky130_fd_sc_hd__a21oi_2 _35951_ (.A1(net734),
    .A2(net766),
    .B1(_14868_),
    .Y(_04276_));
 sky130_fd_sc_hd__o21ai_0 _35952_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[7] ),
    .A2(net766),
    .B1(net2027),
    .Y(_14869_));
 sky130_fd_sc_hd__a21oi_2 _35953_ (.A1(net662),
    .A2(net766),
    .B1(_14869_),
    .Y(_04277_));
 sky130_fd_sc_hd__nand2_1 _35954_ (.A(_13083_),
    .B(_13084_),
    .Y(_14870_));
 sky130_fd_sc_hd__o21ai_0 _35955_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[8] ),
    .A2(net767),
    .B1(net2049),
    .Y(_14871_));
 sky130_fd_sc_hd__a21oi_2 _35956_ (.A1(_14870_),
    .A2(net767),
    .B1(_14871_),
    .Y(_04278_));
 sky130_fd_sc_hd__inv_1 _35957_ (.A(_13187_),
    .Y(_14872_));
 sky130_fd_sc_hd__o21ai_0 _35959_ (.A1(\inst$top.soc.cpu.loadstore.dbus__adr[9] ),
    .A2(net764),
    .B1(net2028),
    .Y(_14874_));
 sky130_fd_sc_hd__a21oi_2 _35960_ (.A1(_14872_),
    .A2(net764),
    .B1(_14874_),
    .Y(_04279_));
 sky130_fd_sc_hd__nand2_1 _35961_ (.A(_12693_),
    .B(net2566),
    .Y(_14875_));
 sky130_fd_sc_hd__nand2_1 _35962_ (.A(_14875_),
    .B(\inst$top.soc.cpu.loadstore.dbus__cyc ),
    .Y(_14876_));
 sky130_fd_sc_hd__a21oi_1 _35963_ (.A1(net727),
    .A2(_14876_),
    .B1(net2949),
    .Y(_04280_));
 sky130_fd_sc_hd__o21ai_0 _35964_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[0] ),
    .A2(net769),
    .B1(net2120),
    .Y(_14877_));
 sky130_fd_sc_hd__nand2_1 _35965_ (.A(_09912_),
    .B(\inst$top.soc.cpu.sink__payload$12[143] ),
    .Y(_14878_));
 sky130_fd_sc_hd__nor2_1 _35966_ (.A(net2842),
    .B(_14878_),
    .Y(_14879_));
 sky130_fd_sc_hd__inv_1 _35967_ (.A(_14879_),
    .Y(_14880_));
 sky130_fd_sc_hd__nand2_1 _35968_ (.A(_14880_),
    .B(_03083_),
    .Y(_14881_));
 sky130_fd_sc_hd__inv_1 _35969_ (.A(net1024),
    .Y(_14882_));
 sky130_fd_sc_hd__nand2_1 _35970_ (.A(_13682_),
    .B(_09912_),
    .Y(_14883_));
 sky130_fd_sc_hd__nor2_1 _35971_ (.A(net2842),
    .B(_14883_),
    .Y(_14884_));
 sky130_fd_sc_hd__inv_1 _35972_ (.A(_14884_),
    .Y(_14885_));
 sky130_fd_sc_hd__nor2_1 _35973_ (.A(\inst$top.soc.cpu.d.sink__payload.csr_fmt_i ),
    .B(_12974_),
    .Y(_14886_));
 sky130_fd_sc_hd__inv_1 _35974_ (.A(net1639),
    .Y(_14887_));
 sky130_fd_sc_hd__o21ai_1 _35975_ (.A1(_14882_),
    .A2(_14885_),
    .B1(net1228),
    .Y(_14888_));
 sky130_fd_sc_hd__a21oi_1 _35976_ (.A1(_20376_),
    .A2(_14888_),
    .B1(net728),
    .Y(_14889_));
 sky130_fd_sc_hd__nor2_1 _35977_ (.A(_14877_),
    .B(_14889_),
    .Y(_04281_));
 sky130_fd_sc_hd__nand2_1 _35980_ (.A(_14879_),
    .B(_20058_),
    .Y(_14892_));
 sky130_fd_sc_hd__o21ai_0 _35981_ (.A1(_20113_),
    .A2(_14881_),
    .B1(_14892_),
    .Y(_14893_));
 sky130_fd_sc_hd__a22oi_1 _35982_ (.A1(_20058_),
    .A2(net1640),
    .B1(_14884_),
    .B2(_14893_),
    .Y(_14894_));
 sky130_fd_sc_hd__o21ai_0 _35983_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[10] ),
    .A2(net769),
    .B1(net2120),
    .Y(_14895_));
 sky130_fd_sc_hd__a21oi_2 _35984_ (.A1(net769),
    .A2(_14894_),
    .B1(_14895_),
    .Y(_04282_));
 sky130_fd_sc_hd__a22o_1 _35985_ (.A1(_20053_),
    .A2(_14879_),
    .B1(_14882_),
    .B2(_20104_),
    .X(_14896_));
 sky130_fd_sc_hd__a22oi_1 _35986_ (.A1(_20053_),
    .A2(net1640),
    .B1(_14896_),
    .B2(_14884_),
    .Y(_14897_));
 sky130_fd_sc_hd__o21ai_0 _35987_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[11] ),
    .A2(net770),
    .B1(net2054),
    .Y(_14898_));
 sky130_fd_sc_hd__a21oi_2 _35988_ (.A1(net770),
    .A2(_14897_),
    .B1(_14898_),
    .Y(_04283_));
 sky130_fd_sc_hd__o2bb2ai_1 _35989_ (.A1_N(_20046_),
    .A2_N(_14879_),
    .B1(_20097_),
    .B2(_14881_),
    .Y(_14899_));
 sky130_fd_sc_hd__a22oi_1 _35990_ (.A1(_20046_),
    .A2(net1640),
    .B1(_14899_),
    .B2(_14884_),
    .Y(_14900_));
 sky130_fd_sc_hd__o21ai_0 _35992_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[12] ),
    .A2(net769),
    .B1(net2120),
    .Y(_14902_));
 sky130_fd_sc_hd__a21oi_2 _35993_ (.A1(net769),
    .A2(_14900_),
    .B1(_14902_),
    .Y(_04284_));
 sky130_fd_sc_hd__nand2_1 _35994_ (.A(_14879_),
    .B(_20040_),
    .Y(_14903_));
 sky130_fd_sc_hd__o21ai_0 _35995_ (.A1(_20090_),
    .A2(net1024),
    .B1(_14903_),
    .Y(_14904_));
 sky130_fd_sc_hd__a22oi_1 _35996_ (.A1(_20040_),
    .A2(net1640),
    .B1(_14884_),
    .B2(_14904_),
    .Y(_14905_));
 sky130_fd_sc_hd__o21ai_0 _35997_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[13] ),
    .A2(net773),
    .B1(net2127),
    .Y(_14906_));
 sky130_fd_sc_hd__a21oi_2 _35998_ (.A1(net773),
    .A2(_14905_),
    .B1(_14906_),
    .Y(_04285_));
 sky130_fd_sc_hd__nand2_1 _36001_ (.A(_14879_),
    .B(_20034_),
    .Y(_14909_));
 sky130_fd_sc_hd__o21ai_0 _36002_ (.A1(_20084_),
    .A2(net1024),
    .B1(_14909_),
    .Y(_14910_));
 sky130_fd_sc_hd__a22oi_1 _36003_ (.A1(_20034_),
    .A2(net1639),
    .B1(_14884_),
    .B2(_14910_),
    .Y(_14911_));
 sky130_fd_sc_hd__o21ai_0 _36004_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[14] ),
    .A2(net777),
    .B1(net2061),
    .Y(_14912_));
 sky130_fd_sc_hd__a21oi_2 _36005_ (.A1(net777),
    .A2(_14911_),
    .B1(_14912_),
    .Y(_04286_));
 sky130_fd_sc_hd__nand2_1 _36006_ (.A(_14879_),
    .B(_20027_),
    .Y(_14913_));
 sky130_fd_sc_hd__o21ai_0 _36007_ (.A1(_20078_),
    .A2(net1024),
    .B1(_14913_),
    .Y(_14914_));
 sky130_fd_sc_hd__a22oi_1 _36008_ (.A1(_20027_),
    .A2(net1640),
    .B1(_14884_),
    .B2(_14914_),
    .Y(_14915_));
 sky130_fd_sc_hd__o21ai_0 _36009_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[15] ),
    .A2(net771),
    .B1(net2061),
    .Y(_14916_));
 sky130_fd_sc_hd__a21oi_2 _36010_ (.A1(net771),
    .A2(_14915_),
    .B1(_14916_),
    .Y(_04287_));
 sky130_fd_sc_hd__nor2_1 _36011_ (.A(\inst$top.soc.cpu.sink__payload$12[144] ),
    .B(_13682_),
    .Y(_14917_));
 sky130_fd_sc_hd__inv_1 _36012_ (.A(_14917_),
    .Y(_14918_));
 sky130_fd_sc_hd__nor2_1 _36013_ (.A(net2842),
    .B(_14918_),
    .Y(_14919_));
 sky130_fd_sc_hd__nor2_1 _36016_ (.A(_20021_),
    .B(net1228),
    .Y(_14922_));
 sky130_fd_sc_hd__a31oi_1 _36017_ (.A1(net811),
    .A2(_20376_),
    .A3(_14881_),
    .B1(_14922_),
    .Y(_14923_));
 sky130_fd_sc_hd__o21ai_0 _36018_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[16] ),
    .A2(net773),
    .B1(net2129),
    .Y(_14924_));
 sky130_fd_sc_hd__a21oi_2 _36019_ (.A1(net774),
    .A2(_14923_),
    .B1(_14924_),
    .Y(_04288_));
 sky130_fd_sc_hd__nor2_1 _36020_ (.A(_20016_),
    .B(net1227),
    .Y(_14925_));
 sky130_fd_sc_hd__a31oi_1 _36021_ (.A1(net811),
    .A2(_20127_),
    .A3(_14881_),
    .B1(_14925_),
    .Y(_14926_));
 sky130_fd_sc_hd__o21ai_0 _36022_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[17] ),
    .A2(net775),
    .B1(net2127),
    .Y(_14927_));
 sky130_fd_sc_hd__a21oi_2 _36023_ (.A1(net775),
    .A2(_14926_),
    .B1(_14927_),
    .Y(_04289_));
 sky130_fd_sc_hd__nor2_1 _36024_ (.A(_20011_),
    .B(net1227),
    .Y(_14928_));
 sky130_fd_sc_hd__a31oi_1 _36025_ (.A1(net811),
    .A2(_20112_),
    .A3(net1024),
    .B1(_14928_),
    .Y(_14929_));
 sky130_fd_sc_hd__o21ai_0 _36026_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[18] ),
    .A2(net773),
    .B1(net2130),
    .Y(_14930_));
 sky130_fd_sc_hd__a21oi_2 _36027_ (.A1(net774),
    .A2(_14929_),
    .B1(_14930_),
    .Y(_04290_));
 sky130_fd_sc_hd__nor2_1 _36028_ (.A(_20007_),
    .B(net1227),
    .Y(_14931_));
 sky130_fd_sc_hd__a31oi_1 _36029_ (.A1(net811),
    .A2(_20104_),
    .A3(net1024),
    .B1(_14931_),
    .Y(_14932_));
 sky130_fd_sc_hd__o21ai_0 _36031_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[19] ),
    .A2(net776),
    .B1(net2130),
    .Y(_14934_));
 sky130_fd_sc_hd__a21oi_2 _36032_ (.A1(net775),
    .A2(_14932_),
    .B1(_14934_),
    .Y(_04291_));
 sky130_fd_sc_hd__o21ai_0 _36033_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[1] ),
    .A2(net770),
    .B1(net2055),
    .Y(_14935_));
 sky130_fd_sc_hd__a21oi_1 _36034_ (.A1(_20127_),
    .A2(_14888_),
    .B1(net727),
    .Y(_14936_));
 sky130_fd_sc_hd__nor2_1 _36035_ (.A(_14935_),
    .B(_14936_),
    .Y(_04292_));
 sky130_fd_sc_hd__nor2_1 _36036_ (.A(net1822),
    .B(net1227),
    .Y(_14937_));
 sky130_fd_sc_hd__a31oi_1 _36037_ (.A1(net811),
    .A2(_20096_),
    .A3(net1024),
    .B1(_14937_),
    .Y(_14938_));
 sky130_fd_sc_hd__o21ai_0 _36038_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[20] ),
    .A2(net774),
    .B1(net2129),
    .Y(_14939_));
 sky130_fd_sc_hd__a21oi_2 _36039_ (.A1(net774),
    .A2(_14938_),
    .B1(_14939_),
    .Y(_04293_));
 sky130_fd_sc_hd__nor2_1 _36040_ (.A(_19995_),
    .B(net1227),
    .Y(_14940_));
 sky130_fd_sc_hd__a31oi_1 _36041_ (.A1(net810),
    .A2(_20089_),
    .A3(net1024),
    .B1(_14940_),
    .Y(_14941_));
 sky130_fd_sc_hd__o21ai_0 _36042_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[21] ),
    .A2(net771),
    .B1(net2062),
    .Y(_14942_));
 sky130_fd_sc_hd__a21oi_2 _36043_ (.A1(net771),
    .A2(_14941_),
    .B1(_14942_),
    .Y(_04294_));
 sky130_fd_sc_hd__nor2_1 _36044_ (.A(net1823),
    .B(net1227),
    .Y(_14943_));
 sky130_fd_sc_hd__a31oi_1 _36045_ (.A1(net810),
    .A2(_20083_),
    .A3(net1024),
    .B1(_14943_),
    .Y(_14944_));
 sky130_fd_sc_hd__o21ai_0 _36047_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[22] ),
    .A2(net774),
    .B1(net2126),
    .Y(_14946_));
 sky130_fd_sc_hd__a21oi_2 _36048_ (.A1(net773),
    .A2(_14944_),
    .B1(_14946_),
    .Y(_04295_));
 sky130_fd_sc_hd__nor2_1 _36049_ (.A(net1824),
    .B(net1227),
    .Y(_14947_));
 sky130_fd_sc_hd__a31oi_1 _36050_ (.A1(net810),
    .A2(_20077_),
    .A3(net1024),
    .B1(_14947_),
    .Y(_14948_));
 sky130_fd_sc_hd__o21ai_0 _36051_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[23] ),
    .A2(net775),
    .B1(net2127),
    .Y(_14949_));
 sky130_fd_sc_hd__a21oi_2 _36052_ (.A1(net775),
    .A2(_14948_),
    .B1(_14949_),
    .Y(_04296_));
 sky130_fd_sc_hd__a22o_1 _36054_ (.A1(_20071_),
    .A2(_14879_),
    .B1(_14882_),
    .B2(_20376_),
    .X(_14951_));
 sky130_fd_sc_hd__nor2_1 _36055_ (.A(_19971_),
    .B(net1228),
    .Y(_14952_));
 sky130_fd_sc_hd__a21oi_1 _36056_ (.A1(_14951_),
    .A2(net810),
    .B1(_14952_),
    .Y(_14953_));
 sky130_fd_sc_hd__o21ai_0 _36057_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[24] ),
    .A2(net772),
    .B1(net2127),
    .Y(_14954_));
 sky130_fd_sc_hd__a21oi_2 _36058_ (.A1(net772),
    .A2(_14953_),
    .B1(_14954_),
    .Y(_04297_));
 sky130_fd_sc_hd__nand2_1 _36059_ (.A(net727),
    .B(\inst$top.soc.cpu.loadstore.dbus__dat_w[25] ),
    .Y(_14955_));
 sky130_fd_sc_hd__a21oi_1 _36060_ (.A1(_19965_),
    .A2(_19964_),
    .B1(net1227),
    .Y(_14956_));
 sky130_fd_sc_hd__a22oi_1 _36061_ (.A1(_20065_),
    .A2(_14879_),
    .B1(_14882_),
    .B2(_20127_),
    .Y(_14957_));
 sky130_fd_sc_hd__nor3_1 _36062_ (.A(net2842),
    .B(_14918_),
    .C(_14957_),
    .Y(_14958_));
 sky130_fd_sc_hd__o21ai_0 _36063_ (.A1(_14956_),
    .A2(_14958_),
    .B1(net772),
    .Y(_14959_));
 sky130_fd_sc_hd__a21oi_1 _36064_ (.A1(_14955_),
    .A2(_14959_),
    .B1(net2982),
    .Y(_04298_));
 sky130_fd_sc_hd__a21oi_1 _36065_ (.A1(_19960_),
    .A2(_19959_),
    .B1(net1227),
    .Y(_14960_));
 sky130_fd_sc_hd__a21oi_1 _36066_ (.A1(net810),
    .A2(_14893_),
    .B1(_14960_),
    .Y(_14961_));
 sky130_fd_sc_hd__o21ai_0 _36067_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[26] ),
    .A2(net769),
    .B1(net2120),
    .Y(_14962_));
 sky130_fd_sc_hd__a21oi_2 _36068_ (.A1(net770),
    .A2(_14961_),
    .B1(_14962_),
    .Y(_04299_));
 sky130_fd_sc_hd__a21oi_1 _36069_ (.A1(_19955_),
    .A2(_19954_),
    .B1(net1227),
    .Y(_14963_));
 sky130_fd_sc_hd__a21oi_1 _36070_ (.A1(_14896_),
    .A2(net810),
    .B1(_14963_),
    .Y(_14964_));
 sky130_fd_sc_hd__o21ai_0 _36071_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[27] ),
    .A2(net773),
    .B1(net2126),
    .Y(_14965_));
 sky130_fd_sc_hd__a21oi_2 _36072_ (.A1(net773),
    .A2(_14964_),
    .B1(_14965_),
    .Y(_04300_));
 sky130_fd_sc_hd__a22oi_1 _36073_ (.A1(_19942_),
    .A2(net1639),
    .B1(net810),
    .B2(_14899_),
    .Y(_14966_));
 sky130_fd_sc_hd__o21ai_0 _36074_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[28] ),
    .A2(net769),
    .B1(net2120),
    .Y(_14967_));
 sky130_fd_sc_hd__a21oi_2 _36075_ (.A1(net770),
    .A2(_14966_),
    .B1(_14967_),
    .Y(_04301_));
 sky130_fd_sc_hd__a22oi_1 _36076_ (.A1(_19928_),
    .A2(net1639),
    .B1(net810),
    .B2(_14904_),
    .Y(_14968_));
 sky130_fd_sc_hd__o21ai_0 _36077_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[29] ),
    .A2(net773),
    .B1(net2126),
    .Y(_14969_));
 sky130_fd_sc_hd__a21oi_2 _36078_ (.A1(net773),
    .A2(_14968_),
    .B1(_14969_),
    .Y(_04302_));
 sky130_fd_sc_hd__o21ai_0 _36079_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[2] ),
    .A2(net772),
    .B1(net2062),
    .Y(_14970_));
 sky130_fd_sc_hd__a21oi_1 _36080_ (.A1(_20112_),
    .A2(_14888_),
    .B1(net727),
    .Y(_14971_));
 sky130_fd_sc_hd__nor2_1 _36081_ (.A(_14970_),
    .B(_14971_),
    .Y(_04303_));
 sky130_fd_sc_hd__a22oi_1 _36082_ (.A1(_19916_),
    .A2(net1639),
    .B1(net810),
    .B2(_14910_),
    .Y(_14972_));
 sky130_fd_sc_hd__o21ai_0 _36083_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[30] ),
    .A2(net771),
    .B1(net2061),
    .Y(_14973_));
 sky130_fd_sc_hd__a21oi_1 _36084_ (.A1(net771),
    .A2(_14972_),
    .B1(_14973_),
    .Y(_04304_));
 sky130_fd_sc_hd__nand2_1 _36085_ (.A(_19893_),
    .B(_19896_),
    .Y(_14974_));
 sky130_fd_sc_hd__a22oi_1 _36086_ (.A1(_14974_),
    .A2(net1639),
    .B1(net810),
    .B2(_14914_),
    .Y(_14975_));
 sky130_fd_sc_hd__o21ai_0 _36087_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[31] ),
    .A2(net775),
    .B1(net2127),
    .Y(_14976_));
 sky130_fd_sc_hd__a21oi_1 _36088_ (.A1(net776),
    .A2(_14975_),
    .B1(_14976_),
    .Y(_04305_));
 sky130_fd_sc_hd__o21ai_0 _36089_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[3] ),
    .A2(net775),
    .B1(net2127),
    .Y(_14977_));
 sky130_fd_sc_hd__a21oi_1 _36090_ (.A1(_20104_),
    .A2(_14888_),
    .B1(net727),
    .Y(_14978_));
 sky130_fd_sc_hd__nor2_1 _36091_ (.A(_14977_),
    .B(_14978_),
    .Y(_04306_));
 sky130_fd_sc_hd__o21ai_0 _36092_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[4] ),
    .A2(net769),
    .B1(net2120),
    .Y(_14979_));
 sky130_fd_sc_hd__a21oi_1 _36093_ (.A1(_20096_),
    .A2(_14888_),
    .B1(net727),
    .Y(_14980_));
 sky130_fd_sc_hd__nor2_1 _36094_ (.A(_14979_),
    .B(_14980_),
    .Y(_04307_));
 sky130_fd_sc_hd__o21ai_0 _36095_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[5] ),
    .A2(net769),
    .B1(net2120),
    .Y(_14981_));
 sky130_fd_sc_hd__a21oi_1 _36096_ (.A1(_20089_),
    .A2(_14888_),
    .B1(net727),
    .Y(_14982_));
 sky130_fd_sc_hd__nor2_1 _36097_ (.A(_14981_),
    .B(_14982_),
    .Y(_04308_));
 sky130_fd_sc_hd__o21ai_0 _36099_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[6] ),
    .A2(net775),
    .B1(net2127),
    .Y(_14984_));
 sky130_fd_sc_hd__a21oi_1 _36100_ (.A1(_20083_),
    .A2(_14888_),
    .B1(net727),
    .Y(_14985_));
 sky130_fd_sc_hd__nor2_1 _36101_ (.A(_14984_),
    .B(_14985_),
    .Y(_04309_));
 sky130_fd_sc_hd__o21ai_0 _36102_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[7] ),
    .A2(net769),
    .B1(net2120),
    .Y(_14986_));
 sky130_fd_sc_hd__a21oi_1 _36103_ (.A1(_20077_),
    .A2(_14888_),
    .B1(net727),
    .Y(_14987_));
 sky130_fd_sc_hd__nor2_1 _36104_ (.A(_14986_),
    .B(_14987_),
    .Y(_04310_));
 sky130_fd_sc_hd__a22oi_1 _36105_ (.A1(_20071_),
    .A2(net1639),
    .B1(_14951_),
    .B2(_14884_),
    .Y(_14988_));
 sky130_fd_sc_hd__o21ai_0 _36106_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[8] ),
    .A2(net771),
    .B1(net2126),
    .Y(_14989_));
 sky130_fd_sc_hd__a21oi_1 _36107_ (.A1(net773),
    .A2(_14988_),
    .B1(_14989_),
    .Y(_04311_));
 sky130_fd_sc_hd__nor2_1 _36108_ (.A(_14885_),
    .B(_14957_),
    .Y(_14990_));
 sky130_fd_sc_hd__a21oi_1 _36109_ (.A1(_20065_),
    .A2(net1639),
    .B1(_14990_),
    .Y(_14991_));
 sky130_fd_sc_hd__o21ai_0 _36112_ (.A1(\inst$top.soc.cpu.loadstore.dbus__dat_w[9] ),
    .A2(net770),
    .B1(net2055),
    .Y(_14994_));
 sky130_fd_sc_hd__a21oi_1 _36113_ (.A1(net770),
    .A2(_14991_),
    .B1(_14994_),
    .Y(_04312_));
 sky130_fd_sc_hd__inv_1 _36114_ (.A(_03083_),
    .Y(_14995_));
 sky130_fd_sc_hd__nand3_1 _36115_ (.A(_13682_),
    .B(_09912_),
    .C(_14995_),
    .Y(_14996_));
 sky130_fd_sc_hd__o21ai_0 _36116_ (.A1(\inst$top.soc.cpu.loadstore.dbus__sel[0] ),
    .A2(net772),
    .B1(net2076),
    .Y(_14997_));
 sky130_fd_sc_hd__a31oi_1 _36117_ (.A1(net772),
    .A2(net1228),
    .A3(_14996_),
    .B1(_14997_),
    .Y(_04313_));
 sky130_fd_sc_hd__nand2_1 _36118_ (.A(_14878_),
    .B(_14995_),
    .Y(_14998_));
 sky130_fd_sc_hd__a31oi_1 _36119_ (.A1(_13682_),
    .A2(_14998_),
    .A3(_09912_),
    .B1(net1639),
    .Y(_14999_));
 sky130_fd_sc_hd__o21ai_0 _36120_ (.A1(\inst$top.soc.cpu.loadstore.dbus__sel[1] ),
    .A2(net772),
    .B1(net2062),
    .Y(_15000_));
 sky130_fd_sc_hd__a21oi_1 _36121_ (.A1(net772),
    .A2(_14999_),
    .B1(_15000_),
    .Y(_04314_));
 sky130_fd_sc_hd__nor2_1 _36122_ (.A(_14995_),
    .B(_14878_),
    .Y(_15001_));
 sky130_fd_sc_hd__o22ai_1 _36123_ (.A1(_14995_),
    .A2(_13682_),
    .B1(_15001_),
    .B2(_14917_),
    .Y(_15002_));
 sky130_fd_sc_hd__o21ai_0 _36124_ (.A1(\inst$top.soc.cpu.loadstore.dbus__sel[2] ),
    .A2(net772),
    .B1(net2076),
    .Y(_15003_));
 sky130_fd_sc_hd__a31oi_1 _36125_ (.A1(net771),
    .A2(net1228),
    .A3(_15002_),
    .B1(_15003_),
    .Y(_04315_));
 sky130_fd_sc_hd__a21oi_1 _36126_ (.A1(_14917_),
    .A2(_14998_),
    .B1(net1639),
    .Y(_15004_));
 sky130_fd_sc_hd__o21ai_0 _36127_ (.A1(\inst$top.soc.cpu.loadstore.dbus__sel[3] ),
    .A2(net771),
    .B1(net2061),
    .Y(_15005_));
 sky130_fd_sc_hd__a21oi_1 _36128_ (.A1(net771),
    .A2(_15004_),
    .B1(_15005_),
    .Y(_04316_));
 sky130_fd_sc_hd__nand2_1 _36129_ (.A(_12693_),
    .B(_09339_),
    .Y(_15006_));
 sky130_fd_sc_hd__nand2_1 _36131_ (.A(net1767),
    .B(\inst$top.soc.cpu.loadstore.dbus__stb ),
    .Y(_15008_));
 sky130_fd_sc_hd__a21oi_1 _36132_ (.A1(net727),
    .A2(_15008_),
    .B1(net2950),
    .Y(_04317_));
 sky130_fd_sc_hd__nand2_1 _36133_ (.A(_14811_),
    .B(\inst$top.soc.cpu.loadstore.dbus__we ),
    .Y(_15009_));
 sky130_fd_sc_hd__a21oi_1 _36135_ (.A1(_15009_),
    .A2(_14812_),
    .B1(net2955),
    .Y(_04318_));
 sky130_fd_sc_hd__inv_1 _36138_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[0] ),
    .Y(_15013_));
 sky130_fd_sc_hd__a21oi_1 _36139_ (.A1(net1768),
    .A2(_15013_),
    .B1(net2980),
    .Y(_15014_));
 sky130_fd_sc_hd__o21ai_0 _36140_ (.A1(net1767),
    .A2(_12713_),
    .B1(_15014_),
    .Y(_15015_));
 sky130_fd_sc_hd__inv_2 _36141_ (.A(_15015_),
    .Y(_04319_));
 sky130_fd_sc_hd__inv_1 _36142_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[10] ),
    .Y(_15016_));
 sky130_fd_sc_hd__a21oi_1 _36143_ (.A1(net1768),
    .A2(_15016_),
    .B1(net2980),
    .Y(_15017_));
 sky130_fd_sc_hd__o21ai_0 _36144_ (.A1(net1767),
    .A2(_12725_),
    .B1(_15017_),
    .Y(_15018_));
 sky130_fd_sc_hd__inv_2 _36145_ (.A(_15018_),
    .Y(_04320_));
 sky130_fd_sc_hd__inv_1 _36146_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[11] ),
    .Y(_15019_));
 sky130_fd_sc_hd__a21oi_1 _36147_ (.A1(net1770),
    .A2(_15019_),
    .B1(net2980),
    .Y(_15020_));
 sky130_fd_sc_hd__o21ai_0 _36148_ (.A1(net1770),
    .A2(_12732_),
    .B1(_15020_),
    .Y(_15021_));
 sky130_fd_sc_hd__inv_2 _36149_ (.A(_15021_),
    .Y(_04321_));
 sky130_fd_sc_hd__inv_1 _36150_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[12] ),
    .Y(_15022_));
 sky130_fd_sc_hd__a21oi_1 _36152_ (.A1(net1770),
    .A2(_15022_),
    .B1(net2980),
    .Y(_15024_));
 sky130_fd_sc_hd__o21ai_0 _36153_ (.A1(net1770),
    .A2(_12739_),
    .B1(_15024_),
    .Y(_15025_));
 sky130_fd_sc_hd__inv_2 _36154_ (.A(_15025_),
    .Y(_04322_));
 sky130_fd_sc_hd__inv_1 _36155_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[13] ),
    .Y(_15026_));
 sky130_fd_sc_hd__a21oi_1 _36156_ (.A1(net1772),
    .A2(_15026_),
    .B1(net2990),
    .Y(_15027_));
 sky130_fd_sc_hd__o21ai_0 _36157_ (.A1(net1773),
    .A2(_12746_),
    .B1(_15027_),
    .Y(_15028_));
 sky130_fd_sc_hd__inv_2 _36158_ (.A(_15028_),
    .Y(_04323_));
 sky130_fd_sc_hd__inv_1 _36159_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[14] ),
    .Y(_15029_));
 sky130_fd_sc_hd__a21oi_1 _36160_ (.A1(net1773),
    .A2(_15029_),
    .B1(net2990),
    .Y(_15030_));
 sky130_fd_sc_hd__o21ai_0 _36161_ (.A1(net1771),
    .A2(_12753_),
    .B1(_15030_),
    .Y(_15031_));
 sky130_fd_sc_hd__inv_2 _36162_ (.A(_15031_),
    .Y(_04324_));
 sky130_fd_sc_hd__inv_1 _36163_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[15] ),
    .Y(_15032_));
 sky130_fd_sc_hd__a21oi_1 _36164_ (.A1(net1769),
    .A2(_15032_),
    .B1(net2988),
    .Y(_15033_));
 sky130_fd_sc_hd__o21ai_0 _36165_ (.A1(net1769),
    .A2(_12761_),
    .B1(_15033_),
    .Y(_15034_));
 sky130_fd_sc_hd__inv_2 _36166_ (.A(_15034_),
    .Y(_04325_));
 sky130_fd_sc_hd__inv_1 _36167_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[16] ),
    .Y(_15035_));
 sky130_fd_sc_hd__a21oi_1 _36168_ (.A1(net1772),
    .A2(_15035_),
    .B1(net2989),
    .Y(_15036_));
 sky130_fd_sc_hd__o21ai_0 _36169_ (.A1(net1772),
    .A2(_12768_),
    .B1(_15036_),
    .Y(_15037_));
 sky130_fd_sc_hd__inv_2 _36170_ (.A(_15037_),
    .Y(_04326_));
 sky130_fd_sc_hd__inv_1 _36172_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[17] ),
    .Y(_15039_));
 sky130_fd_sc_hd__a21oi_1 _36173_ (.A1(net1772),
    .A2(_15039_),
    .B1(net2990),
    .Y(_15040_));
 sky130_fd_sc_hd__o21ai_0 _36174_ (.A1(net1772),
    .A2(_12775_),
    .B1(_15040_),
    .Y(_15041_));
 sky130_fd_sc_hd__inv_2 _36175_ (.A(_15041_),
    .Y(_04327_));
 sky130_fd_sc_hd__inv_1 _36176_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[18] ),
    .Y(_15042_));
 sky130_fd_sc_hd__a21oi_1 _36177_ (.A1(net1769),
    .A2(_15042_),
    .B1(net2988),
    .Y(_15043_));
 sky130_fd_sc_hd__o21ai_0 _36178_ (.A1(net1769),
    .A2(_12783_),
    .B1(_15043_),
    .Y(_15044_));
 sky130_fd_sc_hd__inv_2 _36179_ (.A(_15044_),
    .Y(_04328_));
 sky130_fd_sc_hd__inv_1 _36181_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[19] ),
    .Y(_15046_));
 sky130_fd_sc_hd__a21oi_1 _36182_ (.A1(net1772),
    .A2(_15046_),
    .B1(net2990),
    .Y(_15047_));
 sky130_fd_sc_hd__o21ai_0 _36183_ (.A1(net1772),
    .A2(_12793_),
    .B1(_15047_),
    .Y(_15048_));
 sky130_fd_sc_hd__inv_2 _36184_ (.A(_15048_),
    .Y(_04329_));
 sky130_fd_sc_hd__inv_1 _36185_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[1] ),
    .Y(_15049_));
 sky130_fd_sc_hd__a21oi_1 _36186_ (.A1(net1770),
    .A2(_15049_),
    .B1(net2980),
    .Y(_15050_));
 sky130_fd_sc_hd__o21ai_0 _36187_ (.A1(net1770),
    .A2(_12800_),
    .B1(_15050_),
    .Y(_15051_));
 sky130_fd_sc_hd__inv_2 _36188_ (.A(_15051_),
    .Y(_04330_));
 sky130_fd_sc_hd__inv_1 _36189_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[20] ),
    .Y(_15052_));
 sky130_fd_sc_hd__a21oi_1 _36190_ (.A1(net1771),
    .A2(_15052_),
    .B1(net2988),
    .Y(_15053_));
 sky130_fd_sc_hd__o21ai_0 _36191_ (.A1(net1769),
    .A2(_12807_),
    .B1(_15053_),
    .Y(_15054_));
 sky130_fd_sc_hd__inv_2 _36192_ (.A(_15054_),
    .Y(_04331_));
 sky130_fd_sc_hd__inv_1 _36193_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[21] ),
    .Y(_15055_));
 sky130_fd_sc_hd__a21oi_1 _36195_ (.A1(net1771),
    .A2(_15055_),
    .B1(net2989),
    .Y(_15057_));
 sky130_fd_sc_hd__o21ai_0 _36196_ (.A1(net1771),
    .A2(_12814_),
    .B1(_15057_),
    .Y(_15058_));
 sky130_fd_sc_hd__inv_2 _36197_ (.A(_15058_),
    .Y(_04332_));
 sky130_fd_sc_hd__inv_1 _36198_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[22] ),
    .Y(_15059_));
 sky130_fd_sc_hd__a21oi_1 _36199_ (.A1(net1771),
    .A2(_15059_),
    .B1(net2989),
    .Y(_15060_));
 sky130_fd_sc_hd__o21ai_0 _36200_ (.A1(net1771),
    .A2(_12821_),
    .B1(_15060_),
    .Y(_15061_));
 sky130_fd_sc_hd__inv_2 _36201_ (.A(_15061_),
    .Y(_04333_));
 sky130_fd_sc_hd__inv_1 _36202_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[23] ),
    .Y(_15062_));
 sky130_fd_sc_hd__a21oi_1 _36203_ (.A1(net1769),
    .A2(_15062_),
    .B1(net2988),
    .Y(_15063_));
 sky130_fd_sc_hd__o21ai_0 _36204_ (.A1(net1769),
    .A2(_12828_),
    .B1(_15063_),
    .Y(_15064_));
 sky130_fd_sc_hd__inv_2 _36205_ (.A(_15064_),
    .Y(_04334_));
 sky130_fd_sc_hd__inv_1 _36206_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[24] ),
    .Y(_15065_));
 sky130_fd_sc_hd__a21oi_1 _36207_ (.A1(net1771),
    .A2(_15065_),
    .B1(net2990),
    .Y(_15066_));
 sky130_fd_sc_hd__o21ai_0 _36208_ (.A1(net1771),
    .A2(net3038),
    .B1(_15066_),
    .Y(_15067_));
 sky130_fd_sc_hd__inv_2 _36209_ (.A(_15067_),
    .Y(_04335_));
 sky130_fd_sc_hd__inv_1 _36210_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[25] ),
    .Y(_15068_));
 sky130_fd_sc_hd__a21oi_1 _36211_ (.A1(net1769),
    .A2(_15068_),
    .B1(net2988),
    .Y(_15069_));
 sky130_fd_sc_hd__o21ai_0 _36212_ (.A1(net1774),
    .A2(_12843_),
    .B1(_15069_),
    .Y(_15070_));
 sky130_fd_sc_hd__inv_2 _36213_ (.A(_15070_),
    .Y(_04336_));
 sky130_fd_sc_hd__inv_1 _36215_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[26] ),
    .Y(_15072_));
 sky130_fd_sc_hd__a21oi_1 _36216_ (.A1(net1774),
    .A2(_15072_),
    .B1(net2988),
    .Y(_15073_));
 sky130_fd_sc_hd__o21ai_0 _36217_ (.A1(net1769),
    .A2(net3037),
    .B1(_15073_),
    .Y(_15074_));
 sky130_fd_sc_hd__inv_2 _36218_ (.A(_15074_),
    .Y(_04337_));
 sky130_fd_sc_hd__inv_1 _36219_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[27] ),
    .Y(_15075_));
 sky130_fd_sc_hd__a21oi_1 _36220_ (.A1(net1768),
    .A2(_15075_),
    .B1(net2982),
    .Y(_15076_));
 sky130_fd_sc_hd__o21ai_0 _36221_ (.A1(net1768),
    .A2(_12858_),
    .B1(_15076_),
    .Y(_15077_));
 sky130_fd_sc_hd__inv_2 _36222_ (.A(_15077_),
    .Y(_04338_));
 sky130_fd_sc_hd__inv_1 _36224_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[28] ),
    .Y(_15079_));
 sky130_fd_sc_hd__a21oi_1 _36225_ (.A1(net1768),
    .A2(_15079_),
    .B1(net2980),
    .Y(_15080_));
 sky130_fd_sc_hd__o21ai_0 _36226_ (.A1(net1768),
    .A2(_12866_),
    .B1(_15080_),
    .Y(_15081_));
 sky130_fd_sc_hd__inv_2 _36227_ (.A(_15081_),
    .Y(_04339_));
 sky130_fd_sc_hd__inv_1 _36228_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[29] ),
    .Y(_15082_));
 sky130_fd_sc_hd__a21oi_1 _36229_ (.A1(net1772),
    .A2(_15082_),
    .B1(net2990),
    .Y(_15083_));
 sky130_fd_sc_hd__o21ai_0 _36230_ (.A1(net1772),
    .A2(net3041),
    .B1(_15083_),
    .Y(_15084_));
 sky130_fd_sc_hd__inv_2 _36231_ (.A(_15084_),
    .Y(_04340_));
 sky130_fd_sc_hd__inv_1 _36232_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[2] ),
    .Y(_15085_));
 sky130_fd_sc_hd__a21oi_1 _36233_ (.A1(net1767),
    .A2(_15085_),
    .B1(net2982),
    .Y(_15086_));
 sky130_fd_sc_hd__o21ai_0 _36234_ (.A1(net1767),
    .A2(_12880_),
    .B1(_15086_),
    .Y(_15087_));
 sky130_fd_sc_hd__inv_2 _36235_ (.A(_15087_),
    .Y(_04341_));
 sky130_fd_sc_hd__inv_1 _36236_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[30] ),
    .Y(_15088_));
 sky130_fd_sc_hd__a21oi_1 _36238_ (.A1(net1772),
    .A2(_15088_),
    .B1(net2990),
    .Y(_15090_));
 sky130_fd_sc_hd__o21ai_0 _36239_ (.A1(net1773),
    .A2(net3040),
    .B1(_15090_),
    .Y(_15091_));
 sky130_fd_sc_hd__inv_2 _36240_ (.A(_15091_),
    .Y(_04342_));
 sky130_fd_sc_hd__inv_1 _36241_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[31] ),
    .Y(_15092_));
 sky130_fd_sc_hd__a21oi_1 _36242_ (.A1(net1770),
    .A2(_15092_),
    .B1(net2991),
    .Y(_15093_));
 sky130_fd_sc_hd__o21ai_0 _36243_ (.A1(net1770),
    .A2(_12894_),
    .B1(_15093_),
    .Y(_15094_));
 sky130_fd_sc_hd__inv_2 _36244_ (.A(_15094_),
    .Y(_04343_));
 sky130_fd_sc_hd__inv_1 _36245_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[3] ),
    .Y(_15095_));
 sky130_fd_sc_hd__a21oi_1 _36246_ (.A1(net1767),
    .A2(_15095_),
    .B1(net2982),
    .Y(_15096_));
 sky130_fd_sc_hd__o21ai_0 _36247_ (.A1(net1767),
    .A2(_12901_),
    .B1(_15096_),
    .Y(_15097_));
 sky130_fd_sc_hd__inv_2 _36248_ (.A(_15097_),
    .Y(_04344_));
 sky130_fd_sc_hd__inv_1 _36249_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[4] ),
    .Y(_15098_));
 sky130_fd_sc_hd__a21oi_1 _36250_ (.A1(net1767),
    .A2(_15098_),
    .B1(net2982),
    .Y(_15099_));
 sky130_fd_sc_hd__o21ai_0 _36251_ (.A1(net1767),
    .A2(_12909_),
    .B1(_15099_),
    .Y(_15100_));
 sky130_fd_sc_hd__inv_2 _36252_ (.A(_15100_),
    .Y(_04345_));
 sky130_fd_sc_hd__inv_1 _36253_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[5] ),
    .Y(_15101_));
 sky130_fd_sc_hd__a21oi_1 _36254_ (.A1(net1774),
    .A2(_15101_),
    .B1(net2991),
    .Y(_15102_));
 sky130_fd_sc_hd__o21ai_0 _36255_ (.A1(net1770),
    .A2(_12916_),
    .B1(_15102_),
    .Y(_15103_));
 sky130_fd_sc_hd__inv_2 _36256_ (.A(_15103_),
    .Y(_04346_));
 sky130_fd_sc_hd__inv_1 _36257_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[6] ),
    .Y(_15104_));
 sky130_fd_sc_hd__a21oi_1 _36258_ (.A1(net1773),
    .A2(_15104_),
    .B1(net2990),
    .Y(_15105_));
 sky130_fd_sc_hd__o21ai_0 _36259_ (.A1(net1773),
    .A2(_12923_),
    .B1(_15105_),
    .Y(_15106_));
 sky130_fd_sc_hd__inv_2 _36260_ (.A(_15106_),
    .Y(_04347_));
 sky130_fd_sc_hd__inv_1 _36261_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[7] ),
    .Y(_15107_));
 sky130_fd_sc_hd__a21oi_1 _36262_ (.A1(net1769),
    .A2(_15107_),
    .B1(net2991),
    .Y(_15108_));
 sky130_fd_sc_hd__o21ai_0 _36263_ (.A1(net1774),
    .A2(net3039),
    .B1(_15108_),
    .Y(_15109_));
 sky130_fd_sc_hd__inv_2 _36264_ (.A(_15109_),
    .Y(_04348_));
 sky130_fd_sc_hd__inv_1 _36265_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[8] ),
    .Y(_15110_));
 sky130_fd_sc_hd__a21oi_1 _36266_ (.A1(net1767),
    .A2(_15110_),
    .B1(net2981),
    .Y(_15111_));
 sky130_fd_sc_hd__o21ai_0 _36267_ (.A1(net1768),
    .A2(_12937_),
    .B1(_15111_),
    .Y(_15112_));
 sky130_fd_sc_hd__inv_2 _36268_ (.A(_15112_),
    .Y(_04349_));
 sky130_fd_sc_hd__inv_1 _36269_ (.A(\inst$top.soc.cpu.loadstore.m_load_data[9] ),
    .Y(_15113_));
 sky130_fd_sc_hd__a21oi_1 _36270_ (.A1(net1771),
    .A2(_15113_),
    .B1(net2991),
    .Y(_15114_));
 sky130_fd_sc_hd__o21ai_0 _36271_ (.A1(net1771),
    .A2(_12944_),
    .B1(_15114_),
    .Y(_15115_));
 sky130_fd_sc_hd__inv_2 _36272_ (.A(_15115_),
    .Y(_04350_));
 sky130_fd_sc_hd__nand2_1 _36273_ (.A(net2029),
    .B(\inst$top.soc.cpu.x.source__valid ),
    .Y(_15116_));
 sky130_fd_sc_hd__nor2_1 _36274_ (.A(_15116_),
    .B(net1881),
    .Y(_04351_));
 sky130_fd_sc_hd__nor2_1 _36275_ (.A(\inst$top.soc.cpu.multiplier.x_low ),
    .B(net1914),
    .Y(_15117_));
 sky130_fd_sc_hd__o21ai_0 _36278_ (.A1(\inst$top.soc.cpu.multiplier.m_low ),
    .A2(net2279),
    .B1(net2155),
    .Y(_15120_));
 sky130_fd_sc_hd__nor2_1 _36279_ (.A(_15117_),
    .B(_15120_),
    .Y(_04352_));
 sky130_fd_sc_hd__o21ai_0 _36280_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[0] ),
    .A2(net2282),
    .B1(net2177),
    .Y(_15121_));
 sky130_fd_sc_hd__a21oi_1 _36281_ (.A1(_00162_),
    .A2(net2282),
    .B1(_15121_),
    .Y(_04353_));
 sky130_fd_sc_hd__inv_1 _36284_ (.A(_03409_),
    .Y(_15124_));
 sky130_fd_sc_hd__a21oi_1 _36285_ (.A1(_03387_),
    .A2(_03379_),
    .B1(_03386_),
    .Y(_15125_));
 sky130_fd_sc_hd__nand3_1 _36286_ (.A(_02547_),
    .B(_02915_),
    .C(_03387_),
    .Y(_15126_));
 sky130_fd_sc_hd__nand2_1 _36287_ (.A(_15125_),
    .B(_15126_),
    .Y(_15127_));
 sky130_fd_sc_hd__nand2_1 _36288_ (.A(_03393_),
    .B(_03402_),
    .Y(_15128_));
 sky130_fd_sc_hd__inv_1 _36289_ (.A(_15128_),
    .Y(_15129_));
 sky130_fd_sc_hd__nand2_1 _36290_ (.A(_03402_),
    .B(_03392_),
    .Y(_15130_));
 sky130_fd_sc_hd__inv_1 _36291_ (.A(_03401_),
    .Y(_15131_));
 sky130_fd_sc_hd__nand2_1 _36292_ (.A(_15130_),
    .B(_15131_),
    .Y(_15132_));
 sky130_fd_sc_hd__a21oi_1 _36293_ (.A1(_15127_),
    .A2(_15129_),
    .B1(_15132_),
    .Y(_15133_));
 sky130_fd_sc_hd__xor2_1 _36294_ (.A(_15124_),
    .B(_15133_),
    .X(_15134_));
 sky130_fd_sc_hd__nor2_1 _36295_ (.A(\inst$top.soc.cpu.multiplier.m_prod[10] ),
    .B(net2300),
    .Y(_15135_));
 sky130_fd_sc_hd__nor2_1 _36296_ (.A(net3009),
    .B(_15135_),
    .Y(_15136_));
 sky130_fd_sc_hd__o21ai_0 _36297_ (.A1(net1922),
    .A2(_15134_),
    .B1(_15136_),
    .Y(_15137_));
 sky130_fd_sc_hd__inv_2 _36298_ (.A(_15137_),
    .Y(_04354_));
 sky130_fd_sc_hd__a21oi_1 _36299_ (.A1(_03393_),
    .A2(_03386_),
    .B1(_03392_),
    .Y(_15138_));
 sky130_fd_sc_hd__nand3_1 _36300_ (.A(_02548_),
    .B(_03387_),
    .C(_03393_),
    .Y(_15139_));
 sky130_fd_sc_hd__nand2_1 _36301_ (.A(_15138_),
    .B(_15139_),
    .Y(_15140_));
 sky130_fd_sc_hd__nand2_1 _36302_ (.A(_03402_),
    .B(_03409_),
    .Y(_15141_));
 sky130_fd_sc_hd__inv_1 _36303_ (.A(_15141_),
    .Y(_15142_));
 sky130_fd_sc_hd__o21bai_1 _36304_ (.A1(_15124_),
    .A2(_15131_),
    .B1_N(_03408_),
    .Y(_15143_));
 sky130_fd_sc_hd__a21oi_1 _36305_ (.A1(_15140_),
    .A2(_15142_),
    .B1(_15143_),
    .Y(_15144_));
 sky130_fd_sc_hd__xnor2_1 _36306_ (.A(_03414_),
    .B(_15144_),
    .Y(_15145_));
 sky130_fd_sc_hd__nor2_1 _36308_ (.A(\inst$top.soc.cpu.multiplier.m_prod[11] ),
    .B(net2300),
    .Y(_15147_));
 sky130_fd_sc_hd__nor2_1 _36309_ (.A(net3009),
    .B(_15147_),
    .Y(_15148_));
 sky130_fd_sc_hd__o21ai_0 _36310_ (.A1(net1922),
    .A2(_15145_),
    .B1(_15148_),
    .Y(_15149_));
 sky130_fd_sc_hd__inv_2 _36311_ (.A(_15149_),
    .Y(_04355_));
 sky130_fd_sc_hd__nand2_1 _36312_ (.A(_03409_),
    .B(_03414_),
    .Y(_15150_));
 sky130_fd_sc_hd__a21oi_1 _36313_ (.A1(_03414_),
    .A2(_03408_),
    .B1(_03413_),
    .Y(_15151_));
 sky130_fd_sc_hd__o21ai_1 _36314_ (.A1(_15150_),
    .A2(_15133_),
    .B1(_15151_),
    .Y(_15152_));
 sky130_fd_sc_hd__xor2_1 _36315_ (.A(_03420_),
    .B(net601),
    .X(_15153_));
 sky130_fd_sc_hd__nor2_1 _36316_ (.A(\inst$top.soc.cpu.multiplier.m_prod[12] ),
    .B(net2301),
    .Y(_15154_));
 sky130_fd_sc_hd__nor2_1 _36317_ (.A(net3007),
    .B(_15154_),
    .Y(_15155_));
 sky130_fd_sc_hd__o21ai_0 _36318_ (.A1(net1921),
    .A2(_15153_),
    .B1(_15155_),
    .Y(_15156_));
 sky130_fd_sc_hd__inv_2 _36319_ (.A(_15156_),
    .Y(_04356_));
 sky130_fd_sc_hd__nand2_1 _36320_ (.A(_03414_),
    .B(_03420_),
    .Y(_15157_));
 sky130_fd_sc_hd__a21oi_1 _36321_ (.A1(_03420_),
    .A2(_03413_),
    .B1(_03419_),
    .Y(_15158_));
 sky130_fd_sc_hd__o21ai_1 _36322_ (.A1(_15157_),
    .A2(_15144_),
    .B1(_15158_),
    .Y(_15159_));
 sky130_fd_sc_hd__xor2_1 _36323_ (.A(_03427_),
    .B(_15159_),
    .X(_15160_));
 sky130_fd_sc_hd__nor2_1 _36324_ (.A(\inst$top.soc.cpu.multiplier.m_prod[13] ),
    .B(net2301),
    .Y(_15161_));
 sky130_fd_sc_hd__nor2_1 _36325_ (.A(net3007),
    .B(_15161_),
    .Y(_15162_));
 sky130_fd_sc_hd__o21ai_0 _36326_ (.A1(net1921),
    .A2(_15160_),
    .B1(_15162_),
    .Y(_15163_));
 sky130_fd_sc_hd__inv_2 _36327_ (.A(_15163_),
    .Y(_04357_));
 sky130_fd_sc_hd__inv_1 _36328_ (.A(_03433_),
    .Y(_15164_));
 sky130_fd_sc_hd__nand2_1 _36329_ (.A(_03427_),
    .B(_03419_),
    .Y(_15165_));
 sky130_fd_sc_hd__inv_1 _36330_ (.A(_03426_),
    .Y(_15166_));
 sky130_fd_sc_hd__nand2_1 _36331_ (.A(_15165_),
    .B(_15166_),
    .Y(_15167_));
 sky130_fd_sc_hd__a31oi_1 _36332_ (.A1(net601),
    .A2(_03420_),
    .A3(_03427_),
    .B1(_15167_),
    .Y(_15168_));
 sky130_fd_sc_hd__xor2_1 _36333_ (.A(_15164_),
    .B(_15168_),
    .X(_15169_));
 sky130_fd_sc_hd__nor2_1 _36334_ (.A(\inst$top.soc.cpu.multiplier.m_prod[14] ),
    .B(net2301),
    .Y(_15170_));
 sky130_fd_sc_hd__nor2_1 _36335_ (.A(net3009),
    .B(_15170_),
    .Y(_15171_));
 sky130_fd_sc_hd__o21ai_0 _36336_ (.A1(net1921),
    .A2(_15169_),
    .B1(_15171_),
    .Y(_15172_));
 sky130_fd_sc_hd__inv_2 _36337_ (.A(_15172_),
    .Y(_04358_));
 sky130_fd_sc_hd__inv_1 _36338_ (.A(_03443_),
    .Y(_15173_));
 sky130_fd_sc_hd__inv_1 _36339_ (.A(_03432_),
    .Y(_15174_));
 sky130_fd_sc_hd__o21ai_0 _36340_ (.A1(_15164_),
    .A2(_15166_),
    .B1(_15174_),
    .Y(_15175_));
 sky130_fd_sc_hd__a31oi_1 _36341_ (.A1(_15159_),
    .A2(_03427_),
    .A3(_03433_),
    .B1(_15175_),
    .Y(_15176_));
 sky130_fd_sc_hd__xor2_1 _36342_ (.A(_15173_),
    .B(_15176_),
    .X(_15177_));
 sky130_fd_sc_hd__nor2_1 _36343_ (.A(\inst$top.soc.cpu.multiplier.m_prod[15] ),
    .B(net2300),
    .Y(_15178_));
 sky130_fd_sc_hd__nor2_1 _36344_ (.A(net3007),
    .B(_15178_),
    .Y(_15179_));
 sky130_fd_sc_hd__o21ai_0 _36345_ (.A1(net1921),
    .A2(_15177_),
    .B1(_15179_),
    .Y(_15180_));
 sky130_fd_sc_hd__inv_2 _36346_ (.A(_15180_),
    .Y(_04359_));
 sky130_fd_sc_hd__inv_1 _36347_ (.A(_03455_),
    .Y(_15181_));
 sky130_fd_sc_hd__nand2_1 _36348_ (.A(_03420_),
    .B(_03427_),
    .Y(_15182_));
 sky130_fd_sc_hd__nand2_1 _36349_ (.A(_03433_),
    .B(_03443_),
    .Y(_15183_));
 sky130_fd_sc_hd__nor2_1 _36350_ (.A(_15182_),
    .B(_15183_),
    .Y(_15184_));
 sky130_fd_sc_hd__nand2_1 _36351_ (.A(net601),
    .B(_15184_),
    .Y(_15185_));
 sky130_fd_sc_hd__inv_1 _36352_ (.A(_03442_),
    .Y(_15186_));
 sky130_fd_sc_hd__o21ai_0 _36353_ (.A1(_15173_),
    .A2(_15174_),
    .B1(_15186_),
    .Y(_15187_));
 sky130_fd_sc_hd__a31oi_1 _36354_ (.A1(_15167_),
    .A2(_03433_),
    .A3(_03443_),
    .B1(_15187_),
    .Y(_15188_));
 sky130_fd_sc_hd__nand2_1 _36355_ (.A(_15185_),
    .B(_15188_),
    .Y(_15189_));
 sky130_fd_sc_hd__nor2_1 _36356_ (.A(_15181_),
    .B(_15189_),
    .Y(_15190_));
 sky130_fd_sc_hd__nand2_1 _36357_ (.A(_15189_),
    .B(_15181_),
    .Y(_15191_));
 sky130_fd_sc_hd__nand2_1 _36358_ (.A(_15191_),
    .B(net2305),
    .Y(_15192_));
 sky130_fd_sc_hd__o221ai_1 _36359_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[16] ),
    .A2(net2305),
    .B1(_15190_),
    .B2(_15192_),
    .C1(net2184),
    .Y(_15193_));
 sky130_fd_sc_hd__inv_2 _36360_ (.A(_15193_),
    .Y(_04360_));
 sky130_fd_sc_hd__inv_1 _36361_ (.A(_03464_),
    .Y(_15194_));
 sky130_fd_sc_hd__nand2_1 _36362_ (.A(_03427_),
    .B(_03433_),
    .Y(_15195_));
 sky130_fd_sc_hd__nand2_1 _36363_ (.A(_03443_),
    .B(_03455_),
    .Y(_15196_));
 sky130_fd_sc_hd__nor2_1 _36364_ (.A(_15195_),
    .B(_15196_),
    .Y(_15197_));
 sky130_fd_sc_hd__nand2_1 _36365_ (.A(_15159_),
    .B(_15197_),
    .Y(_15198_));
 sky130_fd_sc_hd__inv_1 _36366_ (.A(_03454_),
    .Y(_15199_));
 sky130_fd_sc_hd__o21ai_0 _36367_ (.A1(_15181_),
    .A2(_15186_),
    .B1(_15199_),
    .Y(_15200_));
 sky130_fd_sc_hd__a31oi_1 _36368_ (.A1(_15175_),
    .A2(_03443_),
    .A3(_03455_),
    .B1(_15200_),
    .Y(_15201_));
 sky130_fd_sc_hd__nand2_1 _36369_ (.A(_15198_),
    .B(_15201_),
    .Y(_15202_));
 sky130_fd_sc_hd__nor2_1 _36370_ (.A(_15194_),
    .B(_15202_),
    .Y(_15203_));
 sky130_fd_sc_hd__nand2_1 _36371_ (.A(_15202_),
    .B(_15194_),
    .Y(_15204_));
 sky130_fd_sc_hd__nand2_1 _36372_ (.A(_15204_),
    .B(net2305),
    .Y(_15205_));
 sky130_fd_sc_hd__o221ai_1 _36374_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[17] ),
    .A2(net2305),
    .B1(_15203_),
    .B2(_15205_),
    .C1(net2184),
    .Y(_15207_));
 sky130_fd_sc_hd__inv_2 _36375_ (.A(_15207_),
    .Y(_04361_));
 sky130_fd_sc_hd__inv_1 _36377_ (.A(_03476_),
    .Y(_15209_));
 sky130_fd_sc_hd__nand2_1 _36378_ (.A(_03464_),
    .B(_03455_),
    .Y(_15210_));
 sky130_fd_sc_hd__inv_1 _36379_ (.A(_15210_),
    .Y(_15211_));
 sky130_fd_sc_hd__inv_1 _36380_ (.A(_03463_),
    .Y(_15212_));
 sky130_fd_sc_hd__o21ai_0 _36381_ (.A1(_15194_),
    .A2(_15199_),
    .B1(_15212_),
    .Y(_15213_));
 sky130_fd_sc_hd__a21oi_1 _36382_ (.A1(_15189_),
    .A2(_15211_),
    .B1(_15213_),
    .Y(_15214_));
 sky130_fd_sc_hd__inv_1 _36383_ (.A(_15214_),
    .Y(_15215_));
 sky130_fd_sc_hd__nor2_1 _36384_ (.A(_15209_),
    .B(_15215_),
    .Y(_15216_));
 sky130_fd_sc_hd__o21ai_0 _36385_ (.A1(_03476_),
    .A2(_15214_),
    .B1(net2305),
    .Y(_15217_));
 sky130_fd_sc_hd__o221ai_1 _36386_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[18] ),
    .A2(net2305),
    .B1(_15216_),
    .B2(_15217_),
    .C1(net2180),
    .Y(_15218_));
 sky130_fd_sc_hd__inv_2 _36387_ (.A(_15218_),
    .Y(_04362_));
 sky130_fd_sc_hd__inv_1 _36388_ (.A(_03487_),
    .Y(_15219_));
 sky130_fd_sc_hd__nand2_1 _36389_ (.A(_03476_),
    .B(_03464_),
    .Y(_15220_));
 sky130_fd_sc_hd__inv_1 _36390_ (.A(_15220_),
    .Y(_15221_));
 sky130_fd_sc_hd__inv_1 _36391_ (.A(_03475_),
    .Y(_15222_));
 sky130_fd_sc_hd__o21ai_0 _36392_ (.A1(_15209_),
    .A2(_15212_),
    .B1(_15222_),
    .Y(_15223_));
 sky130_fd_sc_hd__a21oi_1 _36393_ (.A1(_15202_),
    .A2(_15221_),
    .B1(_15223_),
    .Y(_15224_));
 sky130_fd_sc_hd__inv_1 _36394_ (.A(_15224_),
    .Y(_15225_));
 sky130_fd_sc_hd__nor2_1 _36395_ (.A(_15219_),
    .B(_15225_),
    .Y(_15226_));
 sky130_fd_sc_hd__o21ai_0 _36396_ (.A1(_03487_),
    .A2(_15224_),
    .B1(net2306),
    .Y(_15227_));
 sky130_fd_sc_hd__o221ai_1 _36397_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[19] ),
    .A2(net2306),
    .B1(_15226_),
    .B2(_15227_),
    .C1(net2184),
    .Y(_15228_));
 sky130_fd_sc_hd__inv_2 _36398_ (.A(_15228_),
    .Y(_04363_));
 sky130_fd_sc_hd__nor2_1 _36399_ (.A(\inst$top.soc.cpu.multiplier.x_prod[1] ),
    .B(net1922),
    .Y(_15229_));
 sky130_fd_sc_hd__o21ai_0 _36400_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[1] ),
    .A2(net2299),
    .B1(net2179),
    .Y(_15230_));
 sky130_fd_sc_hd__nor2_1 _36401_ (.A(_15229_),
    .B(_15230_),
    .Y(_04364_));
 sky130_fd_sc_hd__inv_1 _36402_ (.A(_03496_),
    .Y(_15231_));
 sky130_fd_sc_hd__nand2_1 _36403_ (.A(_03476_),
    .B(_03487_),
    .Y(_15232_));
 sky130_fd_sc_hd__nor2_1 _36404_ (.A(_15210_),
    .B(_15232_),
    .Y(_15233_));
 sky130_fd_sc_hd__inv_1 _36405_ (.A(_15232_),
    .Y(_15234_));
 sky130_fd_sc_hd__inv_1 _36406_ (.A(_03486_),
    .Y(_15235_));
 sky130_fd_sc_hd__o21ai_0 _36407_ (.A1(_15219_),
    .A2(_15222_),
    .B1(_15235_),
    .Y(_15236_));
 sky130_fd_sc_hd__a21oi_1 _36408_ (.A1(_15213_),
    .A2(_15234_),
    .B1(_15236_),
    .Y(_15237_));
 sky130_fd_sc_hd__inv_1 _36409_ (.A(_15237_),
    .Y(_15238_));
 sky130_fd_sc_hd__a21oi_1 _36410_ (.A1(_15189_),
    .A2(_15233_),
    .B1(_15238_),
    .Y(_15239_));
 sky130_fd_sc_hd__inv_1 _36411_ (.A(_15239_),
    .Y(_15240_));
 sky130_fd_sc_hd__nor2_1 _36412_ (.A(_15231_),
    .B(_15240_),
    .Y(_15241_));
 sky130_fd_sc_hd__o21ai_0 _36413_ (.A1(_03496_),
    .A2(_15239_),
    .B1(net2307),
    .Y(_15242_));
 sky130_fd_sc_hd__o221ai_1 _36414_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[20] ),
    .A2(net2307),
    .B1(_15241_),
    .B2(_15242_),
    .C1(net2184),
    .Y(_15243_));
 sky130_fd_sc_hd__inv_2 _36415_ (.A(_15243_),
    .Y(_04365_));
 sky130_fd_sc_hd__inv_1 _36416_ (.A(_03508_),
    .Y(_15244_));
 sky130_fd_sc_hd__nand2_1 _36417_ (.A(_03487_),
    .B(_03496_),
    .Y(_15245_));
 sky130_fd_sc_hd__inv_1 _36418_ (.A(_15245_),
    .Y(_15246_));
 sky130_fd_sc_hd__o21bai_1 _36419_ (.A1(_15231_),
    .A2(_15235_),
    .B1_N(_03495_),
    .Y(_15247_));
 sky130_fd_sc_hd__a21oi_1 _36420_ (.A1(_15225_),
    .A2(_15246_),
    .B1(_15247_),
    .Y(_15248_));
 sky130_fd_sc_hd__inv_1 _36421_ (.A(_15248_),
    .Y(_15249_));
 sky130_fd_sc_hd__nor2_1 _36422_ (.A(_15244_),
    .B(_15249_),
    .Y(_15250_));
 sky130_fd_sc_hd__o21ai_0 _36423_ (.A1(_03508_),
    .A2(_15248_),
    .B1(net2307),
    .Y(_15251_));
 sky130_fd_sc_hd__o221ai_1 _36424_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[21] ),
    .A2(net2307),
    .B1(_15250_),
    .B2(_15251_),
    .C1(net2184),
    .Y(_15252_));
 sky130_fd_sc_hd__inv_2 _36425_ (.A(_15252_),
    .Y(_04366_));
 sky130_fd_sc_hd__nand2_1 _36426_ (.A(_03496_),
    .B(_03508_),
    .Y(_15253_));
 sky130_fd_sc_hd__a21oi_1 _36427_ (.A1(_03508_),
    .A2(_03495_),
    .B1(_03507_),
    .Y(_15254_));
 sky130_fd_sc_hd__o21ai_0 _36428_ (.A1(_15253_),
    .A2(_15239_),
    .B1(_15254_),
    .Y(_15255_));
 sky130_fd_sc_hd__xor2_1 _36429_ (.A(_03522_),
    .B(_15255_),
    .X(_15256_));
 sky130_fd_sc_hd__nor2_1 _36430_ (.A(\inst$top.soc.cpu.multiplier.m_prod[22] ),
    .B(net2309),
    .Y(_15257_));
 sky130_fd_sc_hd__nor2_1 _36431_ (.A(net3013),
    .B(_15257_),
    .Y(_15258_));
 sky130_fd_sc_hd__o21ai_0 _36432_ (.A1(net1930),
    .A2(_15256_),
    .B1(_15258_),
    .Y(_15259_));
 sky130_fd_sc_hd__inv_2 _36433_ (.A(_15259_),
    .Y(_04367_));
 sky130_fd_sc_hd__inv_1 _36434_ (.A(_03533_),
    .Y(_15260_));
 sky130_fd_sc_hd__nand2_1 _36435_ (.A(_03508_),
    .B(_03522_),
    .Y(_15261_));
 sky130_fd_sc_hd__nor2_1 _36436_ (.A(_15245_),
    .B(_15261_),
    .Y(_15262_));
 sky130_fd_sc_hd__nand2_1 _36437_ (.A(_15225_),
    .B(_15262_),
    .Y(_15263_));
 sky130_fd_sc_hd__inv_1 _36438_ (.A(_15261_),
    .Y(_15264_));
 sky130_fd_sc_hd__a21oi_1 _36439_ (.A1(_03522_),
    .A2(_03507_),
    .B1(_03521_),
    .Y(_15265_));
 sky130_fd_sc_hd__inv_1 _36440_ (.A(_15265_),
    .Y(_15266_));
 sky130_fd_sc_hd__a21oi_1 _36441_ (.A1(_15247_),
    .A2(_15264_),
    .B1(_15266_),
    .Y(_15267_));
 sky130_fd_sc_hd__nand2_1 _36442_ (.A(_15263_),
    .B(_15267_),
    .Y(_15268_));
 sky130_fd_sc_hd__nor2_1 _36443_ (.A(_15260_),
    .B(_15268_),
    .Y(_15269_));
 sky130_fd_sc_hd__nand2_1 _36444_ (.A(_15268_),
    .B(_15260_),
    .Y(_15270_));
 sky130_fd_sc_hd__nand2_1 _36445_ (.A(_15270_),
    .B(net2309),
    .Y(_15271_));
 sky130_fd_sc_hd__o221ai_1 _36446_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[23] ),
    .A2(net2309),
    .B1(_15269_),
    .B2(_15271_),
    .C1(net2186),
    .Y(_15272_));
 sky130_fd_sc_hd__inv_2 _36447_ (.A(_15272_),
    .Y(_04368_));
 sky130_fd_sc_hd__nand2_1 _36448_ (.A(_03522_),
    .B(_03533_),
    .Y(_15273_));
 sky130_fd_sc_hd__nor2_1 _36449_ (.A(_15253_),
    .B(_15273_),
    .Y(_15274_));
 sky130_fd_sc_hd__a21oi_1 _36450_ (.A1(_03533_),
    .A2(_03521_),
    .B1(_03532_),
    .Y(_15275_));
 sky130_fd_sc_hd__o21ai_0 _36451_ (.A1(_15273_),
    .A2(_15254_),
    .B1(_15275_),
    .Y(_15276_));
 sky130_fd_sc_hd__a21oi_1 _36452_ (.A1(_15240_),
    .A2(_15274_),
    .B1(_15276_),
    .Y(_15277_));
 sky130_fd_sc_hd__xnor2_1 _36453_ (.A(_03546_),
    .B(_15277_),
    .Y(_15278_));
 sky130_fd_sc_hd__nor2_1 _36455_ (.A(\inst$top.soc.cpu.multiplier.m_prod[24] ),
    .B(net2307),
    .Y(_15280_));
 sky130_fd_sc_hd__nor2_1 _36456_ (.A(net3012),
    .B(_15280_),
    .Y(_15281_));
 sky130_fd_sc_hd__o21ai_0 _36457_ (.A1(net1928),
    .A2(_15278_),
    .B1(_15281_),
    .Y(_15282_));
 sky130_fd_sc_hd__inv_2 _36458_ (.A(_15282_),
    .Y(_04369_));
 sky130_fd_sc_hd__nand2_1 _36460_ (.A(_03533_),
    .B(_03546_),
    .Y(_15284_));
 sky130_fd_sc_hd__inv_1 _36461_ (.A(_15284_),
    .Y(_15285_));
 sky130_fd_sc_hd__a21oi_1 _36462_ (.A1(_03546_),
    .A2(_03532_),
    .B1(_03545_),
    .Y(_15286_));
 sky130_fd_sc_hd__a21boi_0 _36463_ (.A1(_15268_),
    .A2(_15285_),
    .B1_N(_15286_),
    .Y(_15287_));
 sky130_fd_sc_hd__xnor2_1 _36464_ (.A(_03558_),
    .B(_15287_),
    .Y(_15288_));
 sky130_fd_sc_hd__nor2_1 _36465_ (.A(\inst$top.soc.cpu.multiplier.m_prod[25] ),
    .B(net2309),
    .Y(_15289_));
 sky130_fd_sc_hd__nor2_1 _36466_ (.A(net3013),
    .B(_15289_),
    .Y(_15290_));
 sky130_fd_sc_hd__o21ai_0 _36467_ (.A1(net1931),
    .A2(_15288_),
    .B1(_15290_),
    .Y(_15291_));
 sky130_fd_sc_hd__inv_2 _36468_ (.A(_15291_),
    .Y(_04370_));
 sky130_fd_sc_hd__nand2_1 _36469_ (.A(_03546_),
    .B(_03558_),
    .Y(_15292_));
 sky130_fd_sc_hd__a21oi_1 _36470_ (.A1(_03558_),
    .A2(_03545_),
    .B1(_03557_),
    .Y(_15293_));
 sky130_fd_sc_hd__o21ai_0 _36471_ (.A1(_15292_),
    .A2(_15277_),
    .B1(_15293_),
    .Y(_15294_));
 sky130_fd_sc_hd__xor2_1 _36472_ (.A(_03570_),
    .B(_15294_),
    .X(_15295_));
 sky130_fd_sc_hd__nor2_1 _36473_ (.A(\inst$top.soc.cpu.multiplier.m_prod[26] ),
    .B(net2306),
    .Y(_15296_));
 sky130_fd_sc_hd__nor2_1 _36474_ (.A(net3012),
    .B(_15296_),
    .Y(_15297_));
 sky130_fd_sc_hd__o21ai_0 _36475_ (.A1(net1928),
    .A2(_15295_),
    .B1(_15297_),
    .Y(_15298_));
 sky130_fd_sc_hd__inv_2 _36476_ (.A(_15298_),
    .Y(_04371_));
 sky130_fd_sc_hd__nand2_1 _36477_ (.A(_03558_),
    .B(_03570_),
    .Y(_15299_));
 sky130_fd_sc_hd__a21oi_1 _36478_ (.A1(_03570_),
    .A2(_03557_),
    .B1(_03569_),
    .Y(_15300_));
 sky130_fd_sc_hd__o21ai_0 _36479_ (.A1(_15299_),
    .A2(_15287_),
    .B1(_15300_),
    .Y(_15301_));
 sky130_fd_sc_hd__xor2_1 _36480_ (.A(_03582_),
    .B(_15301_),
    .X(_15302_));
 sky130_fd_sc_hd__nor2_1 _36481_ (.A(\inst$top.soc.cpu.multiplier.m_prod[27] ),
    .B(net2306),
    .Y(_15303_));
 sky130_fd_sc_hd__nor2_1 _36482_ (.A(net3007),
    .B(_15303_),
    .Y(_15304_));
 sky130_fd_sc_hd__o21ai_0 _36483_ (.A1(net1928),
    .A2(_15302_),
    .B1(_15304_),
    .Y(_15305_));
 sky130_fd_sc_hd__inv_2 _36484_ (.A(_15305_),
    .Y(_04372_));
 sky130_fd_sc_hd__inv_1 _36485_ (.A(_15233_),
    .Y(_15306_));
 sky130_fd_sc_hd__nand2_1 _36486_ (.A(_03570_),
    .B(_03582_),
    .Y(_15307_));
 sky130_fd_sc_hd__nor2_1 _36487_ (.A(_15292_),
    .B(_15307_),
    .Y(_15308_));
 sky130_fd_sc_hd__nand2_1 _36488_ (.A(_15274_),
    .B(_15308_),
    .Y(_15309_));
 sky130_fd_sc_hd__nor4_1 _36489_ (.A(_15182_),
    .B(_15183_),
    .C(_15306_),
    .D(_15309_),
    .Y(_15310_));
 sky130_fd_sc_hd__nor2_1 _36490_ (.A(_15306_),
    .B(_15188_),
    .Y(_15311_));
 sky130_fd_sc_hd__nor2_1 _36491_ (.A(_15238_),
    .B(_15311_),
    .Y(_15312_));
 sky130_fd_sc_hd__a21oi_1 _36492_ (.A1(_03582_),
    .A2(_03569_),
    .B1(_03581_),
    .Y(_15313_));
 sky130_fd_sc_hd__o21ai_0 _36493_ (.A1(_15307_),
    .A2(_15293_),
    .B1(_15313_),
    .Y(_15314_));
 sky130_fd_sc_hd__a21oi_1 _36494_ (.A1(_15276_),
    .A2(_15308_),
    .B1(_15314_),
    .Y(_15315_));
 sky130_fd_sc_hd__o21ai_0 _36495_ (.A1(_15309_),
    .A2(_15312_),
    .B1(_15315_),
    .Y(_15316_));
 sky130_fd_sc_hd__a21o_1 _36496_ (.A1(net601),
    .A2(_15310_),
    .B1(_15316_),
    .X(_15317_));
 sky130_fd_sc_hd__xor2_1 _36497_ (.A(_03595_),
    .B(_15317_),
    .X(_15318_));
 sky130_fd_sc_hd__nor2_1 _36498_ (.A(\inst$top.soc.cpu.multiplier.m_prod[28] ),
    .B(net2310),
    .Y(_15319_));
 sky130_fd_sc_hd__nor2_1 _36499_ (.A(net3013),
    .B(_15319_),
    .Y(_15320_));
 sky130_fd_sc_hd__o21ai_0 _36500_ (.A1(net1930),
    .A2(_15318_),
    .B1(_15320_),
    .Y(_15321_));
 sky130_fd_sc_hd__inv_2 _36501_ (.A(_15321_),
    .Y(_04373_));
 sky130_fd_sc_hd__nor2_1 _36502_ (.A(_15220_),
    .B(_15245_),
    .Y(_15322_));
 sky130_fd_sc_hd__nor2_1 _36503_ (.A(_15261_),
    .B(_15284_),
    .Y(_15323_));
 sky130_fd_sc_hd__nand2_1 _36504_ (.A(_03582_),
    .B(_03595_),
    .Y(_15324_));
 sky130_fd_sc_hd__nor2_1 _36505_ (.A(_15299_),
    .B(_15324_),
    .Y(_15325_));
 sky130_fd_sc_hd__nand2_1 _36506_ (.A(_15323_),
    .B(_15325_),
    .Y(_15326_));
 sky130_fd_sc_hd__inv_1 _36507_ (.A(_15326_),
    .Y(_15327_));
 sky130_fd_sc_hd__nand4_1 _36508_ (.A(_15159_),
    .B(_15197_),
    .C(_15322_),
    .D(_15327_),
    .Y(_15328_));
 sky130_fd_sc_hd__inv_1 _36509_ (.A(_15322_),
    .Y(_15329_));
 sky130_fd_sc_hd__a21oi_1 _36510_ (.A1(_15223_),
    .A2(_15246_),
    .B1(_15247_),
    .Y(_15330_));
 sky130_fd_sc_hd__o21ai_0 _36511_ (.A1(_15329_),
    .A2(_15201_),
    .B1(_15330_),
    .Y(_15331_));
 sky130_fd_sc_hd__nand2_1 _36512_ (.A(_15331_),
    .B(_15327_),
    .Y(_15332_));
 sky130_fd_sc_hd__o21ai_0 _36513_ (.A1(_15284_),
    .A2(_15265_),
    .B1(_15286_),
    .Y(_15333_));
 sky130_fd_sc_hd__a21oi_1 _36514_ (.A1(_03595_),
    .A2(_03581_),
    .B1(_03594_),
    .Y(_15334_));
 sky130_fd_sc_hd__o21ai_0 _36515_ (.A1(_15324_),
    .A2(_15300_),
    .B1(_15334_),
    .Y(_15335_));
 sky130_fd_sc_hd__a21oi_1 _36516_ (.A1(_15333_),
    .A2(_15325_),
    .B1(_15335_),
    .Y(_15336_));
 sky130_fd_sc_hd__nand3_1 _36517_ (.A(_15328_),
    .B(_15332_),
    .C(_15336_),
    .Y(_15337_));
 sky130_fd_sc_hd__xor2_1 _36518_ (.A(_03604_),
    .B(_15337_),
    .X(_15338_));
 sky130_fd_sc_hd__nor2_1 _36519_ (.A(\inst$top.soc.cpu.multiplier.m_prod[29] ),
    .B(net2309),
    .Y(_15339_));
 sky130_fd_sc_hd__nor2_1 _36520_ (.A(net3013),
    .B(_15339_),
    .Y(_15340_));
 sky130_fd_sc_hd__o21ai_0 _36521_ (.A1(net1930),
    .A2(_15338_),
    .B1(_15340_),
    .Y(_15341_));
 sky130_fd_sc_hd__inv_2 _36522_ (.A(_15341_),
    .Y(_04374_));
 sky130_fd_sc_hd__nor2_1 _36523_ (.A(\inst$top.soc.cpu.multiplier.x_prod[2] ),
    .B(net1922),
    .Y(_15342_));
 sky130_fd_sc_hd__o21ai_0 _36524_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[2] ),
    .A2(net2299),
    .B1(net2179),
    .Y(_15343_));
 sky130_fd_sc_hd__nor2_1 _36525_ (.A(_15342_),
    .B(_15343_),
    .Y(_04375_));
 sky130_fd_sc_hd__inv_1 _36526_ (.A(_03615_),
    .Y(_15344_));
 sky130_fd_sc_hd__a21oi_1 _36527_ (.A1(_03604_),
    .A2(_03594_),
    .B1(_03603_),
    .Y(_15345_));
 sky130_fd_sc_hd__inv_1 _36528_ (.A(_15345_),
    .Y(_15346_));
 sky130_fd_sc_hd__a31oi_1 _36529_ (.A1(_15317_),
    .A2(_03595_),
    .A3(_03604_),
    .B1(_15346_),
    .Y(_15347_));
 sky130_fd_sc_hd__inv_1 _36530_ (.A(_15347_),
    .Y(_15348_));
 sky130_fd_sc_hd__nor2_1 _36531_ (.A(_15344_),
    .B(_15348_),
    .Y(_15349_));
 sky130_fd_sc_hd__o21ai_0 _36532_ (.A1(_03615_),
    .A2(_15347_),
    .B1(net2310),
    .Y(_15350_));
 sky130_fd_sc_hd__o221ai_1 _36533_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[30] ),
    .A2(net2310),
    .B1(_15349_),
    .B2(_15350_),
    .C1(net2186),
    .Y(_15351_));
 sky130_fd_sc_hd__inv_2 _36534_ (.A(_15351_),
    .Y(_04376_));
 sky130_fd_sc_hd__inv_1 _36535_ (.A(_03627_),
    .Y(_15352_));
 sky130_fd_sc_hd__a21oi_1 _36536_ (.A1(_03615_),
    .A2(_03603_),
    .B1(_03614_),
    .Y(_15353_));
 sky130_fd_sc_hd__inv_1 _36537_ (.A(_15353_),
    .Y(_15354_));
 sky130_fd_sc_hd__a31oi_1 _36538_ (.A1(_15337_),
    .A2(_03604_),
    .A3(_03615_),
    .B1(_15354_),
    .Y(_15355_));
 sky130_fd_sc_hd__inv_1 _36539_ (.A(_15355_),
    .Y(_15356_));
 sky130_fd_sc_hd__nor2_1 _36540_ (.A(_15352_),
    .B(_15356_),
    .Y(_15357_));
 sky130_fd_sc_hd__o21ai_0 _36541_ (.A1(_03627_),
    .A2(_15355_),
    .B1(net2309),
    .Y(_15358_));
 sky130_fd_sc_hd__o221ai_1 _36542_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[31] ),
    .A2(net2310),
    .B1(_15357_),
    .B2(_15358_),
    .C1(net2186),
    .Y(_15359_));
 sky130_fd_sc_hd__inv_2 _36543_ (.A(_15359_),
    .Y(_04377_));
 sky130_fd_sc_hd__nand2_1 _36544_ (.A(_03595_),
    .B(_03604_),
    .Y(_15360_));
 sky130_fd_sc_hd__nand2_1 _36545_ (.A(_03615_),
    .B(_03627_),
    .Y(_15361_));
 sky130_fd_sc_hd__nor2_1 _36546_ (.A(_15360_),
    .B(_15361_),
    .Y(_15362_));
 sky130_fd_sc_hd__nand2_1 _36547_ (.A(_15308_),
    .B(_15362_),
    .Y(_15363_));
 sky130_fd_sc_hd__nor4_1 _36548_ (.A(_15253_),
    .B(_15273_),
    .C(_15306_),
    .D(_15363_),
    .Y(_15364_));
 sky130_fd_sc_hd__a21oi_1 _36549_ (.A1(_15238_),
    .A2(_15274_),
    .B1(_15276_),
    .Y(_15365_));
 sky130_fd_sc_hd__a21oi_1 _36550_ (.A1(_03627_),
    .A2(_03614_),
    .B1(_03626_),
    .Y(_15366_));
 sky130_fd_sc_hd__inv_1 _36551_ (.A(_15366_),
    .Y(_15367_));
 sky130_fd_sc_hd__a31oi_1 _36552_ (.A1(_15346_),
    .A2(_03615_),
    .A3(_03627_),
    .B1(_15367_),
    .Y(_15368_));
 sky130_fd_sc_hd__nand2_1 _36553_ (.A(_15314_),
    .B(_15362_),
    .Y(_15369_));
 sky130_fd_sc_hd__o211ai_1 _36554_ (.A1(_15363_),
    .A2(_15365_),
    .B1(_15368_),
    .C1(_15369_),
    .Y(_15370_));
 sky130_fd_sc_hd__a21oi_1 _36555_ (.A1(_15189_),
    .A2(_15364_),
    .B1(_15370_),
    .Y(_15371_));
 sky130_fd_sc_hd__xnor2_1 _36556_ (.A(_03635_),
    .B(_15371_),
    .Y(_15372_));
 sky130_fd_sc_hd__inv_1 _36558_ (.A(\inst$top.soc.cpu.multiplier.m_prod[32] ),
    .Y(_15374_));
 sky130_fd_sc_hd__a21oi_1 _36559_ (.A1(net1930),
    .A2(_15374_),
    .B1(net3012),
    .Y(_15375_));
 sky130_fd_sc_hd__o21ai_0 _36560_ (.A1(net1930),
    .A2(_15372_),
    .B1(_15375_),
    .Y(_15376_));
 sky130_fd_sc_hd__inv_2 _36561_ (.A(_15376_),
    .Y(_04378_));
 sky130_fd_sc_hd__nand2_1 _36562_ (.A(_03604_),
    .B(_03615_),
    .Y(_15377_));
 sky130_fd_sc_hd__nand2_1 _36563_ (.A(_03627_),
    .B(_03635_),
    .Y(_15378_));
 sky130_fd_sc_hd__nor2_1 _36564_ (.A(_15377_),
    .B(_15378_),
    .Y(_15379_));
 sky130_fd_sc_hd__a21oi_1 _36565_ (.A1(_03635_),
    .A2(_03626_),
    .B1(_03634_),
    .Y(_15380_));
 sky130_fd_sc_hd__inv_1 _36566_ (.A(_15380_),
    .Y(_15381_));
 sky130_fd_sc_hd__a31oi_1 _36567_ (.A1(_15354_),
    .A2(_03627_),
    .A3(_03635_),
    .B1(_15381_),
    .Y(_15382_));
 sky130_fd_sc_hd__inv_1 _36568_ (.A(_15382_),
    .Y(_15383_));
 sky130_fd_sc_hd__a21oi_1 _36569_ (.A1(_15337_),
    .A2(_15379_),
    .B1(_15383_),
    .Y(_15384_));
 sky130_fd_sc_hd__xnor2_1 _36570_ (.A(_03641_),
    .B(_15384_),
    .Y(_15385_));
 sky130_fd_sc_hd__inv_1 _36571_ (.A(\inst$top.soc.cpu.multiplier.m_prod[33] ),
    .Y(_15386_));
 sky130_fd_sc_hd__a21oi_1 _36573_ (.A1(net1919),
    .A2(_15386_),
    .B1(net3007),
    .Y(_15388_));
 sky130_fd_sc_hd__o21ai_0 _36574_ (.A1(net1920),
    .A2(_15385_),
    .B1(_15388_),
    .Y(_15389_));
 sky130_fd_sc_hd__inv_2 _36575_ (.A(_15389_),
    .Y(_04379_));
 sky130_fd_sc_hd__nor2_1 _36576_ (.A(_15307_),
    .B(_15360_),
    .Y(_15390_));
 sky130_fd_sc_hd__nand2_1 _36577_ (.A(_03635_),
    .B(_03641_),
    .Y(_15391_));
 sky130_fd_sc_hd__nor2_1 _36578_ (.A(_15361_),
    .B(_15391_),
    .Y(_15392_));
 sky130_fd_sc_hd__nand2_1 _36579_ (.A(_15390_),
    .B(_15392_),
    .Y(_15393_));
 sky130_fd_sc_hd__nor2_1 _36580_ (.A(_15273_),
    .B(_15292_),
    .Y(_15394_));
 sky130_fd_sc_hd__inv_1 _36581_ (.A(_15253_),
    .Y(_15395_));
 sky130_fd_sc_hd__nand3_1 _36582_ (.A(_15394_),
    .B(_15234_),
    .C(_15395_),
    .Y(_15396_));
 sky130_fd_sc_hd__nor2_1 _36583_ (.A(_15393_),
    .B(_15396_),
    .Y(_15397_));
 sky130_fd_sc_hd__o21ai_0 _36584_ (.A1(_15360_),
    .A2(_15313_),
    .B1(_15345_),
    .Y(_15398_));
 sky130_fd_sc_hd__inv_1 _36585_ (.A(_15398_),
    .Y(_15399_));
 sky130_fd_sc_hd__inv_1 _36586_ (.A(_15392_),
    .Y(_15400_));
 sky130_fd_sc_hd__a21boi_0 _36587_ (.A1(_15236_),
    .A2(_15395_),
    .B1_N(_15254_),
    .Y(_15401_));
 sky130_fd_sc_hd__inv_1 _36588_ (.A(_15401_),
    .Y(_15402_));
 sky130_fd_sc_hd__o21ai_0 _36589_ (.A1(_15292_),
    .A2(_15275_),
    .B1(_15293_),
    .Y(_15403_));
 sky130_fd_sc_hd__a21oi_1 _36590_ (.A1(_15402_),
    .A2(_15394_),
    .B1(_15403_),
    .Y(_15404_));
 sky130_fd_sc_hd__a21oi_1 _36591_ (.A1(_03641_),
    .A2(_03634_),
    .B1(_03640_),
    .Y(_15405_));
 sky130_fd_sc_hd__inv_1 _36592_ (.A(_15405_),
    .Y(_15406_));
 sky130_fd_sc_hd__a31oi_1 _36593_ (.A1(_15367_),
    .A2(_03635_),
    .A3(_03641_),
    .B1(_15406_),
    .Y(_15407_));
 sky130_fd_sc_hd__o221ai_1 _36594_ (.A1(_15399_),
    .A2(_15400_),
    .B1(_15393_),
    .B2(_15404_),
    .C1(_15407_),
    .Y(_15408_));
 sky130_fd_sc_hd__a21oi_1 _36595_ (.A1(_15215_),
    .A2(_15397_),
    .B1(_15408_),
    .Y(_15409_));
 sky130_fd_sc_hd__xnor2_1 _36596_ (.A(_03647_),
    .B(_15409_),
    .Y(_15410_));
 sky130_fd_sc_hd__inv_1 _36597_ (.A(\inst$top.soc.cpu.multiplier.m_prod[34] ),
    .Y(_15411_));
 sky130_fd_sc_hd__a21oi_1 _36598_ (.A1(net1930),
    .A2(_15411_),
    .B1(net3013),
    .Y(_15412_));
 sky130_fd_sc_hd__o21ai_0 _36599_ (.A1(net1930),
    .A2(_15410_),
    .B1(_15412_),
    .Y(_15413_));
 sky130_fd_sc_hd__inv_2 _36600_ (.A(_15413_),
    .Y(_04380_));
 sky130_fd_sc_hd__nor2_1 _36601_ (.A(_15284_),
    .B(_15299_),
    .Y(_15414_));
 sky130_fd_sc_hd__nand2_1 _36602_ (.A(_15262_),
    .B(_15414_),
    .Y(_15415_));
 sky130_fd_sc_hd__nor2_1 _36603_ (.A(_15324_),
    .B(_15377_),
    .Y(_15416_));
 sky130_fd_sc_hd__nand2_1 _36604_ (.A(_03641_),
    .B(_03647_),
    .Y(_15417_));
 sky130_fd_sc_hd__nor2_1 _36605_ (.A(_15378_),
    .B(_15417_),
    .Y(_15418_));
 sky130_fd_sc_hd__nand2_1 _36606_ (.A(_15416_),
    .B(_15418_),
    .Y(_15419_));
 sky130_fd_sc_hd__nor2_1 _36607_ (.A(_15415_),
    .B(_15419_),
    .Y(_15420_));
 sky130_fd_sc_hd__inv_1 _36608_ (.A(_15267_),
    .Y(_15421_));
 sky130_fd_sc_hd__o21ai_0 _36609_ (.A1(_15299_),
    .A2(_15286_),
    .B1(_15300_),
    .Y(_15422_));
 sky130_fd_sc_hd__a21oi_1 _36610_ (.A1(_15421_),
    .A2(_15414_),
    .B1(_15422_),
    .Y(_15423_));
 sky130_fd_sc_hd__o21ai_0 _36611_ (.A1(_15377_),
    .A2(_15334_),
    .B1(_15353_),
    .Y(_15424_));
 sky130_fd_sc_hd__a21oi_1 _36612_ (.A1(_03647_),
    .A2(_03640_),
    .B1(_03646_),
    .Y(_15425_));
 sky130_fd_sc_hd__inv_1 _36613_ (.A(_15425_),
    .Y(_15426_));
 sky130_fd_sc_hd__a31oi_1 _36614_ (.A1(_15381_),
    .A2(_03641_),
    .A3(_03647_),
    .B1(_15426_),
    .Y(_15427_));
 sky130_fd_sc_hd__inv_1 _36615_ (.A(_15427_),
    .Y(_15428_));
 sky130_fd_sc_hd__a21oi_1 _36616_ (.A1(_15424_),
    .A2(_15418_),
    .B1(_15428_),
    .Y(_15429_));
 sky130_fd_sc_hd__o21ai_0 _36617_ (.A1(_15419_),
    .A2(_15423_),
    .B1(_15429_),
    .Y(_15430_));
 sky130_fd_sc_hd__a21oi_1 _36618_ (.A1(_15225_),
    .A2(_15420_),
    .B1(_15430_),
    .Y(_15431_));
 sky130_fd_sc_hd__xnor2_2 _36619_ (.A(_03653_),
    .B(_15431_),
    .Y(_15432_));
 sky130_fd_sc_hd__inv_1 _36620_ (.A(\inst$top.soc.cpu.multiplier.m_prod[35] ),
    .Y(_15433_));
 sky130_fd_sc_hd__a21oi_1 _36621_ (.A1(net1923),
    .A2(_15433_),
    .B1(net3008),
    .Y(_15434_));
 sky130_fd_sc_hd__o21ai_0 _36622_ (.A1(net1923),
    .A2(_15432_),
    .B1(_15434_),
    .Y(_15435_));
 sky130_fd_sc_hd__inv_2 _36623_ (.A(_15435_),
    .Y(_04381_));
 sky130_fd_sc_hd__a21oi_1 _36624_ (.A1(_03653_),
    .A2(_03646_),
    .B1(_03652_),
    .Y(_15436_));
 sky130_fd_sc_hd__inv_1 _36625_ (.A(_15436_),
    .Y(_15437_));
 sky130_fd_sc_hd__nand2_1 _36626_ (.A(_03647_),
    .B(_03653_),
    .Y(_15438_));
 sky130_fd_sc_hd__nor2_1 _36627_ (.A(_15438_),
    .B(_15409_),
    .Y(_15439_));
 sky130_fd_sc_hd__nor2_1 _36628_ (.A(_15437_),
    .B(_15439_),
    .Y(_15440_));
 sky130_fd_sc_hd__xnor2_2 _36629_ (.A(_03659_),
    .B(_15440_),
    .Y(_15441_));
 sky130_fd_sc_hd__inv_1 _36630_ (.A(\inst$top.soc.cpu.multiplier.m_prod[36] ),
    .Y(_15442_));
 sky130_fd_sc_hd__a21oi_1 _36631_ (.A1(net1921),
    .A2(_15442_),
    .B1(net3008),
    .Y(_15443_));
 sky130_fd_sc_hd__o21ai_0 _36632_ (.A1(net1921),
    .A2(_15441_),
    .B1(_15443_),
    .Y(_15444_));
 sky130_fd_sc_hd__inv_2 _36633_ (.A(_15444_),
    .Y(_04382_));
 sky130_fd_sc_hd__nand2_1 _36635_ (.A(_03653_),
    .B(_03659_),
    .Y(_15446_));
 sky130_fd_sc_hd__nor2_1 _36636_ (.A(_15417_),
    .B(_15446_),
    .Y(_15447_));
 sky130_fd_sc_hd__nand2_1 _36637_ (.A(_15379_),
    .B(_15447_),
    .Y(_15448_));
 sky130_fd_sc_hd__nor2_1 _36638_ (.A(_15326_),
    .B(_15448_),
    .Y(_15449_));
 sky130_fd_sc_hd__inv_1 _36639_ (.A(_15446_),
    .Y(_15450_));
 sky130_fd_sc_hd__a21oi_1 _36640_ (.A1(_03659_),
    .A2(_03652_),
    .B1(_03658_),
    .Y(_15451_));
 sky130_fd_sc_hd__inv_1 _36641_ (.A(_15451_),
    .Y(_15452_));
 sky130_fd_sc_hd__a21oi_1 _36642_ (.A1(_15426_),
    .A2(_15450_),
    .B1(_15452_),
    .Y(_15453_));
 sky130_fd_sc_hd__a21boi_0 _36643_ (.A1(_15383_),
    .A2(_15447_),
    .B1_N(_15453_),
    .Y(_15454_));
 sky130_fd_sc_hd__o21ai_0 _36644_ (.A1(_15448_),
    .A2(_15336_),
    .B1(_15454_),
    .Y(_15455_));
 sky130_fd_sc_hd__a21oi_1 _36645_ (.A1(_15249_),
    .A2(_15449_),
    .B1(_15455_),
    .Y(_15456_));
 sky130_fd_sc_hd__xnor2_1 _36646_ (.A(_03665_),
    .B(_15456_),
    .Y(_15457_));
 sky130_fd_sc_hd__inv_1 _36647_ (.A(\inst$top.soc.cpu.multiplier.m_prod[37] ),
    .Y(_15458_));
 sky130_fd_sc_hd__a21oi_1 _36648_ (.A1(net1930),
    .A2(_15458_),
    .B1(net3013),
    .Y(_15459_));
 sky130_fd_sc_hd__o21ai_0 _36649_ (.A1(net1930),
    .A2(_15457_),
    .B1(_15459_),
    .Y(_15460_));
 sky130_fd_sc_hd__inv_2 _36650_ (.A(_15460_),
    .Y(_04383_));
 sky130_fd_sc_hd__nand2_1 _36651_ (.A(_03659_),
    .B(_03665_),
    .Y(_15461_));
 sky130_fd_sc_hd__nor2_1 _36652_ (.A(_15438_),
    .B(_15461_),
    .Y(_15462_));
 sky130_fd_sc_hd__inv_1 _36653_ (.A(_15462_),
    .Y(_15463_));
 sky130_fd_sc_hd__a21oi_1 _36654_ (.A1(_03665_),
    .A2(_03658_),
    .B1(_03664_),
    .Y(_15464_));
 sky130_fd_sc_hd__inv_1 _36655_ (.A(_15464_),
    .Y(_15465_));
 sky130_fd_sc_hd__a31oi_1 _36656_ (.A1(_15437_),
    .A2(_03659_),
    .A3(_03665_),
    .B1(_15465_),
    .Y(_15466_));
 sky130_fd_sc_hd__o21ai_0 _36657_ (.A1(_15463_),
    .A2(_15409_),
    .B1(_15466_),
    .Y(_15467_));
 sky130_fd_sc_hd__xor2_1 _36658_ (.A(_03671_),
    .B(_15467_),
    .X(_15468_));
 sky130_fd_sc_hd__inv_1 _36659_ (.A(\inst$top.soc.cpu.multiplier.m_prod[38] ),
    .Y(_15469_));
 sky130_fd_sc_hd__a21oi_1 _36660_ (.A1(net1919),
    .A2(_15469_),
    .B1(net3007),
    .Y(_15470_));
 sky130_fd_sc_hd__o21ai_0 _36661_ (.A1(net1919),
    .A2(_15468_),
    .B1(_15470_),
    .Y(_15471_));
 sky130_fd_sc_hd__inv_2 _36662_ (.A(_15471_),
    .Y(_04384_));
 sky130_fd_sc_hd__nand2_1 _36663_ (.A(_03665_),
    .B(_03671_),
    .Y(_15472_));
 sky130_fd_sc_hd__nor2_1 _36664_ (.A(_15446_),
    .B(_15472_),
    .Y(_15473_));
 sky130_fd_sc_hd__inv_1 _36665_ (.A(_15473_),
    .Y(_15474_));
 sky130_fd_sc_hd__inv_1 _36666_ (.A(_15472_),
    .Y(_15475_));
 sky130_fd_sc_hd__a21oi_1 _36667_ (.A1(_03671_),
    .A2(_03664_),
    .B1(_03670_),
    .Y(_15476_));
 sky130_fd_sc_hd__inv_1 _36668_ (.A(_15476_),
    .Y(_15477_));
 sky130_fd_sc_hd__a21oi_1 _36669_ (.A1(_15452_),
    .A2(_15475_),
    .B1(_15477_),
    .Y(_15478_));
 sky130_fd_sc_hd__o21ai_0 _36670_ (.A1(_15474_),
    .A2(_15431_),
    .B1(_15478_),
    .Y(_15479_));
 sky130_fd_sc_hd__xor2_1 _36671_ (.A(_02554_),
    .B(_15479_),
    .X(_15480_));
 sky130_fd_sc_hd__inv_1 _36672_ (.A(\inst$top.soc.cpu.multiplier.m_prod[39] ),
    .Y(_15481_));
 sky130_fd_sc_hd__a21oi_1 _36673_ (.A1(net1921),
    .A2(_15481_),
    .B1(net3007),
    .Y(_15482_));
 sky130_fd_sc_hd__o21ai_0 _36674_ (.A1(net1921),
    .A2(_15480_),
    .B1(_15482_),
    .Y(_15483_));
 sky130_fd_sc_hd__inv_2 _36675_ (.A(_15483_),
    .Y(_04385_));
 sky130_fd_sc_hd__nor2_1 _36676_ (.A(\inst$top.soc.cpu.multiplier.x_prod[3] ),
    .B(net1922),
    .Y(_15484_));
 sky130_fd_sc_hd__o21ai_0 _36677_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[3] ),
    .A2(net2299),
    .B1(net2179),
    .Y(_15485_));
 sky130_fd_sc_hd__nor2_1 _36678_ (.A(_15484_),
    .B(_15485_),
    .Y(_04386_));
 sky130_fd_sc_hd__nand2_1 _36679_ (.A(_02554_),
    .B(_03671_),
    .Y(_15486_));
 sky130_fd_sc_hd__nor2_1 _36680_ (.A(_15461_),
    .B(_15486_),
    .Y(_15487_));
 sky130_fd_sc_hd__inv_1 _36681_ (.A(_15487_),
    .Y(_15488_));
 sky130_fd_sc_hd__a21oi_1 _36682_ (.A1(_02554_),
    .A2(_03670_),
    .B1(_02553_),
    .Y(_15489_));
 sky130_fd_sc_hd__inv_1 _36683_ (.A(_15489_),
    .Y(_15490_));
 sky130_fd_sc_hd__a31oi_1 _36684_ (.A1(_15465_),
    .A2(_02554_),
    .A3(_03671_),
    .B1(_15490_),
    .Y(_15491_));
 sky130_fd_sc_hd__o21ai_0 _36685_ (.A1(_15488_),
    .A2(_15440_),
    .B1(_15491_),
    .Y(_15492_));
 sky130_fd_sc_hd__xor2_1 _36686_ (.A(_02560_),
    .B(_15492_),
    .X(_15493_));
 sky130_fd_sc_hd__inv_1 _36688_ (.A(\inst$top.soc.cpu.multiplier.m_prod[40] ),
    .Y(_15495_));
 sky130_fd_sc_hd__a21oi_1 _36689_ (.A1(net1928),
    .A2(_15495_),
    .B1(net3012),
    .Y(_15496_));
 sky130_fd_sc_hd__o21ai_0 _36690_ (.A1(net1928),
    .A2(_15493_),
    .B1(_15496_),
    .Y(_15497_));
 sky130_fd_sc_hd__inv_2 _36691_ (.A(_15497_),
    .Y(_04387_));
 sky130_fd_sc_hd__nand2_1 _36692_ (.A(_02554_),
    .B(_02560_),
    .Y(_15498_));
 sky130_fd_sc_hd__nor2_1 _36693_ (.A(_15472_),
    .B(_15498_),
    .Y(_15499_));
 sky130_fd_sc_hd__inv_1 _36694_ (.A(_15499_),
    .Y(_15500_));
 sky130_fd_sc_hd__a21oi_1 _36695_ (.A1(_02560_),
    .A2(_02553_),
    .B1(_02559_),
    .Y(_15501_));
 sky130_fd_sc_hd__inv_1 _36696_ (.A(_15501_),
    .Y(_15502_));
 sky130_fd_sc_hd__a31oi_1 _36697_ (.A1(_15477_),
    .A2(_02554_),
    .A3(_02560_),
    .B1(_15502_),
    .Y(_15503_));
 sky130_fd_sc_hd__o21ai_0 _36698_ (.A1(_15500_),
    .A2(_15456_),
    .B1(_15503_),
    .Y(_15504_));
 sky130_fd_sc_hd__xor2_1 _36699_ (.A(_02566_),
    .B(_15504_),
    .X(_15505_));
 sky130_fd_sc_hd__inv_1 _36700_ (.A(\inst$top.soc.cpu.multiplier.m_prod[41] ),
    .Y(_15506_));
 sky130_fd_sc_hd__a21oi_1 _36701_ (.A1(net1928),
    .A2(_15506_),
    .B1(net3012),
    .Y(_15507_));
 sky130_fd_sc_hd__o21ai_0 _36702_ (.A1(net1928),
    .A2(_15505_),
    .B1(_15507_),
    .Y(_15508_));
 sky130_fd_sc_hd__inv_2 _36703_ (.A(_15508_),
    .Y(_04388_));
 sky130_fd_sc_hd__nand2_1 _36704_ (.A(_02560_),
    .B(_02566_),
    .Y(_15509_));
 sky130_fd_sc_hd__nor2_1 _36705_ (.A(_15486_),
    .B(_15509_),
    .Y(_15510_));
 sky130_fd_sc_hd__nand2_1 _36706_ (.A(_15467_),
    .B(_15510_),
    .Y(_15511_));
 sky130_fd_sc_hd__a21oi_1 _36707_ (.A1(_02566_),
    .A2(_02559_),
    .B1(_02565_),
    .Y(_15512_));
 sky130_fd_sc_hd__inv_1 _36708_ (.A(_15512_),
    .Y(_15513_));
 sky130_fd_sc_hd__a31oi_1 _36709_ (.A1(_15490_),
    .A2(_02560_),
    .A3(_02566_),
    .B1(_15513_),
    .Y(_15514_));
 sky130_fd_sc_hd__nand2_1 _36710_ (.A(_15511_),
    .B(_15514_),
    .Y(_15515_));
 sky130_fd_sc_hd__xor2_1 _36711_ (.A(_02572_),
    .B(_15515_),
    .X(_15516_));
 sky130_fd_sc_hd__inv_1 _36712_ (.A(\inst$top.soc.cpu.multiplier.m_prod[42] ),
    .Y(_15517_));
 sky130_fd_sc_hd__a21oi_1 _36713_ (.A1(net1919),
    .A2(_15517_),
    .B1(net3007),
    .Y(_15518_));
 sky130_fd_sc_hd__o21ai_0 _36714_ (.A1(net1919),
    .A2(_15516_),
    .B1(_15518_),
    .Y(_15519_));
 sky130_fd_sc_hd__inv_2 _36715_ (.A(_15519_),
    .Y(_04389_));
 sky130_fd_sc_hd__nand2_1 _36716_ (.A(_02566_),
    .B(_02572_),
    .Y(_15520_));
 sky130_fd_sc_hd__nor2_1 _36717_ (.A(_15498_),
    .B(_15520_),
    .Y(_15521_));
 sky130_fd_sc_hd__inv_1 _36718_ (.A(_15520_),
    .Y(_15522_));
 sky130_fd_sc_hd__a21oi_1 _36719_ (.A1(_02572_),
    .A2(_02565_),
    .B1(_02571_),
    .Y(_15523_));
 sky130_fd_sc_hd__inv_1 _36720_ (.A(_15523_),
    .Y(_15524_));
 sky130_fd_sc_hd__a21oi_1 _36721_ (.A1(_15502_),
    .A2(_15522_),
    .B1(_15524_),
    .Y(_15525_));
 sky130_fd_sc_hd__a21boi_0 _36722_ (.A1(_15479_),
    .A2(_15521_),
    .B1_N(_15525_),
    .Y(_15526_));
 sky130_fd_sc_hd__or2_2 _36723_ (.A(_02578_),
    .B(_15526_),
    .X(_15527_));
 sky130_fd_sc_hd__nand2_1 _36725_ (.A(_15526_),
    .B(_02578_),
    .Y(_15529_));
 sky130_fd_sc_hd__nand3_1 _36726_ (.A(_15527_),
    .B(net2310),
    .C(_15529_),
    .Y(_15530_));
 sky130_fd_sc_hd__o211ai_1 _36727_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[43] ),
    .A2(net2300),
    .B1(net2179),
    .C1(_15530_),
    .Y(_15531_));
 sky130_fd_sc_hd__inv_2 _36728_ (.A(_15531_),
    .Y(_04390_));
 sky130_fd_sc_hd__inv_1 _36729_ (.A(_15438_),
    .Y(_15532_));
 sky130_fd_sc_hd__a21oi_1 _36730_ (.A1(_15406_),
    .A2(_15532_),
    .B1(_15437_),
    .Y(_15533_));
 sky130_fd_sc_hd__o31ai_1 _36731_ (.A1(_15391_),
    .A2(_15438_),
    .A3(_15368_),
    .B1(_15533_),
    .Y(_15534_));
 sky130_fd_sc_hd__nand2_1 _36732_ (.A(_02572_),
    .B(_02578_),
    .Y(_15535_));
 sky130_fd_sc_hd__nor2_1 _36733_ (.A(_15509_),
    .B(_15535_),
    .Y(_15536_));
 sky130_fd_sc_hd__inv_1 _36734_ (.A(_15536_),
    .Y(_15537_));
 sky130_fd_sc_hd__nor2_1 _36735_ (.A(_15488_),
    .B(_15537_),
    .Y(_15538_));
 sky130_fd_sc_hd__a21oi_1 _36736_ (.A1(_02578_),
    .A2(_02571_),
    .B1(_02577_),
    .Y(_15539_));
 sky130_fd_sc_hd__inv_1 _36737_ (.A(_15539_),
    .Y(_15540_));
 sky130_fd_sc_hd__a31oi_1 _36738_ (.A1(_15513_),
    .A2(_02572_),
    .A3(_02578_),
    .B1(_15540_),
    .Y(_15541_));
 sky130_fd_sc_hd__o21ai_0 _36739_ (.A1(_15537_),
    .A2(_15491_),
    .B1(_15541_),
    .Y(_15542_));
 sky130_fd_sc_hd__a21oi_1 _36740_ (.A1(_15534_),
    .A2(_15538_),
    .B1(_15542_),
    .Y(_15543_));
 sky130_fd_sc_hd__nor2_1 _36741_ (.A(_15391_),
    .B(_15438_),
    .Y(_15544_));
 sky130_fd_sc_hd__and3_1 _36742_ (.A(_15538_),
    .B(_15362_),
    .C(_15544_),
    .X(_15545_));
 sky130_fd_sc_hd__nand2_1 _36743_ (.A(_15316_),
    .B(_15545_),
    .Y(_15546_));
 sky130_fd_sc_hd__nand3_1 _36744_ (.A(net601),
    .B(_15310_),
    .C(_15545_),
    .Y(_15547_));
 sky130_fd_sc_hd__nand3_1 _36745_ (.A(_15543_),
    .B(_15546_),
    .C(_15547_),
    .Y(_15548_));
 sky130_fd_sc_hd__xor2_1 _36746_ (.A(_02584_),
    .B(_15548_),
    .X(_15549_));
 sky130_fd_sc_hd__inv_1 _36747_ (.A(\inst$top.soc.cpu.multiplier.m_prod[44] ),
    .Y(_15550_));
 sky130_fd_sc_hd__a21oi_1 _36749_ (.A1(net1928),
    .A2(_15550_),
    .B1(net3012),
    .Y(_15552_));
 sky130_fd_sc_hd__o21ai_0 _36750_ (.A1(net1928),
    .A2(_15549_),
    .B1(_15552_),
    .Y(_15553_));
 sky130_fd_sc_hd__inv_2 _36751_ (.A(_15553_),
    .Y(_04391_));
 sky130_fd_sc_hd__nand2_1 _36752_ (.A(_02578_),
    .B(_02584_),
    .Y(_15554_));
 sky130_fd_sc_hd__nor2_1 _36753_ (.A(_15520_),
    .B(_15554_),
    .Y(_15555_));
 sky130_fd_sc_hd__nand2_1 _36754_ (.A(_15504_),
    .B(_15555_),
    .Y(_15556_));
 sky130_fd_sc_hd__a21oi_1 _36755_ (.A1(_02584_),
    .A2(_02577_),
    .B1(_02583_),
    .Y(_15557_));
 sky130_fd_sc_hd__inv_1 _36756_ (.A(_15557_),
    .Y(_15558_));
 sky130_fd_sc_hd__a31oi_1 _36757_ (.A1(_15524_),
    .A2(_02578_),
    .A3(_02584_),
    .B1(_15558_),
    .Y(_15559_));
 sky130_fd_sc_hd__nand2_1 _36758_ (.A(_15556_),
    .B(_15559_),
    .Y(_15560_));
 sky130_fd_sc_hd__xor2_1 _36759_ (.A(_02590_),
    .B(_15560_),
    .X(_15561_));
 sky130_fd_sc_hd__inv_1 _36760_ (.A(\inst$top.soc.cpu.multiplier.m_prod[45] ),
    .Y(_15562_));
 sky130_fd_sc_hd__a21oi_1 _36761_ (.A1(net1920),
    .A2(_15562_),
    .B1(net3008),
    .Y(_15563_));
 sky130_fd_sc_hd__o21ai_0 _36762_ (.A1(net1919),
    .A2(_15561_),
    .B1(_15563_),
    .Y(_15564_));
 sky130_fd_sc_hd__inv_2 _36763_ (.A(_15564_),
    .Y(_04392_));
 sky130_fd_sc_hd__inv_1 _36764_ (.A(_15510_),
    .Y(_15565_));
 sky130_fd_sc_hd__nand2_1 _36765_ (.A(_02584_),
    .B(_02590_),
    .Y(_15566_));
 sky130_fd_sc_hd__nor2_1 _36766_ (.A(_15535_),
    .B(_15566_),
    .Y(_15567_));
 sky130_fd_sc_hd__inv_1 _36767_ (.A(_15567_),
    .Y(_15568_));
 sky130_fd_sc_hd__nor2_1 _36768_ (.A(_15565_),
    .B(_15568_),
    .Y(_15569_));
 sky130_fd_sc_hd__a21oi_1 _36769_ (.A1(_02590_),
    .A2(_02583_),
    .B1(_02589_),
    .Y(_15570_));
 sky130_fd_sc_hd__inv_1 _36770_ (.A(_15570_),
    .Y(_15571_));
 sky130_fd_sc_hd__a31oi_1 _36771_ (.A1(_15540_),
    .A2(_02584_),
    .A3(_02590_),
    .B1(_15571_),
    .Y(_15572_));
 sky130_fd_sc_hd__o21ai_0 _36772_ (.A1(_15568_),
    .A2(_15514_),
    .B1(_15572_),
    .Y(_15573_));
 sky130_fd_sc_hd__a21oi_1 _36773_ (.A1(_15467_),
    .A2(_15569_),
    .B1(_15573_),
    .Y(_15574_));
 sky130_fd_sc_hd__or2_2 _36774_ (.A(_02596_),
    .B(_15574_),
    .X(_15575_));
 sky130_fd_sc_hd__nand2_1 _36775_ (.A(_15574_),
    .B(_02596_),
    .Y(_15576_));
 sky130_fd_sc_hd__nand3_1 _36776_ (.A(_15575_),
    .B(net2310),
    .C(_15576_),
    .Y(_15577_));
 sky130_fd_sc_hd__o211ai_1 _36777_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[46] ),
    .A2(net2305),
    .B1(net2179),
    .C1(_15577_),
    .Y(_15578_));
 sky130_fd_sc_hd__inv_2 _36778_ (.A(_15578_),
    .Y(_04393_));
 sky130_fd_sc_hd__inv_1 _36779_ (.A(_15521_),
    .Y(_15579_));
 sky130_fd_sc_hd__nand2_1 _36780_ (.A(_02590_),
    .B(_02596_),
    .Y(_15580_));
 sky130_fd_sc_hd__nor2_1 _36781_ (.A(_15554_),
    .B(_15580_),
    .Y(_15581_));
 sky130_fd_sc_hd__inv_1 _36782_ (.A(_15581_),
    .Y(_15582_));
 sky130_fd_sc_hd__nor2_1 _36783_ (.A(_15579_),
    .B(_15582_),
    .Y(_15583_));
 sky130_fd_sc_hd__nand2_1 _36784_ (.A(_15479_),
    .B(_15583_),
    .Y(_15584_));
 sky130_fd_sc_hd__a21oi_1 _36785_ (.A1(_02596_),
    .A2(_02589_),
    .B1(_02595_),
    .Y(_15585_));
 sky130_fd_sc_hd__inv_1 _36786_ (.A(_15585_),
    .Y(_15586_));
 sky130_fd_sc_hd__a31oi_1 _36787_ (.A1(_15558_),
    .A2(_02590_),
    .A3(_02596_),
    .B1(_15586_),
    .Y(_15587_));
 sky130_fd_sc_hd__o21ai_0 _36788_ (.A1(_15582_),
    .A2(_15525_),
    .B1(_15587_),
    .Y(_15588_));
 sky130_fd_sc_hd__inv_1 _36789_ (.A(_15588_),
    .Y(_15589_));
 sky130_fd_sc_hd__nand2_1 _36790_ (.A(_15584_),
    .B(_15589_),
    .Y(_15590_));
 sky130_fd_sc_hd__xor2_1 _36791_ (.A(_02602_),
    .B(_15590_),
    .X(_15591_));
 sky130_fd_sc_hd__inv_1 _36792_ (.A(\inst$top.soc.cpu.multiplier.m_prod[47] ),
    .Y(_15592_));
 sky130_fd_sc_hd__a21oi_1 _36793_ (.A1(net1919),
    .A2(_15592_),
    .B1(net3008),
    .Y(_15593_));
 sky130_fd_sc_hd__o21ai_0 _36794_ (.A1(net1919),
    .A2(_15591_),
    .B1(_15593_),
    .Y(_15594_));
 sky130_fd_sc_hd__inv_2 _36795_ (.A(_15594_),
    .Y(_04394_));
 sky130_fd_sc_hd__nand2_1 _36796_ (.A(_02596_),
    .B(_02602_),
    .Y(_15595_));
 sky130_fd_sc_hd__nor2_1 _36797_ (.A(_15566_),
    .B(_15595_),
    .Y(_15596_));
 sky130_fd_sc_hd__inv_1 _36798_ (.A(_15596_),
    .Y(_15597_));
 sky130_fd_sc_hd__nor2_1 _36799_ (.A(_15537_),
    .B(_15597_),
    .Y(_15598_));
 sky130_fd_sc_hd__and3_1 _36800_ (.A(_15598_),
    .B(_15544_),
    .C(_15487_),
    .X(_15599_));
 sky130_fd_sc_hd__nand2_1 _36801_ (.A(_15370_),
    .B(_15599_),
    .Y(_15600_));
 sky130_fd_sc_hd__o21ai_0 _36802_ (.A1(_15488_),
    .A2(_15533_),
    .B1(_15491_),
    .Y(_15601_));
 sky130_fd_sc_hd__a21oi_1 _36803_ (.A1(_02602_),
    .A2(_02595_),
    .B1(_02601_),
    .Y(_15602_));
 sky130_fd_sc_hd__inv_1 _36804_ (.A(_15602_),
    .Y(_15603_));
 sky130_fd_sc_hd__a31oi_1 _36805_ (.A1(_15571_),
    .A2(_02596_),
    .A3(_02602_),
    .B1(_15603_),
    .Y(_15604_));
 sky130_fd_sc_hd__o21ai_0 _36806_ (.A1(_15597_),
    .A2(_15541_),
    .B1(_15604_),
    .Y(_15605_));
 sky130_fd_sc_hd__a21oi_1 _36807_ (.A1(_15601_),
    .A2(_15598_),
    .B1(_15605_),
    .Y(_15606_));
 sky130_fd_sc_hd__nand3_1 _36808_ (.A(_15189_),
    .B(_15364_),
    .C(_15599_),
    .Y(_15607_));
 sky130_fd_sc_hd__nand3_1 _36809_ (.A(_15600_),
    .B(_15606_),
    .C(_15607_),
    .Y(_15608_));
 sky130_fd_sc_hd__nor2_1 _36810_ (.A(_02609_),
    .B(_15608_),
    .Y(_15609_));
 sky130_fd_sc_hd__nand2_1 _36811_ (.A(_15608_),
    .B(_02609_),
    .Y(_15610_));
 sky130_fd_sc_hd__inv_1 _36812_ (.A(_15610_),
    .Y(_15611_));
 sky130_fd_sc_hd__o21ai_0 _36813_ (.A1(_15609_),
    .A2(_15611_),
    .B1(net2308),
    .Y(_15612_));
 sky130_fd_sc_hd__o211ai_1 _36814_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[48] ),
    .A2(net2305),
    .B1(net2184),
    .C1(_15612_),
    .Y(_15613_));
 sky130_fd_sc_hd__inv_2 _36815_ (.A(_15613_),
    .Y(_04395_));
 sky130_fd_sc_hd__inv_1 _36816_ (.A(_15555_),
    .Y(_15614_));
 sky130_fd_sc_hd__nand2_1 _36817_ (.A(_02602_),
    .B(_02609_),
    .Y(_15615_));
 sky130_fd_sc_hd__nor2_1 _36818_ (.A(_15580_),
    .B(_15615_),
    .Y(_15616_));
 sky130_fd_sc_hd__inv_1 _36819_ (.A(_15616_),
    .Y(_15617_));
 sky130_fd_sc_hd__nor2_1 _36820_ (.A(_15614_),
    .B(_15617_),
    .Y(_15618_));
 sky130_fd_sc_hd__nand2_1 _36821_ (.A(_15504_),
    .B(_15618_),
    .Y(_15619_));
 sky130_fd_sc_hd__a21oi_1 _36822_ (.A1(_02609_),
    .A2(_02601_),
    .B1(_02608_),
    .Y(_15620_));
 sky130_fd_sc_hd__inv_1 _36823_ (.A(_15620_),
    .Y(_15621_));
 sky130_fd_sc_hd__a31oi_1 _36824_ (.A1(_15586_),
    .A2(_02602_),
    .A3(_02609_),
    .B1(_15621_),
    .Y(_15622_));
 sky130_fd_sc_hd__o21ai_0 _36825_ (.A1(_15617_),
    .A2(_15559_),
    .B1(_15622_),
    .Y(_15623_));
 sky130_fd_sc_hd__inv_1 _36826_ (.A(_15623_),
    .Y(_15624_));
 sky130_fd_sc_hd__nand2_1 _36827_ (.A(_15619_),
    .B(_15624_),
    .Y(_15625_));
 sky130_fd_sc_hd__xor2_1 _36828_ (.A(_02615_),
    .B(_15625_),
    .X(_15626_));
 sky130_fd_sc_hd__inv_1 _36829_ (.A(\inst$top.soc.cpu.multiplier.m_prod[49] ),
    .Y(_15627_));
 sky130_fd_sc_hd__a21oi_1 _36830_ (.A1(net1931),
    .A2(_15627_),
    .B1(net3013),
    .Y(_15628_));
 sky130_fd_sc_hd__o21ai_0 _36831_ (.A1(net1931),
    .A2(_15626_),
    .B1(_15628_),
    .Y(_15629_));
 sky130_fd_sc_hd__inv_2 _36832_ (.A(_15629_),
    .Y(_04396_));
 sky130_fd_sc_hd__nor2_1 _36833_ (.A(\inst$top.soc.cpu.multiplier.x_prod[4] ),
    .B(net1922),
    .Y(_15630_));
 sky130_fd_sc_hd__o21ai_0 _36836_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[4] ),
    .A2(net2299),
    .B1(net2179),
    .Y(_15633_));
 sky130_fd_sc_hd__nor2_1 _36837_ (.A(_15630_),
    .B(_15633_),
    .Y(_04397_));
 sky130_fd_sc_hd__nand2_1 _36839_ (.A(_02609_),
    .B(_02615_),
    .Y(_15635_));
 sky130_fd_sc_hd__nor2_1 _36840_ (.A(_15595_),
    .B(_15635_),
    .Y(_15636_));
 sky130_fd_sc_hd__inv_1 _36841_ (.A(_15636_),
    .Y(_15637_));
 sky130_fd_sc_hd__nor4_1 _36842_ (.A(_15463_),
    .B(_15565_),
    .C(_15568_),
    .D(_15637_),
    .Y(_15638_));
 sky130_fd_sc_hd__nand3_1 _36843_ (.A(_15215_),
    .B(_15397_),
    .C(_15638_),
    .Y(_15639_));
 sky130_fd_sc_hd__o21ai_0 _36844_ (.A1(_15565_),
    .A2(_15466_),
    .B1(_15514_),
    .Y(_15640_));
 sky130_fd_sc_hd__nor2_1 _36845_ (.A(_15568_),
    .B(_15637_),
    .Y(_15641_));
 sky130_fd_sc_hd__inv_1 _36846_ (.A(_15635_),
    .Y(_15642_));
 sky130_fd_sc_hd__a21oi_1 _36847_ (.A1(_02615_),
    .A2(_02608_),
    .B1(_02614_),
    .Y(_15643_));
 sky130_fd_sc_hd__inv_1 _36848_ (.A(_15643_),
    .Y(_15644_));
 sky130_fd_sc_hd__a21oi_1 _36849_ (.A1(_15603_),
    .A2(_15642_),
    .B1(_15644_),
    .Y(_15645_));
 sky130_fd_sc_hd__o21ai_0 _36850_ (.A1(_15637_),
    .A2(_15572_),
    .B1(_15645_),
    .Y(_15646_));
 sky130_fd_sc_hd__a21oi_1 _36851_ (.A1(_15640_),
    .A2(_15641_),
    .B1(_15646_),
    .Y(_15647_));
 sky130_fd_sc_hd__nand2_1 _36852_ (.A(_15408_),
    .B(_15638_),
    .Y(_15648_));
 sky130_fd_sc_hd__nand3_1 _36853_ (.A(_15639_),
    .B(_15647_),
    .C(_15648_),
    .Y(_15649_));
 sky130_fd_sc_hd__xor2_1 _36854_ (.A(_02622_),
    .B(_15649_),
    .X(_15650_));
 sky130_fd_sc_hd__inv_1 _36855_ (.A(\inst$top.soc.cpu.multiplier.m_prod[50] ),
    .Y(_15651_));
 sky130_fd_sc_hd__a21oi_1 _36856_ (.A1(net1920),
    .A2(_15651_),
    .B1(net3007),
    .Y(_15652_));
 sky130_fd_sc_hd__o21ai_0 _36857_ (.A1(net1920),
    .A2(_15650_),
    .B1(_15652_),
    .Y(_15653_));
 sky130_fd_sc_hd__inv_2 _36858_ (.A(_15653_),
    .Y(_04398_));
 sky130_fd_sc_hd__nand2_1 _36859_ (.A(_02615_),
    .B(_02622_),
    .Y(_15654_));
 sky130_fd_sc_hd__nor2_1 _36860_ (.A(_15615_),
    .B(_15654_),
    .Y(_15655_));
 sky130_fd_sc_hd__inv_1 _36861_ (.A(_15655_),
    .Y(_15656_));
 sky130_fd_sc_hd__nor4_1 _36862_ (.A(_15474_),
    .B(_15579_),
    .C(_15582_),
    .D(_15656_),
    .Y(_15657_));
 sky130_fd_sc_hd__nand3_1 _36863_ (.A(_15225_),
    .B(_15420_),
    .C(_15657_),
    .Y(_15658_));
 sky130_fd_sc_hd__o21ai_0 _36864_ (.A1(_15579_),
    .A2(_15478_),
    .B1(_15525_),
    .Y(_15659_));
 sky130_fd_sc_hd__nor2_1 _36865_ (.A(_15582_),
    .B(_15656_),
    .Y(_15660_));
 sky130_fd_sc_hd__nand2_1 _36866_ (.A(_02622_),
    .B(_02614_),
    .Y(_15661_));
 sky130_fd_sc_hd__inv_1 _36867_ (.A(_02621_),
    .Y(_15662_));
 sky130_fd_sc_hd__nand2_1 _36868_ (.A(_15661_),
    .B(_15662_),
    .Y(_15663_));
 sky130_fd_sc_hd__a31oi_1 _36869_ (.A1(_15621_),
    .A2(_02615_),
    .A3(_02622_),
    .B1(_15663_),
    .Y(_15664_));
 sky130_fd_sc_hd__o21ai_0 _36870_ (.A1(_15656_),
    .A2(_15587_),
    .B1(_15664_),
    .Y(_15665_));
 sky130_fd_sc_hd__a21oi_1 _36871_ (.A1(_15659_),
    .A2(_15660_),
    .B1(_15665_),
    .Y(_15666_));
 sky130_fd_sc_hd__nand2_1 _36872_ (.A(_15430_),
    .B(_15657_),
    .Y(_15667_));
 sky130_fd_sc_hd__nand3_1 _36873_ (.A(_15658_),
    .B(_15666_),
    .C(_15667_),
    .Y(_15668_));
 sky130_fd_sc_hd__nor2_1 _36874_ (.A(_02628_),
    .B(_15668_),
    .Y(_15669_));
 sky130_fd_sc_hd__nand2_1 _36875_ (.A(_15668_),
    .B(_02628_),
    .Y(_15670_));
 sky130_fd_sc_hd__inv_1 _36876_ (.A(_15670_),
    .Y(_15671_));
 sky130_fd_sc_hd__o21ai_0 _36877_ (.A1(_15669_),
    .A2(_15671_),
    .B1(net2308),
    .Y(_15672_));
 sky130_fd_sc_hd__o211ai_1 _36878_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[51] ),
    .A2(net2305),
    .B1(net2184),
    .C1(_15672_),
    .Y(_15673_));
 sky130_fd_sc_hd__inv_2 _36879_ (.A(_15673_),
    .Y(_04399_));
 sky130_fd_sc_hd__nand2_1 _36880_ (.A(_02622_),
    .B(_02628_),
    .Y(_15674_));
 sky130_fd_sc_hd__inv_1 _36881_ (.A(_15674_),
    .Y(_15675_));
 sky130_fd_sc_hd__nand2_1 _36882_ (.A(_15642_),
    .B(_15675_),
    .Y(_15676_));
 sky130_fd_sc_hd__nor2_1 _36883_ (.A(_15676_),
    .B(_15597_),
    .Y(_15677_));
 sky130_fd_sc_hd__a21oi_1 _36884_ (.A1(_02628_),
    .A2(_02621_),
    .B1(_02627_),
    .Y(_15678_));
 sky130_fd_sc_hd__inv_1 _36885_ (.A(_15678_),
    .Y(_15679_));
 sky130_fd_sc_hd__a21oi_1 _36886_ (.A1(_15644_),
    .A2(_15675_),
    .B1(_15679_),
    .Y(_15680_));
 sky130_fd_sc_hd__o21ai_0 _36887_ (.A1(_15676_),
    .A2(_15604_),
    .B1(_15680_),
    .Y(_15681_));
 sky130_fd_sc_hd__a21o_1 _36888_ (.A1(_15548_),
    .A2(_15677_),
    .B1(_15681_),
    .X(_15682_));
 sky130_fd_sc_hd__xor2_1 _36889_ (.A(_02634_),
    .B(_15682_),
    .X(_15683_));
 sky130_fd_sc_hd__inv_1 _36890_ (.A(\inst$top.soc.cpu.multiplier.m_prod[52] ),
    .Y(_15684_));
 sky130_fd_sc_hd__a21oi_1 _36891_ (.A1(net1929),
    .A2(_15684_),
    .B1(net3012),
    .Y(_15685_));
 sky130_fd_sc_hd__o21ai_0 _36892_ (.A1(net1929),
    .A2(_15683_),
    .B1(_15685_),
    .Y(_15686_));
 sky130_fd_sc_hd__inv_2 _36893_ (.A(_15686_),
    .Y(_04400_));
 sky130_fd_sc_hd__nand2_1 _36894_ (.A(_02628_),
    .B(_02634_),
    .Y(_15687_));
 sky130_fd_sc_hd__nor2_1 _36895_ (.A(_15654_),
    .B(_15687_),
    .Y(_15688_));
 sky130_fd_sc_hd__inv_1 _36896_ (.A(_15688_),
    .Y(_15689_));
 sky130_fd_sc_hd__nor2_1 _36897_ (.A(_15500_),
    .B(_15614_),
    .Y(_15690_));
 sky130_fd_sc_hd__inv_1 _36898_ (.A(_15690_),
    .Y(_15691_));
 sky130_fd_sc_hd__nor3_1 _36899_ (.A(_15617_),
    .B(_15689_),
    .C(_15691_),
    .Y(_15692_));
 sky130_fd_sc_hd__nand3_1 _36900_ (.A(_15249_),
    .B(_15449_),
    .C(_15692_),
    .Y(_15693_));
 sky130_fd_sc_hd__o21ai_0 _36901_ (.A1(_15614_),
    .A2(_15503_),
    .B1(_15559_),
    .Y(_15694_));
 sky130_fd_sc_hd__nor2_1 _36902_ (.A(_15617_),
    .B(_15689_),
    .Y(_15695_));
 sky130_fd_sc_hd__nand2_1 _36903_ (.A(_02634_),
    .B(_02627_),
    .Y(_15696_));
 sky130_fd_sc_hd__inv_1 _36904_ (.A(_02633_),
    .Y(_15697_));
 sky130_fd_sc_hd__nand2_1 _36905_ (.A(_15696_),
    .B(_15697_),
    .Y(_15698_));
 sky130_fd_sc_hd__a31oi_1 _36906_ (.A1(_15663_),
    .A2(_02628_),
    .A3(_02634_),
    .B1(_15698_),
    .Y(_15699_));
 sky130_fd_sc_hd__o21ai_0 _36907_ (.A1(_15689_),
    .A2(_15622_),
    .B1(_15699_),
    .Y(_15700_));
 sky130_fd_sc_hd__a21oi_1 _36908_ (.A1(_15694_),
    .A2(_15695_),
    .B1(_15700_),
    .Y(_15701_));
 sky130_fd_sc_hd__nand2_1 _36909_ (.A(_15455_),
    .B(_15692_),
    .Y(_15702_));
 sky130_fd_sc_hd__nand3_1 _36910_ (.A(_15693_),
    .B(_15701_),
    .C(_15702_),
    .Y(_15703_));
 sky130_fd_sc_hd__xor2_1 _36911_ (.A(_02640_),
    .B(_15703_),
    .X(_15704_));
 sky130_fd_sc_hd__inv_1 _36912_ (.A(\inst$top.soc.cpu.multiplier.m_prod[53] ),
    .Y(_15705_));
 sky130_fd_sc_hd__a21oi_1 _36913_ (.A1(net1929),
    .A2(_15705_),
    .B1(net3012),
    .Y(_15706_));
 sky130_fd_sc_hd__o21ai_0 _36914_ (.A1(net1929),
    .A2(_15704_),
    .B1(_15706_),
    .Y(_15707_));
 sky130_fd_sc_hd__inv_2 _36915_ (.A(_15707_),
    .Y(_04401_));
 sky130_fd_sc_hd__nand2_1 _36916_ (.A(_15394_),
    .B(_15390_),
    .Y(_15708_));
 sky130_fd_sc_hd__nor2_1 _36917_ (.A(_15400_),
    .B(_15463_),
    .Y(_15709_));
 sky130_fd_sc_hd__inv_1 _36918_ (.A(_15709_),
    .Y(_15710_));
 sky130_fd_sc_hd__inv_1 _36919_ (.A(_15569_),
    .Y(_15711_));
 sky130_fd_sc_hd__nand2_1 _36920_ (.A(_02634_),
    .B(_02640_),
    .Y(_15712_));
 sky130_fd_sc_hd__nor2_1 _36921_ (.A(_15674_),
    .B(_15712_),
    .Y(_15713_));
 sky130_fd_sc_hd__inv_1 _36922_ (.A(_15713_),
    .Y(_15714_));
 sky130_fd_sc_hd__nor2_1 _36923_ (.A(_15637_),
    .B(_15714_),
    .Y(_15715_));
 sky130_fd_sc_hd__inv_1 _36924_ (.A(_15715_),
    .Y(_15716_));
 sky130_fd_sc_hd__nor2_1 _36925_ (.A(_15711_),
    .B(_15716_),
    .Y(_15717_));
 sky130_fd_sc_hd__inv_1 _36926_ (.A(_15717_),
    .Y(_15718_));
 sky130_fd_sc_hd__nor3_1 _36927_ (.A(_15708_),
    .B(_15710_),
    .C(_15718_),
    .Y(_15719_));
 sky130_fd_sc_hd__nand2_1 _36928_ (.A(_15255_),
    .B(_15719_),
    .Y(_15720_));
 sky130_fd_sc_hd__a21oi_1 _36929_ (.A1(_02640_),
    .A2(_02633_),
    .B1(_02639_),
    .Y(_15721_));
 sky130_fd_sc_hd__inv_1 _36930_ (.A(_15721_),
    .Y(_15722_));
 sky130_fd_sc_hd__a31oi_1 _36931_ (.A1(_15679_),
    .A2(_02634_),
    .A3(_02640_),
    .B1(_15722_),
    .Y(_15723_));
 sky130_fd_sc_hd__o21ai_0 _36932_ (.A1(_15714_),
    .A2(_15645_),
    .B1(_15723_),
    .Y(_15724_));
 sky130_fd_sc_hd__a21oi_1 _36933_ (.A1(_15573_),
    .A2(_15715_),
    .B1(_15724_),
    .Y(_15725_));
 sky130_fd_sc_hd__nand2_1 _36934_ (.A(_15403_),
    .B(_15390_),
    .Y(_15726_));
 sky130_fd_sc_hd__a21oi_1 _36935_ (.A1(_15726_),
    .A2(_15399_),
    .B1(_15710_),
    .Y(_15727_));
 sky130_fd_sc_hd__o21ai_0 _36936_ (.A1(_15463_),
    .A2(_15407_),
    .B1(_15466_),
    .Y(_15728_));
 sky130_fd_sc_hd__o21ai_0 _36937_ (.A1(_15727_),
    .A2(_15728_),
    .B1(_15717_),
    .Y(_15729_));
 sky130_fd_sc_hd__nand3_1 _36938_ (.A(_15720_),
    .B(_15725_),
    .C(_15729_),
    .Y(_15730_));
 sky130_fd_sc_hd__xor2_1 _36939_ (.A(_02647_),
    .B(_15730_),
    .X(_15731_));
 sky130_fd_sc_hd__inv_1 _36940_ (.A(\inst$top.soc.cpu.multiplier.m_prod[54] ),
    .Y(_15732_));
 sky130_fd_sc_hd__a21oi_1 _36941_ (.A1(net1930),
    .A2(_15732_),
    .B1(net3012),
    .Y(_15733_));
 sky130_fd_sc_hd__o21ai_0 _36942_ (.A1(net1931),
    .A2(_15731_),
    .B1(_15733_),
    .Y(_15734_));
 sky130_fd_sc_hd__inv_2 _36943_ (.A(_15734_),
    .Y(_04402_));
 sky130_fd_sc_hd__a21oi_1 _36945_ (.A1(_15422_),
    .A2(_15416_),
    .B1(_15424_),
    .Y(_15736_));
 sky130_fd_sc_hd__nand2_1 _36946_ (.A(_15418_),
    .B(_15473_),
    .Y(_15737_));
 sky130_fd_sc_hd__o21a_1 _36947_ (.A1(_15474_),
    .A2(_15427_),
    .B1(_15478_),
    .X(_15738_));
 sky130_fd_sc_hd__o21a_1 _36948_ (.A1(_15736_),
    .A2(_15737_),
    .B1(_15738_),
    .X(_15739_));
 sky130_fd_sc_hd__inv_1 _36949_ (.A(_15583_),
    .Y(_15740_));
 sky130_fd_sc_hd__nand2_1 _36950_ (.A(_02640_),
    .B(_02647_),
    .Y(_15741_));
 sky130_fd_sc_hd__nor2_1 _36951_ (.A(_15687_),
    .B(_15741_),
    .Y(_15742_));
 sky130_fd_sc_hd__inv_1 _36952_ (.A(_15742_),
    .Y(_15743_));
 sky130_fd_sc_hd__nor2_1 _36953_ (.A(_15656_),
    .B(_15743_),
    .Y(_15744_));
 sky130_fd_sc_hd__inv_1 _36954_ (.A(_15744_),
    .Y(_15745_));
 sky130_fd_sc_hd__nor2_1 _36955_ (.A(_15740_),
    .B(_15745_),
    .Y(_15746_));
 sky130_fd_sc_hd__inv_1 _36956_ (.A(_15746_),
    .Y(_15747_));
 sky130_fd_sc_hd__a21oi_1 _36957_ (.A1(_02647_),
    .A2(_02639_),
    .B1(_02646_),
    .Y(_15748_));
 sky130_fd_sc_hd__inv_1 _36958_ (.A(_15748_),
    .Y(_15749_));
 sky130_fd_sc_hd__a31oi_1 _36959_ (.A1(_02640_),
    .A2(_15698_),
    .A3(_02647_),
    .B1(_15749_),
    .Y(_15750_));
 sky130_fd_sc_hd__o21ai_0 _36960_ (.A1(_15743_),
    .A2(_15664_),
    .B1(_15750_),
    .Y(_15751_));
 sky130_fd_sc_hd__a21oi_1 _36961_ (.A1(_15588_),
    .A2(_15744_),
    .B1(_15751_),
    .Y(_15752_));
 sky130_fd_sc_hd__nand2_1 _36962_ (.A(_15414_),
    .B(_15416_),
    .Y(_15753_));
 sky130_fd_sc_hd__nor3_1 _36963_ (.A(_15753_),
    .B(_15737_),
    .C(_15747_),
    .Y(_15754_));
 sky130_fd_sc_hd__nand2_1 _36964_ (.A(_15268_),
    .B(_15754_),
    .Y(_15755_));
 sky130_fd_sc_hd__o211ai_1 _36965_ (.A1(_15739_),
    .A2(_15747_),
    .B1(_15752_),
    .C1(_15755_),
    .Y(_15756_));
 sky130_fd_sc_hd__nor2_1 _36966_ (.A(_02653_),
    .B(_15756_),
    .Y(_15757_));
 sky130_fd_sc_hd__and2_1 _36967_ (.A(_15756_),
    .B(_02653_),
    .X(_15758_));
 sky130_fd_sc_hd__o21ai_0 _36968_ (.A1(_15757_),
    .A2(_15758_),
    .B1(net2307),
    .Y(_15759_));
 sky130_fd_sc_hd__o211ai_1 _36969_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[55] ),
    .A2(net2307),
    .B1(net2184),
    .C1(_15759_),
    .Y(_15760_));
 sky130_fd_sc_hd__inv_2 _36970_ (.A(_15760_),
    .Y(_04403_));
 sky130_fd_sc_hd__nand2_1 _36971_ (.A(_02647_),
    .B(_02653_),
    .Y(_15761_));
 sky130_fd_sc_hd__nor2_1 _36972_ (.A(_15712_),
    .B(_15761_),
    .Y(_15762_));
 sky130_fd_sc_hd__inv_1 _36973_ (.A(_15762_),
    .Y(_15763_));
 sky130_fd_sc_hd__nand2_1 _36974_ (.A(_02653_),
    .B(_02646_),
    .Y(_15764_));
 sky130_fd_sc_hd__inv_1 _36975_ (.A(_02652_),
    .Y(_15765_));
 sky130_fd_sc_hd__nand2_1 _36976_ (.A(_15764_),
    .B(_15765_),
    .Y(_15766_));
 sky130_fd_sc_hd__a31oi_1 _36977_ (.A1(_15722_),
    .A2(_02647_),
    .A3(_02653_),
    .B1(_15766_),
    .Y(_15767_));
 sky130_fd_sc_hd__nand4_1 _36978_ (.A(_15608_),
    .B(_15642_),
    .C(_15675_),
    .D(_15762_),
    .Y(_15768_));
 sky130_fd_sc_hd__o211ai_1 _36979_ (.A1(_15680_),
    .A2(_15763_),
    .B1(_15767_),
    .C1(_15768_),
    .Y(_15769_));
 sky130_fd_sc_hd__nor2_1 _36980_ (.A(_02659_),
    .B(_15769_),
    .Y(_15770_));
 sky130_fd_sc_hd__and2_1 _36981_ (.A(_15769_),
    .B(_02659_),
    .X(_15771_));
 sky130_fd_sc_hd__o21ai_0 _36982_ (.A1(_15770_),
    .A2(_15771_),
    .B1(net2307),
    .Y(_15772_));
 sky130_fd_sc_hd__o211ai_1 _36983_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[56] ),
    .A2(net2308),
    .B1(net2184),
    .C1(_15772_),
    .Y(_15773_));
 sky130_fd_sc_hd__inv_2 _36984_ (.A(_15773_),
    .Y(_04404_));
 sky130_fd_sc_hd__nand2_1 _36985_ (.A(_15325_),
    .B(_15379_),
    .Y(_15774_));
 sky130_fd_sc_hd__nand2_1 _36986_ (.A(_15447_),
    .B(_15499_),
    .Y(_15775_));
 sky130_fd_sc_hd__nor2_1 _36987_ (.A(_15774_),
    .B(_15775_),
    .Y(_15776_));
 sky130_fd_sc_hd__nand2_1 _36988_ (.A(_02653_),
    .B(_02659_),
    .Y(_15777_));
 sky130_fd_sc_hd__nor2_1 _36989_ (.A(_15741_),
    .B(_15777_),
    .Y(_15778_));
 sky130_fd_sc_hd__inv_1 _36990_ (.A(_15778_),
    .Y(_15779_));
 sky130_fd_sc_hd__nor2_1 _36991_ (.A(_15689_),
    .B(_15779_),
    .Y(_15780_));
 sky130_fd_sc_hd__inv_1 _36992_ (.A(_15780_),
    .Y(_15781_));
 sky130_fd_sc_hd__nor3_1 _36993_ (.A(_15614_),
    .B(_15617_),
    .C(_15781_),
    .Y(_15782_));
 sky130_fd_sc_hd__nand3b_1 _36994_ (.A_N(_15287_),
    .B(_15776_),
    .C(_15782_),
    .Y(_15783_));
 sky130_fd_sc_hd__a21oi_1 _36995_ (.A1(_15335_),
    .A2(_15379_),
    .B1(_15383_),
    .Y(_15784_));
 sky130_fd_sc_hd__o221ai_1 _36996_ (.A1(_15453_),
    .A2(_15500_),
    .B1(_15775_),
    .B2(_15784_),
    .C1(_15503_),
    .Y(_15785_));
 sky130_fd_sc_hd__a21oi_1 _36997_ (.A1(_02659_),
    .A2(_02652_),
    .B1(_02658_),
    .Y(_15786_));
 sky130_fd_sc_hd__o21a_1 _36998_ (.A1(_15777_),
    .A2(_15748_),
    .B1(_15786_),
    .X(_15787_));
 sky130_fd_sc_hd__o221ai_1 _36999_ (.A1(_15699_),
    .A2(_15779_),
    .B1(_15781_),
    .B2(_15624_),
    .C1(_15787_),
    .Y(_15788_));
 sky130_fd_sc_hd__a21oi_1 _37000_ (.A1(_15785_),
    .A2(_15782_),
    .B1(_15788_),
    .Y(_15789_));
 sky130_fd_sc_hd__a21oi_1 _37001_ (.A1(_15783_),
    .A2(_15789_),
    .B1(_02665_),
    .Y(_15790_));
 sky130_fd_sc_hd__nand3_1 _37002_ (.A(_15783_),
    .B(_02665_),
    .C(_15789_),
    .Y(_15791_));
 sky130_fd_sc_hd__nand2_1 _37003_ (.A(_15791_),
    .B(net2309),
    .Y(_15792_));
 sky130_fd_sc_hd__o221ai_1 _37004_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[57] ),
    .A2(net2309),
    .B1(_15790_),
    .B2(_15792_),
    .C1(net2186),
    .Y(_15793_));
 sky130_fd_sc_hd__inv_2 _37005_ (.A(_15793_),
    .Y(_04405_));
 sky130_fd_sc_hd__nand2_1 _37006_ (.A(_02659_),
    .B(_02665_),
    .Y(_15794_));
 sky130_fd_sc_hd__nor2_1 _37007_ (.A(_15761_),
    .B(_15794_),
    .Y(_15795_));
 sky130_fd_sc_hd__inv_1 _37008_ (.A(_15795_),
    .Y(_15796_));
 sky130_fd_sc_hd__inv_1 _37009_ (.A(_15794_),
    .Y(_15797_));
 sky130_fd_sc_hd__a21oi_1 _37010_ (.A1(_02665_),
    .A2(_02658_),
    .B1(_02664_),
    .Y(_15798_));
 sky130_fd_sc_hd__a21boi_0 _37011_ (.A1(_15766_),
    .A2(_15797_),
    .B1_N(_15798_),
    .Y(_15799_));
 sky130_fd_sc_hd__o21ai_0 _37012_ (.A1(_15796_),
    .A2(_15723_),
    .B1(_15799_),
    .Y(_15800_));
 sky130_fd_sc_hd__a31oi_1 _37013_ (.A1(_15649_),
    .A2(_15713_),
    .A3(_15795_),
    .B1(_15800_),
    .Y(_15801_));
 sky130_fd_sc_hd__nor2_1 _37014_ (.A(_02671_),
    .B(_15801_),
    .Y(_15802_));
 sky130_fd_sc_hd__nand2_1 _37015_ (.A(_15801_),
    .B(_02671_),
    .Y(_15803_));
 sky130_fd_sc_hd__nand2_1 _37016_ (.A(_15803_),
    .B(net2305),
    .Y(_15804_));
 sky130_fd_sc_hd__o221ai_1 _37017_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[58] ),
    .A2(net2306),
    .B1(_15802_),
    .B2(_15804_),
    .C1(net2184),
    .Y(_15805_));
 sky130_fd_sc_hd__inv_2 _37018_ (.A(_15805_),
    .Y(_04406_));
 sky130_fd_sc_hd__nand2_1 _37019_ (.A(_02665_),
    .B(_02671_),
    .Y(_15806_));
 sky130_fd_sc_hd__nor2_1 _37020_ (.A(_15777_),
    .B(_15806_),
    .Y(_15807_));
 sky130_fd_sc_hd__inv_1 _37021_ (.A(_15807_),
    .Y(_15808_));
 sky130_fd_sc_hd__a21oi_1 _37022_ (.A1(_02671_),
    .A2(_02664_),
    .B1(_02670_),
    .Y(_15809_));
 sky130_fd_sc_hd__o21ai_0 _37023_ (.A1(_15806_),
    .A2(_15786_),
    .B1(_15809_),
    .Y(_15810_));
 sky130_fd_sc_hd__o21bai_1 _37024_ (.A1(_15808_),
    .A2(_15750_),
    .B1_N(_15810_),
    .Y(_15811_));
 sky130_fd_sc_hd__a31oi_1 _37025_ (.A1(_15668_),
    .A2(_15742_),
    .A3(_15807_),
    .B1(_15811_),
    .Y(_15812_));
 sky130_fd_sc_hd__nor2_1 _37026_ (.A(_02677_),
    .B(_15812_),
    .Y(_15813_));
 sky130_fd_sc_hd__nand2_1 _37027_ (.A(_15812_),
    .B(_02677_),
    .Y(_15814_));
 sky130_fd_sc_hd__nand2_1 _37028_ (.A(_15814_),
    .B(net2300),
    .Y(_15815_));
 sky130_fd_sc_hd__o221ai_1 _37029_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[59] ),
    .A2(net2301),
    .B1(_15813_),
    .B2(_15815_),
    .C1(net2179),
    .Y(_15816_));
 sky130_fd_sc_hd__inv_2 _37030_ (.A(_15816_),
    .Y(_04407_));
 sky130_fd_sc_hd__nor2_1 _37031_ (.A(\inst$top.soc.cpu.multiplier.x_prod[5] ),
    .B(net1922),
    .Y(_15817_));
 sky130_fd_sc_hd__o21ai_0 _37032_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[5] ),
    .A2(net2299),
    .B1(net2179),
    .Y(_15818_));
 sky130_fd_sc_hd__nor2_1 _37033_ (.A(_15817_),
    .B(_15818_),
    .Y(_04408_));
 sky130_fd_sc_hd__inv_1 _37035_ (.A(_02684_),
    .Y(_15820_));
 sky130_fd_sc_hd__nand2_1 _37036_ (.A(_02671_),
    .B(_02677_),
    .Y(_15821_));
 sky130_fd_sc_hd__nand3_1 _37037_ (.A(_15797_),
    .B(_02671_),
    .C(_02677_),
    .Y(_15822_));
 sky130_fd_sc_hd__nor2_1 _37038_ (.A(_15763_),
    .B(_15822_),
    .Y(_15823_));
 sky130_fd_sc_hd__a21oi_1 _37039_ (.A1(_02677_),
    .A2(_02670_),
    .B1(_02676_),
    .Y(_15824_));
 sky130_fd_sc_hd__o21ai_0 _37040_ (.A1(_15822_),
    .A2(_15767_),
    .B1(_15824_),
    .Y(_15825_));
 sky130_fd_sc_hd__a21oi_1 _37041_ (.A1(_15681_),
    .A2(_15823_),
    .B1(_15825_),
    .Y(_15826_));
 sky130_fd_sc_hd__nand3_1 _37042_ (.A(_15548_),
    .B(_15677_),
    .C(_15823_),
    .Y(_15827_));
 sky130_fd_sc_hd__o211ai_1 _37043_ (.A1(_15798_),
    .A2(_15821_),
    .B1(_15826_),
    .C1(_15827_),
    .Y(_15828_));
 sky130_fd_sc_hd__or2_2 _37044_ (.A(_15820_),
    .B(_15828_),
    .X(_15829_));
 sky130_fd_sc_hd__nand2_1 _37045_ (.A(_15828_),
    .B(_15820_),
    .Y(_15830_));
 sky130_fd_sc_hd__nand3_1 _37046_ (.A(_15829_),
    .B(net2307),
    .C(_15830_),
    .Y(_15831_));
 sky130_fd_sc_hd__o211ai_1 _37047_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[60] ),
    .A2(net2308),
    .B1(net2185),
    .C1(_15831_),
    .Y(_15832_));
 sky130_fd_sc_hd__inv_2 _37048_ (.A(_15832_),
    .Y(_04409_));
 sky130_fd_sc_hd__nand2_1 _37049_ (.A(_02677_),
    .B(_02684_),
    .Y(_15833_));
 sky130_fd_sc_hd__nor2_1 _37050_ (.A(_15806_),
    .B(_15833_),
    .Y(_15834_));
 sky130_fd_sc_hd__inv_1 _37051_ (.A(_15834_),
    .Y(_15835_));
 sky130_fd_sc_hd__nor2_1 _37052_ (.A(_15779_),
    .B(_15835_),
    .Y(_15836_));
 sky130_fd_sc_hd__nand2_1 _37053_ (.A(_15703_),
    .B(_15836_),
    .Y(_15837_));
 sky130_fd_sc_hd__a21oi_1 _37054_ (.A1(_02684_),
    .A2(_02676_),
    .B1(_02683_),
    .Y(_15838_));
 sky130_fd_sc_hd__o21ai_0 _37055_ (.A1(_15806_),
    .A2(_15787_),
    .B1(_15809_),
    .Y(_15839_));
 sky130_fd_sc_hd__nand3_1 _37056_ (.A(_15839_),
    .B(_02677_),
    .C(_02684_),
    .Y(_15840_));
 sky130_fd_sc_hd__nand4_1 _37057_ (.A(_15837_),
    .B(_02690_),
    .C(_15838_),
    .D(_15840_),
    .Y(_15841_));
 sky130_fd_sc_hd__nand2_1 _37058_ (.A(_15841_),
    .B(net2307),
    .Y(_15842_));
 sky130_fd_sc_hd__a31oi_1 _37059_ (.A1(_15837_),
    .A2(_15838_),
    .A3(_15840_),
    .B1(_02690_),
    .Y(_15843_));
 sky130_fd_sc_hd__inv_1 _37060_ (.A(\inst$top.soc.cpu.multiplier.m_prod[61] ),
    .Y(_15844_));
 sky130_fd_sc_hd__a21oi_1 _37061_ (.A1(net1928),
    .A2(_15844_),
    .B1(net3012),
    .Y(_15845_));
 sky130_fd_sc_hd__o21ai_0 _37062_ (.A1(_15842_),
    .A2(_15843_),
    .B1(_15845_),
    .Y(_15846_));
 sky130_fd_sc_hd__inv_2 _37063_ (.A(_15846_),
    .Y(_04410_));
 sky130_fd_sc_hd__inv_1 _37064_ (.A(_02690_),
    .Y(_15847_));
 sky130_fd_sc_hd__nor3_1 _37065_ (.A(_15820_),
    .B(_15847_),
    .C(_15821_),
    .Y(_15848_));
 sky130_fd_sc_hd__inv_1 _37066_ (.A(_15848_),
    .Y(_15849_));
 sky130_fd_sc_hd__nor2_1 _37067_ (.A(_15796_),
    .B(_15849_),
    .Y(_15850_));
 sky130_fd_sc_hd__nor2_1 _37068_ (.A(_15849_),
    .B(_15799_),
    .Y(_15851_));
 sky130_fd_sc_hd__a21oi_1 _37069_ (.A1(_02690_),
    .A2(_02683_),
    .B1(_02689_),
    .Y(_15852_));
 sky130_fd_sc_hd__o31ai_1 _37070_ (.A1(_15820_),
    .A2(_15847_),
    .A3(_15824_),
    .B1(_15852_),
    .Y(_15853_));
 sky130_fd_sc_hd__inv_1 _37071_ (.A(_15850_),
    .Y(_15854_));
 sky130_fd_sc_hd__a21oi_1 _37072_ (.A1(_15728_),
    .A2(_15569_),
    .B1(_15573_),
    .Y(_15855_));
 sky130_fd_sc_hd__nor3_1 _37073_ (.A(_15716_),
    .B(_15854_),
    .C(_15855_),
    .Y(_15856_));
 sky130_fd_sc_hd__a2111oi_0 _37074_ (.A1(_15724_),
    .A2(_15850_),
    .B1(_15851_),
    .C1(_15853_),
    .D1(_15856_),
    .Y(_15857_));
 sky130_fd_sc_hd__nor4_1 _37075_ (.A(_15710_),
    .B(_15711_),
    .C(_15716_),
    .D(_15854_),
    .Y(_15858_));
 sky130_fd_sc_hd__nand2_1 _37076_ (.A(_15348_),
    .B(_15858_),
    .Y(_15859_));
 sky130_fd_sc_hd__a21oi_1 _37077_ (.A1(_15857_),
    .A2(_15859_),
    .B1(_02698_),
    .Y(_15860_));
 sky130_fd_sc_hd__nand3_1 _37078_ (.A(_15857_),
    .B(_02698_),
    .C(_15859_),
    .Y(_15861_));
 sky130_fd_sc_hd__nand2_1 _37079_ (.A(_15861_),
    .B(net2309),
    .Y(_15862_));
 sky130_fd_sc_hd__o221ai_1 _37080_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[62] ),
    .A2(net2309),
    .B1(_15860_),
    .B2(_15862_),
    .C1(net2186),
    .Y(_15863_));
 sky130_fd_sc_hd__inv_2 _37081_ (.A(_15863_),
    .Y(_04411_));
 sky130_fd_sc_hd__o22ai_1 _37082_ (.A1(_06005_),
    .A2(net1482),
    .B1(net1739),
    .B2(net1106),
    .Y(_15864_));
 sky130_fd_sc_hd__xnor2_1 _37083_ (.A(_02536_),
    .B(_02338_),
    .Y(_15865_));
 sky130_fd_sc_hd__xnor2_1 _37084_ (.A(_02526_),
    .B(_02337_),
    .Y(_15866_));
 sky130_fd_sc_hd__xnor2_1 _37085_ (.A(_15865_),
    .B(_15866_),
    .Y(_15867_));
 sky130_fd_sc_hd__xnor2_1 _37086_ (.A(_02519_),
    .B(_02514_),
    .Y(_15868_));
 sky130_fd_sc_hd__xor2_1 _37087_ (.A(_02521_),
    .B(_15868_),
    .X(_15869_));
 sky130_fd_sc_hd__xnor2_1 _37088_ (.A(_02398_),
    .B(_02397_),
    .Y(_15870_));
 sky130_fd_sc_hd__xnor2_1 _37089_ (.A(_02534_),
    .B(_02538_),
    .Y(_15871_));
 sky130_fd_sc_hd__xnor2_1 _37090_ (.A(_15870_),
    .B(_15871_),
    .Y(_15872_));
 sky130_fd_sc_hd__xnor2_1 _37091_ (.A(_15869_),
    .B(_15872_),
    .Y(_15873_));
 sky130_fd_sc_hd__xor2_1 _37092_ (.A(_15867_),
    .B(_15873_),
    .X(_15874_));
 sky130_fd_sc_hd__xnor2_1 _37093_ (.A(_15864_),
    .B(_15874_),
    .Y(_15875_));
 sky130_fd_sc_hd__xnor2_1 _37094_ (.A(_02533_),
    .B(net818),
    .Y(_15876_));
 sky130_fd_sc_hd__xor2_1 _37095_ (.A(_02693_),
    .B(_15876_),
    .X(_15877_));
 sky130_fd_sc_hd__xnor2_2 _37096_ (.A(_02176_),
    .B(_02175_),
    .Y(_15878_));
 sky130_fd_sc_hd__xnor2_1 _37097_ (.A(_02532_),
    .B(_02531_),
    .Y(_15879_));
 sky130_fd_sc_hd__xnor2_1 _37098_ (.A(_15878_),
    .B(_15879_),
    .Y(_15880_));
 sky130_fd_sc_hd__xnor2_1 _37099_ (.A(_02516_),
    .B(_02530_),
    .Y(_15881_));
 sky130_fd_sc_hd__xor2_1 _37100_ (.A(_02499_),
    .B(_02523_),
    .X(_15882_));
 sky130_fd_sc_hd__xnor2_1 _37101_ (.A(_15881_),
    .B(_15882_),
    .Y(_15883_));
 sky130_fd_sc_hd__xnor2_1 _37102_ (.A(_15880_),
    .B(_15883_),
    .Y(_15884_));
 sky130_fd_sc_hd__xor2_1 _37103_ (.A(_15877_),
    .B(_15884_),
    .X(_15885_));
 sky130_fd_sc_hd__xor2_1 _37104_ (.A(_02511_),
    .B(_15885_),
    .X(_15886_));
 sky130_fd_sc_hd__xor2_1 _37105_ (.A(_15875_),
    .B(_15886_),
    .X(_15887_));
 sky130_fd_sc_hd__nand2_1 _37106_ (.A(_15590_),
    .B(_15744_),
    .Y(_15888_));
 sky130_fd_sc_hd__inv_1 _37107_ (.A(_02698_),
    .Y(_15889_));
 sky130_fd_sc_hd__nor3_1 _37108_ (.A(_15847_),
    .B(_15889_),
    .C(_15838_),
    .Y(_15890_));
 sky130_fd_sc_hd__a211oi_1 _37109_ (.A1(_02698_),
    .A2(_02689_),
    .B1(_02697_),
    .C1(_15890_),
    .Y(_15891_));
 sky130_fd_sc_hd__nor3_1 _37110_ (.A(_15847_),
    .B(_15889_),
    .C(_15833_),
    .Y(_15892_));
 sky130_fd_sc_hd__nand2_1 _37111_ (.A(_15810_),
    .B(_15892_),
    .Y(_15893_));
 sky130_fd_sc_hd__nand2_1 _37112_ (.A(_15891_),
    .B(_15893_),
    .Y(_15894_));
 sky130_fd_sc_hd__nor2_1 _37113_ (.A(_15751_),
    .B(_15894_),
    .Y(_15895_));
 sky130_fd_sc_hd__nand2_1 _37114_ (.A(_15888_),
    .B(_15895_),
    .Y(_15896_));
 sky130_fd_sc_hd__nand2_1 _37115_ (.A(_15892_),
    .B(_15807_),
    .Y(_15897_));
 sky130_fd_sc_hd__nand3_1 _37116_ (.A(_15891_),
    .B(_15893_),
    .C(_15897_),
    .Y(_15898_));
 sky130_fd_sc_hd__nand2_1 _37117_ (.A(_15896_),
    .B(_15898_),
    .Y(_15899_));
 sky130_fd_sc_hd__xor2_1 _37118_ (.A(_15887_),
    .B(_15899_),
    .X(_15900_));
 sky130_fd_sc_hd__inv_1 _37119_ (.A(\inst$top.soc.cpu.multiplier.m_prod[63] ),
    .Y(_15901_));
 sky130_fd_sc_hd__a21oi_1 _37120_ (.A1(net1919),
    .A2(_15901_),
    .B1(net3007),
    .Y(_15902_));
 sky130_fd_sc_hd__o21ai_0 _37121_ (.A1(net1919),
    .A2(_15900_),
    .B1(_15902_),
    .Y(_15903_));
 sky130_fd_sc_hd__inv_2 _37122_ (.A(_15903_),
    .Y(_04412_));
 sky130_fd_sc_hd__nor2_1 _37124_ (.A(\inst$top.soc.cpu.multiplier.x_prod[6] ),
    .B(net1922),
    .Y(_15905_));
 sky130_fd_sc_hd__o21ai_0 _37126_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[6] ),
    .A2(net2300),
    .B1(net2179),
    .Y(_15907_));
 sky130_fd_sc_hd__nor2_1 _37127_ (.A(_15905_),
    .B(_15907_),
    .Y(_04413_));
 sky130_fd_sc_hd__xnor2_1 _37129_ (.A(_02548_),
    .B(_03387_),
    .Y(_15909_));
 sky130_fd_sc_hd__o21ai_0 _37130_ (.A1(\inst$top.soc.cpu.multiplier.m_prod[7] ),
    .A2(net2300),
    .B1(net2179),
    .Y(_15910_));
 sky130_fd_sc_hd__a21oi_1 _37131_ (.A1(net2300),
    .A2(_15909_),
    .B1(_15910_),
    .Y(_04414_));
 sky130_fd_sc_hd__xor2_1 _37132_ (.A(_03393_),
    .B(_15127_),
    .X(_15911_));
 sky130_fd_sc_hd__nor2_1 _37133_ (.A(\inst$top.soc.cpu.multiplier.m_prod[8] ),
    .B(net2300),
    .Y(_15912_));
 sky130_fd_sc_hd__nor2_1 _37134_ (.A(net3009),
    .B(_15912_),
    .Y(_15913_));
 sky130_fd_sc_hd__o21ai_0 _37135_ (.A1(net1922),
    .A2(_15911_),
    .B1(_15913_),
    .Y(_15914_));
 sky130_fd_sc_hd__inv_2 _37136_ (.A(_15914_),
    .Y(_04415_));
 sky130_fd_sc_hd__xor2_1 _37137_ (.A(_03402_),
    .B(_15140_),
    .X(_15915_));
 sky130_fd_sc_hd__nor2_1 _37138_ (.A(\inst$top.soc.cpu.multiplier.m_prod[9] ),
    .B(net2300),
    .Y(_15916_));
 sky130_fd_sc_hd__nor2_1 _37139_ (.A(net3009),
    .B(_15916_),
    .Y(_15917_));
 sky130_fd_sc_hd__o21ai_0 _37140_ (.A1(net1922),
    .A2(_15915_),
    .B1(_15917_),
    .Y(_15918_));
 sky130_fd_sc_hd__inv_2 _37141_ (.A(_15918_),
    .Y(_04416_));
 sky130_fd_sc_hd__nor2_1 _37144_ (.A(net2881),
    .B(_15374_),
    .Y(_15921_));
 sky130_fd_sc_hd__a21oi_1 _37145_ (.A1(\inst$top.soc.cpu.multiplier.m_low ),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[0] ),
    .B1(_15921_),
    .Y(_15922_));
 sky130_fd_sc_hd__o21ai_0 _37146_ (.A1(\inst$top.soc.cpu.multiplier.w_result[0] ),
    .A2(net2282),
    .B1(net2177),
    .Y(_15923_));
 sky130_fd_sc_hd__a21oi_1 _37147_ (.A1(net2282),
    .A2(_15922_),
    .B1(_15923_),
    .Y(_04417_));
 sky130_fd_sc_hd__nor2_1 _37148_ (.A(net2875),
    .B(_15517_),
    .Y(_15924_));
 sky130_fd_sc_hd__a21oi_1 _37149_ (.A1(net2875),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[10] ),
    .B1(_15924_),
    .Y(_15925_));
 sky130_fd_sc_hd__o21ai_0 _37150_ (.A1(\inst$top.soc.cpu.multiplier.w_result[10] ),
    .A2(net2279),
    .B1(net2154),
    .Y(_15926_));
 sky130_fd_sc_hd__a21oi_1 _37151_ (.A1(net2279),
    .A2(_15925_),
    .B1(_15926_),
    .Y(_04418_));
 sky130_fd_sc_hd__inv_1 _37152_ (.A(\inst$top.soc.cpu.multiplier.m_prod[43] ),
    .Y(_15927_));
 sky130_fd_sc_hd__nor2_1 _37153_ (.A(net2875),
    .B(_15927_),
    .Y(_15928_));
 sky130_fd_sc_hd__a21oi_1 _37154_ (.A1(net2875),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[11] ),
    .B1(_15928_),
    .Y(_15929_));
 sky130_fd_sc_hd__o21ai_0 _37156_ (.A1(\inst$top.soc.cpu.multiplier.w_result[11] ),
    .A2(net2283),
    .B1(net2177),
    .Y(_15931_));
 sky130_fd_sc_hd__a21oi_1 _37157_ (.A1(net2283),
    .A2(_15929_),
    .B1(_15931_),
    .Y(_04419_));
 sky130_fd_sc_hd__nor2_1 _37158_ (.A(net2877),
    .B(_15550_),
    .Y(_15932_));
 sky130_fd_sc_hd__a21oi_1 _37159_ (.A1(net2877),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[12] ),
    .B1(_15932_),
    .Y(_15933_));
 sky130_fd_sc_hd__o21ai_0 _37160_ (.A1(\inst$top.soc.cpu.multiplier.w_result[12] ),
    .A2(net2293),
    .B1(net2181),
    .Y(_15934_));
 sky130_fd_sc_hd__a21oi_1 _37161_ (.A1(net2293),
    .A2(_15933_),
    .B1(_15934_),
    .Y(_04420_));
 sky130_fd_sc_hd__nor2_1 _37162_ (.A(net2874),
    .B(_15562_),
    .Y(_15935_));
 sky130_fd_sc_hd__a21oi_1 _37163_ (.A1(net2874),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[13] ),
    .B1(_15935_),
    .Y(_15936_));
 sky130_fd_sc_hd__o21ai_0 _37164_ (.A1(\inst$top.soc.cpu.multiplier.w_result[13] ),
    .A2(net2283),
    .B1(net2177),
    .Y(_15937_));
 sky130_fd_sc_hd__a21oi_1 _37165_ (.A1(net2282),
    .A2(_15936_),
    .B1(_15937_),
    .Y(_04421_));
 sky130_fd_sc_hd__inv_1 _37166_ (.A(\inst$top.soc.cpu.multiplier.m_prod[46] ),
    .Y(_15938_));
 sky130_fd_sc_hd__nor2_1 _37167_ (.A(net2874),
    .B(_15938_),
    .Y(_15939_));
 sky130_fd_sc_hd__a21oi_1 _37168_ (.A1(net2874),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[14] ),
    .B1(_15939_),
    .Y(_15940_));
 sky130_fd_sc_hd__o21ai_0 _37170_ (.A1(\inst$top.soc.cpu.multiplier.w_result[14] ),
    .A2(net2293),
    .B1(net2177),
    .Y(_15942_));
 sky130_fd_sc_hd__a21oi_1 _37171_ (.A1(net2282),
    .A2(_15940_),
    .B1(_15942_),
    .Y(_04422_));
 sky130_fd_sc_hd__nor2_1 _37172_ (.A(net2875),
    .B(_15592_),
    .Y(_15943_));
 sky130_fd_sc_hd__a21oi_1 _37173_ (.A1(net2875),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[15] ),
    .B1(_15943_),
    .Y(_15944_));
 sky130_fd_sc_hd__o21ai_0 _37174_ (.A1(\inst$top.soc.cpu.multiplier.w_result[15] ),
    .A2(net2301),
    .B1(net2180),
    .Y(_15945_));
 sky130_fd_sc_hd__a21oi_1 _37175_ (.A1(net2301),
    .A2(_15944_),
    .B1(_15945_),
    .Y(_04423_));
 sky130_fd_sc_hd__inv_1 _37177_ (.A(\inst$top.soc.cpu.multiplier.m_prod[48] ),
    .Y(_15947_));
 sky130_fd_sc_hd__nor2_1 _37178_ (.A(net2874),
    .B(_15947_),
    .Y(_15948_));
 sky130_fd_sc_hd__a21oi_1 _37179_ (.A1(net2874),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[16] ),
    .B1(_15948_),
    .Y(_15949_));
 sky130_fd_sc_hd__o21ai_0 _37180_ (.A1(\inst$top.soc.cpu.multiplier.w_result[16] ),
    .A2(net2303),
    .B1(net2178),
    .Y(_15950_));
 sky130_fd_sc_hd__a21oi_1 _37181_ (.A1(net2303),
    .A2(_15949_),
    .B1(_15950_),
    .Y(_04424_));
 sky130_fd_sc_hd__nor2_1 _37182_ (.A(net2878),
    .B(_15627_),
    .Y(_15951_));
 sky130_fd_sc_hd__a21oi_1 _37183_ (.A1(net2878),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[17] ),
    .B1(_15951_),
    .Y(_15952_));
 sky130_fd_sc_hd__o21ai_0 _37184_ (.A1(\inst$top.soc.cpu.multiplier.w_result[17] ),
    .A2(net2303),
    .B1(net2182),
    .Y(_15953_));
 sky130_fd_sc_hd__a21oi_1 _37185_ (.A1(net2303),
    .A2(_15952_),
    .B1(_15953_),
    .Y(_04425_));
 sky130_fd_sc_hd__nor2_1 _37187_ (.A(net2874),
    .B(_15651_),
    .Y(_15955_));
 sky130_fd_sc_hd__a21oi_1 _37188_ (.A1(net2876),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[18] ),
    .B1(_15955_),
    .Y(_15956_));
 sky130_fd_sc_hd__o21ai_0 _37189_ (.A1(\inst$top.soc.cpu.multiplier.w_result[18] ),
    .A2(net2282),
    .B1(net2177),
    .Y(_15957_));
 sky130_fd_sc_hd__a21oi_1 _37190_ (.A1(net2282),
    .A2(_15956_),
    .B1(_15957_),
    .Y(_04426_));
 sky130_fd_sc_hd__inv_1 _37192_ (.A(\inst$top.soc.cpu.multiplier.m_prod[51] ),
    .Y(_15959_));
 sky130_fd_sc_hd__nor2_1 _37193_ (.A(net2877),
    .B(_15959_),
    .Y(_15960_));
 sky130_fd_sc_hd__a21oi_1 _37194_ (.A1(net2877),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[19] ),
    .B1(_15960_),
    .Y(_15961_));
 sky130_fd_sc_hd__o21ai_0 _37195_ (.A1(\inst$top.soc.cpu.multiplier.w_result[19] ),
    .A2(net2303),
    .B1(net2182),
    .Y(_15962_));
 sky130_fd_sc_hd__a21oi_1 _37196_ (.A1(net2303),
    .A2(_15961_),
    .B1(_15962_),
    .Y(_04427_));
 sky130_fd_sc_hd__nor2_1 _37197_ (.A(net2874),
    .B(_15386_),
    .Y(_15963_));
 sky130_fd_sc_hd__a21oi_1 _37198_ (.A1(net2876),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[1] ),
    .B1(_15963_),
    .Y(_15964_));
 sky130_fd_sc_hd__o21ai_0 _37199_ (.A1(\inst$top.soc.cpu.multiplier.w_result[1] ),
    .A2(net2299),
    .B1(net2177),
    .Y(_15965_));
 sky130_fd_sc_hd__a21oi_1 _37200_ (.A1(net2299),
    .A2(_15964_),
    .B1(_15965_),
    .Y(_04428_));
 sky130_fd_sc_hd__nor2_1 _37201_ (.A(net2878),
    .B(_15684_),
    .Y(_15966_));
 sky130_fd_sc_hd__a21oi_1 _37202_ (.A1(net2879),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[20] ),
    .B1(_15966_),
    .Y(_15967_));
 sky130_fd_sc_hd__o21ai_0 _37204_ (.A1(\inst$top.soc.cpu.multiplier.w_result[20] ),
    .A2(net2303),
    .B1(net2182),
    .Y(_15969_));
 sky130_fd_sc_hd__a21oi_1 _37205_ (.A1(net2303),
    .A2(_15967_),
    .B1(_15969_),
    .Y(_04429_));
 sky130_fd_sc_hd__nor2_1 _37206_ (.A(net2877),
    .B(_15705_),
    .Y(_15970_));
 sky130_fd_sc_hd__a21oi_1 _37207_ (.A1(net2877),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[21] ),
    .B1(_15970_),
    .Y(_15971_));
 sky130_fd_sc_hd__o21ai_0 _37208_ (.A1(\inst$top.soc.cpu.multiplier.w_result[21] ),
    .A2(net2311),
    .B1(net2185),
    .Y(_15972_));
 sky130_fd_sc_hd__a21oi_1 _37209_ (.A1(net2304),
    .A2(_15971_),
    .B1(_15972_),
    .Y(_04430_));
 sky130_fd_sc_hd__nor2_1 _37210_ (.A(net2878),
    .B(_15732_),
    .Y(_15973_));
 sky130_fd_sc_hd__a21oi_1 _37211_ (.A1(net2878),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[22] ),
    .B1(_15973_),
    .Y(_15974_));
 sky130_fd_sc_hd__o21ai_0 _37212_ (.A1(\inst$top.soc.cpu.multiplier.w_result[22] ),
    .A2(net2312),
    .B1(net2185),
    .Y(_15975_));
 sky130_fd_sc_hd__a21oi_1 _37213_ (.A1(net2311),
    .A2(_15974_),
    .B1(_15975_),
    .Y(_04431_));
 sky130_fd_sc_hd__inv_1 _37214_ (.A(\inst$top.soc.cpu.multiplier.m_prod[55] ),
    .Y(_15976_));
 sky130_fd_sc_hd__nor2_1 _37215_ (.A(net2879),
    .B(_15976_),
    .Y(_15977_));
 sky130_fd_sc_hd__a21oi_1 _37216_ (.A1(net2879),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[23] ),
    .B1(_15977_),
    .Y(_15978_));
 sky130_fd_sc_hd__o21ai_0 _37218_ (.A1(\inst$top.soc.cpu.multiplier.w_result[23] ),
    .A2(net2304),
    .B1(net2185),
    .Y(_15980_));
 sky130_fd_sc_hd__a21oi_1 _37219_ (.A1(net2304),
    .A2(_15978_),
    .B1(_15980_),
    .Y(_04432_));
 sky130_fd_sc_hd__inv_1 _37220_ (.A(\inst$top.soc.cpu.multiplier.m_prod[56] ),
    .Y(_15981_));
 sky130_fd_sc_hd__nor2_1 _37221_ (.A(net2878),
    .B(_15981_),
    .Y(_15982_));
 sky130_fd_sc_hd__a21oi_1 _37222_ (.A1(net2879),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[24] ),
    .B1(_15982_),
    .Y(_15983_));
 sky130_fd_sc_hd__o21ai_0 _37223_ (.A1(\inst$top.soc.cpu.multiplier.w_result[24] ),
    .A2(net2304),
    .B1(net2185),
    .Y(_15984_));
 sky130_fd_sc_hd__a21oi_1 _37224_ (.A1(net2304),
    .A2(_15983_),
    .B1(_15984_),
    .Y(_04433_));
 sky130_fd_sc_hd__inv_1 _37226_ (.A(\inst$top.soc.cpu.multiplier.m_prod[57] ),
    .Y(_15986_));
 sky130_fd_sc_hd__nor2_1 _37227_ (.A(net2879),
    .B(_15986_),
    .Y(_15987_));
 sky130_fd_sc_hd__a21oi_1 _37228_ (.A1(net2879),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[25] ),
    .B1(_15987_),
    .Y(_15988_));
 sky130_fd_sc_hd__o21ai_0 _37229_ (.A1(\inst$top.soc.cpu.multiplier.w_result[25] ),
    .A2(net2304),
    .B1(net2185),
    .Y(_15989_));
 sky130_fd_sc_hd__a21oi_1 _37230_ (.A1(net2304),
    .A2(_15988_),
    .B1(_15989_),
    .Y(_04434_));
 sky130_fd_sc_hd__inv_1 _37231_ (.A(\inst$top.soc.cpu.multiplier.m_prod[58] ),
    .Y(_15990_));
 sky130_fd_sc_hd__nor2_1 _37232_ (.A(net2880),
    .B(_15990_),
    .Y(_15991_));
 sky130_fd_sc_hd__a21oi_1 _37233_ (.A1(net2880),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[26] ),
    .B1(_15991_),
    .Y(_15992_));
 sky130_fd_sc_hd__o21ai_0 _37234_ (.A1(\inst$top.soc.cpu.multiplier.w_result[26] ),
    .A2(net2304),
    .B1(net2180),
    .Y(_15993_));
 sky130_fd_sc_hd__a21oi_1 _37235_ (.A1(net2304),
    .A2(_15992_),
    .B1(_15993_),
    .Y(_04435_));
 sky130_fd_sc_hd__inv_1 _37237_ (.A(\inst$top.soc.cpu.multiplier.m_prod[59] ),
    .Y(_15995_));
 sky130_fd_sc_hd__nor2_1 _37238_ (.A(net2881),
    .B(_15995_),
    .Y(_15996_));
 sky130_fd_sc_hd__a21oi_1 _37239_ (.A1(net2881),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[27] ),
    .B1(_15996_),
    .Y(_15997_));
 sky130_fd_sc_hd__o21ai_0 _37240_ (.A1(\inst$top.soc.cpu.multiplier.w_result[27] ),
    .A2(net2299),
    .B1(net2178),
    .Y(_15998_));
 sky130_fd_sc_hd__a21oi_1 _37241_ (.A1(net2299),
    .A2(_15997_),
    .B1(_15998_),
    .Y(_04436_));
 sky130_fd_sc_hd__inv_1 _37243_ (.A(\inst$top.soc.cpu.multiplier.m_prod[60] ),
    .Y(_16000_));
 sky130_fd_sc_hd__nor2_1 _37244_ (.A(net2878),
    .B(_16000_),
    .Y(_16001_));
 sky130_fd_sc_hd__a21oi_1 _37245_ (.A1(net2878),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[28] ),
    .B1(_16001_),
    .Y(_16002_));
 sky130_fd_sc_hd__o21ai_0 _37246_ (.A1(\inst$top.soc.cpu.multiplier.w_result[28] ),
    .A2(net2292),
    .B1(net2173),
    .Y(_16003_));
 sky130_fd_sc_hd__a21oi_1 _37247_ (.A1(net2292),
    .A2(_16002_),
    .B1(_16003_),
    .Y(_04437_));
 sky130_fd_sc_hd__nor2_1 _37248_ (.A(net2880),
    .B(_15844_),
    .Y(_16004_));
 sky130_fd_sc_hd__a21oi_1 _37249_ (.A1(net2878),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[29] ),
    .B1(_16004_),
    .Y(_16005_));
 sky130_fd_sc_hd__o21ai_0 _37250_ (.A1(\inst$top.soc.cpu.multiplier.w_result[29] ),
    .A2(net2304),
    .B1(net2185),
    .Y(_16006_));
 sky130_fd_sc_hd__a21oi_1 _37251_ (.A1(net2311),
    .A2(_16005_),
    .B1(_16006_),
    .Y(_04438_));
 sky130_fd_sc_hd__nor2_1 _37252_ (.A(net2876),
    .B(_15411_),
    .Y(_16007_));
 sky130_fd_sc_hd__a21oi_1 _37253_ (.A1(net2876),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[2] ),
    .B1(_16007_),
    .Y(_16008_));
 sky130_fd_sc_hd__o21ai_0 _37255_ (.A1(\inst$top.soc.cpu.multiplier.w_result[2] ),
    .A2(net2302),
    .B1(net2180),
    .Y(_16010_));
 sky130_fd_sc_hd__a21oi_1 _37256_ (.A1(net2302),
    .A2(_16008_),
    .B1(_16010_),
    .Y(_04439_));
 sky130_fd_sc_hd__inv_1 _37257_ (.A(\inst$top.soc.cpu.multiplier.m_prod[62] ),
    .Y(_16011_));
 sky130_fd_sc_hd__nor2_1 _37258_ (.A(net2878),
    .B(_16011_),
    .Y(_16012_));
 sky130_fd_sc_hd__a21oi_1 _37259_ (.A1(net2879),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[30] ),
    .B1(_16012_),
    .Y(_16013_));
 sky130_fd_sc_hd__o21ai_0 _37260_ (.A1(\inst$top.soc.cpu.multiplier.w_result[30] ),
    .A2(net2303),
    .B1(net2182),
    .Y(_16014_));
 sky130_fd_sc_hd__a21oi_1 _37261_ (.A1(net2303),
    .A2(_16013_),
    .B1(_16014_),
    .Y(_04440_));
 sky130_fd_sc_hd__nor2_1 _37262_ (.A(net2874),
    .B(_15901_),
    .Y(_16015_));
 sky130_fd_sc_hd__a21oi_1 _37263_ (.A1(net2874),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[31] ),
    .B1(_16015_),
    .Y(_16016_));
 sky130_fd_sc_hd__o21ai_0 _37264_ (.A1(\inst$top.soc.cpu.multiplier.w_result[31] ),
    .A2(net2302),
    .B1(net2180),
    .Y(_16017_));
 sky130_fd_sc_hd__a21oi_1 _37265_ (.A1(net2299),
    .A2(_16016_),
    .B1(_16017_),
    .Y(_04441_));
 sky130_fd_sc_hd__nor2_1 _37266_ (.A(net2876),
    .B(_15433_),
    .Y(_16018_));
 sky130_fd_sc_hd__a21oi_1 _37267_ (.A1(net2876),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[3] ),
    .B1(_16018_),
    .Y(_16019_));
 sky130_fd_sc_hd__o21ai_0 _37269_ (.A1(\inst$top.soc.cpu.multiplier.w_result[3] ),
    .A2(net2278),
    .B1(net2155),
    .Y(_16021_));
 sky130_fd_sc_hd__a21oi_1 _37270_ (.A1(net2278),
    .A2(_16019_),
    .B1(_16021_),
    .Y(_04442_));
 sky130_fd_sc_hd__nor2_1 _37271_ (.A(net2876),
    .B(_15442_),
    .Y(_16022_));
 sky130_fd_sc_hd__a21oi_1 _37272_ (.A1(net2876),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[4] ),
    .B1(_16022_),
    .Y(_16023_));
 sky130_fd_sc_hd__o21ai_0 _37273_ (.A1(\inst$top.soc.cpu.multiplier.w_result[4] ),
    .A2(net2278),
    .B1(net2155),
    .Y(_16024_));
 sky130_fd_sc_hd__a21oi_1 _37274_ (.A1(net2278),
    .A2(_16023_),
    .B1(_16024_),
    .Y(_04443_));
 sky130_fd_sc_hd__nor2_1 _37275_ (.A(net2881),
    .B(_15458_),
    .Y(_16025_));
 sky130_fd_sc_hd__a21oi_1 _37276_ (.A1(net2876),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[5] ),
    .B1(_16025_),
    .Y(_16026_));
 sky130_fd_sc_hd__o21ai_0 _37277_ (.A1(\inst$top.soc.cpu.multiplier.w_result[5] ),
    .A2(net2283),
    .B1(net2177),
    .Y(_16027_));
 sky130_fd_sc_hd__a21oi_1 _37278_ (.A1(net2283),
    .A2(_16026_),
    .B1(_16027_),
    .Y(_04444_));
 sky130_fd_sc_hd__nor2_1 _37279_ (.A(net2875),
    .B(_15469_),
    .Y(_16028_));
 sky130_fd_sc_hd__a21oi_1 _37280_ (.A1(net2875),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[6] ),
    .B1(_16028_),
    .Y(_16029_));
 sky130_fd_sc_hd__o21ai_0 _37281_ (.A1(\inst$top.soc.cpu.multiplier.w_result[6] ),
    .A2(net2282),
    .B1(net2177),
    .Y(_16030_));
 sky130_fd_sc_hd__a21oi_1 _37282_ (.A1(net2282),
    .A2(_16029_),
    .B1(_16030_),
    .Y(_04445_));
 sky130_fd_sc_hd__nor2_1 _37283_ (.A(net2875),
    .B(_15481_),
    .Y(_16031_));
 sky130_fd_sc_hd__a21oi_1 _37284_ (.A1(net2875),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[7] ),
    .B1(_16031_),
    .Y(_16032_));
 sky130_fd_sc_hd__o21ai_0 _37285_ (.A1(\inst$top.soc.cpu.multiplier.w_result[7] ),
    .A2(net2278),
    .B1(net2155),
    .Y(_16033_));
 sky130_fd_sc_hd__a21oi_1 _37286_ (.A1(net2278),
    .A2(_16032_),
    .B1(_16033_),
    .Y(_04446_));
 sky130_fd_sc_hd__nor2_1 _37287_ (.A(net2877),
    .B(_15495_),
    .Y(_16034_));
 sky130_fd_sc_hd__a21oi_1 _37288_ (.A1(net2877),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[8] ),
    .B1(_16034_),
    .Y(_16035_));
 sky130_fd_sc_hd__o21ai_0 _37289_ (.A1(\inst$top.soc.cpu.multiplier.w_result[8] ),
    .A2(net2293),
    .B1(net2181),
    .Y(_16036_));
 sky130_fd_sc_hd__a21oi_1 _37290_ (.A1(net2293),
    .A2(_16035_),
    .B1(_16036_),
    .Y(_04447_));
 sky130_fd_sc_hd__nor2_1 _37291_ (.A(net2877),
    .B(_15506_),
    .Y(_16037_));
 sky130_fd_sc_hd__a21oi_1 _37292_ (.A1(net2877),
    .A2(\inst$top.soc.cpu.multiplier.m_prod[9] ),
    .B1(_16037_),
    .Y(_16038_));
 sky130_fd_sc_hd__o21ai_0 _37293_ (.A1(\inst$top.soc.cpu.multiplier.w_result[9] ),
    .A2(net2289),
    .B1(net2172),
    .Y(_16039_));
 sky130_fd_sc_hd__a21oi_1 _37294_ (.A1(net2289),
    .A2(_16038_),
    .B1(_16039_),
    .Y(_04448_));
 sky130_fd_sc_hd__nor2_1 _37295_ (.A(\inst$top.soc.cpu.multiplier.x_low ),
    .B(net700),
    .Y(_16040_));
 sky130_fd_sc_hd__nand2_1 _37296_ (.A(_20353_),
    .B(_11908_),
    .Y(_16041_));
 sky130_fd_sc_hd__inv_1 _37297_ (.A(_16041_),
    .Y(_16042_));
 sky130_fd_sc_hd__o21ai_1 _37298_ (.A1(_16042_),
    .A2(net654),
    .B1(net2147),
    .Y(_16043_));
 sky130_fd_sc_hd__nor2_4 _37299_ (.A(_16040_),
    .B(_16043_),
    .Y(_04449_));
 sky130_fd_sc_hd__nor2_1 _37300_ (.A(\inst$top.soc.cpu.multiplier.x_src1_signed ),
    .B(net700),
    .Y(_16044_));
 sky130_fd_sc_hd__nand2_1 _37301_ (.A(\inst$top.soc.cpu.sink__payload$6[45] ),
    .B(\inst$top.soc.cpu.sink__payload$6[44] ),
    .Y(_16045_));
 sky130_fd_sc_hd__inv_1 _37302_ (.A(_16045_),
    .Y(_16046_));
 sky130_fd_sc_hd__nor3_1 _37303_ (.A(\inst$top.soc.cpu.csr_fmt_i ),
    .B(_20353_),
    .C(_16046_),
    .Y(_16047_));
 sky130_fd_sc_hd__o21ai_1 _37304_ (.A1(_16047_),
    .A2(net654),
    .B1(net2147),
    .Y(_16048_));
 sky130_fd_sc_hd__nor2_4 _37305_ (.A(_16044_),
    .B(_16048_),
    .Y(_04450_));
 sky130_fd_sc_hd__nor2_1 _37306_ (.A(\inst$top.soc.cpu.multiplier.x_src2_signed ),
    .B(net699),
    .Y(_16049_));
 sky130_fd_sc_hd__inv_1 _37307_ (.A(\inst$top.soc.cpu.sink__payload$6[44] ),
    .Y(_16050_));
 sky130_fd_sc_hd__nor2_1 _37308_ (.A(\inst$top.soc.cpu.sink__payload$6[45] ),
    .B(_16050_),
    .Y(_16051_));
 sky130_fd_sc_hd__inv_1 _37309_ (.A(_16051_),
    .Y(_16052_));
 sky130_fd_sc_hd__nor2_1 _37310_ (.A(\inst$top.soc.cpu.csr_fmt_i ),
    .B(_16052_),
    .Y(_16053_));
 sky130_fd_sc_hd__o21ai_1 _37311_ (.A1(_16053_),
    .A2(net655),
    .B1(net2178),
    .Y(_16054_));
 sky130_fd_sc_hd__nor2_4 _37312_ (.A(_16049_),
    .B(_16054_),
    .Y(_04451_));
 sky130_fd_sc_hd__clkinv_1 _37313_ (.A(net2857),
    .Y(_16055_));
 sky130_fd_sc_hd__o21ai_0 _37317_ (.A1(net2873),
    .A2(net2294),
    .B1(net2182),
    .Y(_16059_));
 sky130_fd_sc_hd__a21oi_1 _37318_ (.A1(net2000),
    .A2(net2293),
    .B1(_16059_),
    .Y(_04452_));
 sky130_fd_sc_hd__nand2_1 _37322_ (.A(net1466),
    .B(net2857),
    .Y(_16063_));
 sky130_fd_sc_hd__o21ai_0 _37323_ (.A1(net2857),
    .A2(net1368),
    .B1(_16063_),
    .Y(_16064_));
 sky130_fd_sc_hd__nand2_1 _37324_ (.A(net1736),
    .B(net2857),
    .Y(_16065_));
 sky130_fd_sc_hd__o21ai_0 _37325_ (.A1(net2857),
    .A2(net1365),
    .B1(_16065_),
    .Y(_16066_));
 sky130_fd_sc_hd__nand2_1 _37326_ (.A(_16066_),
    .B(net1686),
    .Y(_16067_));
 sky130_fd_sc_hd__o21ai_0 _37327_ (.A1(net1686),
    .A2(_16064_),
    .B1(_16067_),
    .Y(_16068_));
 sky130_fd_sc_hd__nand2_1 _37328_ (.A(_16068_),
    .B(net1701),
    .Y(_16069_));
 sky130_fd_sc_hd__nand2_1 _37331_ (.A(net1481),
    .B(net2857),
    .Y(_16072_));
 sky130_fd_sc_hd__o21ai_0 _37332_ (.A1(net2857),
    .A2(net1695),
    .B1(_16072_),
    .Y(_16073_));
 sky130_fd_sc_hd__nand2_1 _37333_ (.A(net1708),
    .B(net2000),
    .Y(_16074_));
 sky130_fd_sc_hd__o21ai_0 _37334_ (.A1(net2000),
    .A2(net1476),
    .B1(_16074_),
    .Y(_16075_));
 sky130_fd_sc_hd__nand2_1 _37335_ (.A(_16075_),
    .B(net1686),
    .Y(_16076_));
 sky130_fd_sc_hd__o21ai_0 _37336_ (.A1(net1686),
    .A2(_16073_),
    .B1(_16076_),
    .Y(_16077_));
 sky130_fd_sc_hd__nand2_1 _37338_ (.A(_16077_),
    .B(net1382),
    .Y(_16079_));
 sky130_fd_sc_hd__nand2_1 _37339_ (.A(net1117),
    .B(net2857),
    .Y(_16080_));
 sky130_fd_sc_hd__o21ai_0 _37340_ (.A1(net2857),
    .A2(net1360),
    .B1(_16080_),
    .Y(_16081_));
 sky130_fd_sc_hd__nand2_1 _37341_ (.A(net1354),
    .B(net2000),
    .Y(_16082_));
 sky130_fd_sc_hd__o21ai_0 _37342_ (.A1(net2000),
    .A2(net1669),
    .B1(_16082_),
    .Y(_16083_));
 sky130_fd_sc_hd__nand2_1 _37343_ (.A(_16083_),
    .B(net1685),
    .Y(_16084_));
 sky130_fd_sc_hd__o21ai_0 _37344_ (.A1(net1686),
    .A2(_16081_),
    .B1(_16084_),
    .Y(_16085_));
 sky130_fd_sc_hd__nand2_1 _37345_ (.A(net1271),
    .B(net2858),
    .Y(_16086_));
 sky130_fd_sc_hd__o21ai_0 _37346_ (.A1(net2858),
    .A2(_05901_),
    .B1(_16086_),
    .Y(_16087_));
 sky130_fd_sc_hd__nand2_1 _37347_ (.A(net1672),
    .B(net2858),
    .Y(_16088_));
 sky130_fd_sc_hd__o21ai_0 _37348_ (.A1(net2858),
    .A2(net1349),
    .B1(_16088_),
    .Y(_16089_));
 sky130_fd_sc_hd__nand2_1 _37349_ (.A(_16089_),
    .B(net1250),
    .Y(_16090_));
 sky130_fd_sc_hd__o21ai_0 _37350_ (.A1(net1250),
    .A2(_16087_),
    .B1(_16090_),
    .Y(_16091_));
 sky130_fd_sc_hd__nand2_1 _37351_ (.A(_16091_),
    .B(net1700),
    .Y(_16092_));
 sky130_fd_sc_hd__o21ai_0 _37352_ (.A1(net1701),
    .A2(_16085_),
    .B1(_16092_),
    .Y(_16093_));
 sky130_fd_sc_hd__nor2_1 _37353_ (.A(net1388),
    .B(_16093_),
    .Y(_16094_));
 sky130_fd_sc_hd__a31oi_1 _37354_ (.A1(net1388),
    .A2(_16069_),
    .A3(_16079_),
    .B1(_16094_),
    .Y(_16095_));
 sky130_fd_sc_hd__nand2_1 _37356_ (.A(net1146),
    .B(net1999),
    .Y(_16097_));
 sky130_fd_sc_hd__o21ai_0 _37357_ (.A1(net1999),
    .A2(net1296),
    .B1(_16097_),
    .Y(_16098_));
 sky130_fd_sc_hd__nand2_1 _37358_ (.A(net1144),
    .B(net1999),
    .Y(_16099_));
 sky130_fd_sc_hd__o21ai_0 _37359_ (.A1(net1999),
    .A2(net1302),
    .B1(_16099_),
    .Y(_16100_));
 sky130_fd_sc_hd__mux2i_1 _37360_ (.A0(_16098_),
    .A1(_16100_),
    .S(net1688),
    .Y(_16101_));
 sky130_fd_sc_hd__nand2_1 _37361_ (.A(net1151),
    .B(net1999),
    .Y(_16102_));
 sky130_fd_sc_hd__o21ai_0 _37362_ (.A1(net1999),
    .A2(net1288),
    .B1(_16102_),
    .Y(_16103_));
 sky130_fd_sc_hd__nand2_1 _37363_ (.A(net1148),
    .B(net1999),
    .Y(_16104_));
 sky130_fd_sc_hd__o21ai_0 _37364_ (.A1(net1999),
    .A2(net1292),
    .B1(_16104_),
    .Y(_16105_));
 sky130_fd_sc_hd__mux2i_1 _37365_ (.A0(_16103_),
    .A1(_16105_),
    .S(net1688),
    .Y(_16106_));
 sky130_fd_sc_hd__or2_2 _37366_ (.A(net1700),
    .B(_16106_),
    .X(_16107_));
 sky130_fd_sc_hd__o21ai_0 _37367_ (.A1(net1385),
    .A2(_16101_),
    .B1(_16107_),
    .Y(_16108_));
 sky130_fd_sc_hd__nand2_1 _37368_ (.A(net1129),
    .B(net2858),
    .Y(_16109_));
 sky130_fd_sc_hd__o21ai_0 _37369_ (.A1(net2858),
    .A2(net1326),
    .B1(_16109_),
    .Y(_16110_));
 sky130_fd_sc_hd__nand2_1 _37370_ (.A(_16110_),
    .B(net1685),
    .Y(_16111_));
 sky130_fd_sc_hd__nand2_1 _37371_ (.A(net1126),
    .B(net2858),
    .Y(_16112_));
 sky130_fd_sc_hd__o21ai_0 _37372_ (.A1(net2858),
    .A2(net1330),
    .B1(_16112_),
    .Y(_16113_));
 sky130_fd_sc_hd__nand2_1 _37373_ (.A(_16113_),
    .B(net1250),
    .Y(_16114_));
 sky130_fd_sc_hd__nand2_1 _37374_ (.A(_16111_),
    .B(_16114_),
    .Y(_16115_));
 sky130_fd_sc_hd__nand2_1 _37375_ (.A(net1157),
    .B(net2000),
    .Y(_16116_));
 sky130_fd_sc_hd__o21ai_0 _37376_ (.A1(net2000),
    .A2(net1273),
    .B1(_16116_),
    .Y(_16117_));
 sky130_fd_sc_hd__nand2_1 _37377_ (.A(net1677),
    .B(net2858),
    .Y(_16118_));
 sky130_fd_sc_hd__o21ai_0 _37378_ (.A1(net2858),
    .A2(net1334),
    .B1(_16118_),
    .Y(_16119_));
 sky130_fd_sc_hd__mux2i_1 _37379_ (.A0(_16117_),
    .A1(_16119_),
    .S(net1685),
    .Y(_16120_));
 sky130_fd_sc_hd__nand2_1 _37380_ (.A(_16120_),
    .B(net1382),
    .Y(_16121_));
 sky130_fd_sc_hd__o21ai_0 _37381_ (.A1(net1383),
    .A2(_16115_),
    .B1(_16121_),
    .Y(_16122_));
 sky130_fd_sc_hd__nand2_1 _37382_ (.A(_16122_),
    .B(net1386),
    .Y(_16123_));
 sky130_fd_sc_hd__o21ai_0 _37383_ (.A1(net1386),
    .A2(_16108_),
    .B1(_16123_),
    .Y(_16124_));
 sky130_fd_sc_hd__nand2_1 _37384_ (.A(_16124_),
    .B(net1178),
    .Y(_16125_));
 sky130_fd_sc_hd__o21ai_0 _37385_ (.A1(net1178),
    .A2(_16095_),
    .B1(_16125_),
    .Y(_16126_));
 sky130_fd_sc_hd__nand2_1 _37386_ (.A(_16126_),
    .B(net1073),
    .Y(_16127_));
 sky130_fd_sc_hd__nand2_1 _37388_ (.A(_05901_),
    .B(net2860),
    .Y(_16129_));
 sky130_fd_sc_hd__o21ai_0 _37389_ (.A1(net2860),
    .A2(net1270),
    .B1(_16129_),
    .Y(_16130_));
 sky130_fd_sc_hd__nand2_1 _37391_ (.A(net1672),
    .B(net1997),
    .Y(_16132_));
 sky130_fd_sc_hd__o21ai_0 _37392_ (.A1(net1997),
    .A2(net1349),
    .B1(_16132_),
    .Y(_16133_));
 sky130_fd_sc_hd__mux2i_1 _37394_ (.A0(_16130_),
    .A1(_16133_),
    .S(net1689),
    .Y(_16135_));
 sky130_fd_sc_hd__nand2_1 _37395_ (.A(net1117),
    .B(net1998),
    .Y(_16136_));
 sky130_fd_sc_hd__o21ai_0 _37396_ (.A1(net1997),
    .A2(net1360),
    .B1(_16136_),
    .Y(_16137_));
 sky130_fd_sc_hd__nand2_1 _37397_ (.A(net1669),
    .B(net1997),
    .Y(_16138_));
 sky130_fd_sc_hd__o21ai_0 _37398_ (.A1(net1997),
    .A2(net1354),
    .B1(_16138_),
    .Y(_16139_));
 sky130_fd_sc_hd__mux2i_1 _37399_ (.A0(_16137_),
    .A1(_16139_),
    .S(net1251),
    .Y(_16140_));
 sky130_fd_sc_hd__mux2i_1 _37401_ (.A0(_16135_),
    .A1(_16140_),
    .S(net1702),
    .Y(_16142_));
 sky130_fd_sc_hd__nand2_1 _37402_ (.A(net1708),
    .B(net2860),
    .Y(_16143_));
 sky130_fd_sc_hd__o21ai_0 _37403_ (.A1(net2859),
    .A2(net1476),
    .B1(_16143_),
    .Y(_16144_));
 sky130_fd_sc_hd__nor2_1 _37404_ (.A(net1997),
    .B(_03082_),
    .Y(_16145_));
 sky130_fd_sc_hd__o21ai_0 _37405_ (.A1(net2859),
    .A2(net1481),
    .B1(net1687),
    .Y(_16146_));
 sky130_fd_sc_hd__o221ai_1 _37406_ (.A1(net1687),
    .A2(_16144_),
    .B1(_16145_),
    .B2(_16146_),
    .C1(net1704),
    .Y(_16147_));
 sky130_fd_sc_hd__nand2_1 _37408_ (.A(net1466),
    .B(net1997),
    .Y(_16149_));
 sky130_fd_sc_hd__o21ai_0 _37409_ (.A1(net1997),
    .A2(net1368),
    .B1(_16149_),
    .Y(_16150_));
 sky130_fd_sc_hd__nand2_1 _37410_ (.A(net1736),
    .B(net1997),
    .Y(_16151_));
 sky130_fd_sc_hd__o21ai_0 _37411_ (.A1(net1997),
    .A2(net1365),
    .B1(_16151_),
    .Y(_16152_));
 sky130_fd_sc_hd__nand2_1 _37412_ (.A(_16152_),
    .B(net1251),
    .Y(_16153_));
 sky130_fd_sc_hd__o21ai_0 _37413_ (.A1(net1251),
    .A2(_16150_),
    .B1(_16153_),
    .Y(_16154_));
 sky130_fd_sc_hd__nand2_1 _37414_ (.A(_16154_),
    .B(net1384),
    .Y(_16155_));
 sky130_fd_sc_hd__a31oi_1 _37416_ (.A1(_16147_),
    .A2(net1189),
    .A3(_16155_),
    .B1(net1391),
    .Y(_16157_));
 sky130_fd_sc_hd__o21ai_0 _37417_ (.A1(net1187),
    .A2(_16142_),
    .B1(_16157_),
    .Y(_16158_));
 sky130_fd_sc_hd__nand2_1 _37418_ (.A(net1677),
    .B(net1998),
    .Y(_16159_));
 sky130_fd_sc_hd__o21ai_0 _37419_ (.A1(net1998),
    .A2(net1334),
    .B1(_16159_),
    .Y(_16160_));
 sky130_fd_sc_hd__nand2_1 _37420_ (.A(_05903_),
    .B(net2859),
    .Y(_16161_));
 sky130_fd_sc_hd__o21a_1 _37421_ (.A1(net2859),
    .A2(net1273),
    .B1(_16161_),
    .X(_16162_));
 sky130_fd_sc_hd__nand2_1 _37422_ (.A(_16162_),
    .B(net1687),
    .Y(_16163_));
 sky130_fd_sc_hd__o21ai_0 _37423_ (.A1(net1687),
    .A2(_16160_),
    .B1(_16163_),
    .Y(_16164_));
 sky130_fd_sc_hd__nand2_1 _37424_ (.A(_16164_),
    .B(net1702),
    .Y(_16165_));
 sky130_fd_sc_hd__nand2_1 _37425_ (.A(net1129),
    .B(net1998),
    .Y(_16166_));
 sky130_fd_sc_hd__o21ai_0 _37426_ (.A1(net1998),
    .A2(net1325),
    .B1(_16166_),
    .Y(_16167_));
 sky130_fd_sc_hd__nand2_1 _37427_ (.A(net1126),
    .B(net1998),
    .Y(_16168_));
 sky130_fd_sc_hd__o21ai_0 _37428_ (.A1(net1998),
    .A2(net1329),
    .B1(_16168_),
    .Y(_16169_));
 sky130_fd_sc_hd__mux2i_1 _37429_ (.A0(_16167_),
    .A1(_16169_),
    .S(net1688),
    .Y(_16170_));
 sky130_fd_sc_hd__nand2_1 _37430_ (.A(_16170_),
    .B(net1384),
    .Y(_16171_));
 sky130_fd_sc_hd__nand2_1 _37431_ (.A(_16165_),
    .B(_16171_),
    .Y(_16172_));
 sky130_fd_sc_hd__nand2_1 _37432_ (.A(net1141),
    .B(net1999),
    .Y(_16173_));
 sky130_fd_sc_hd__o21ai_0 _37433_ (.A1(net1999),
    .A2(net1306),
    .B1(_16173_),
    .Y(_16174_));
 sky130_fd_sc_hd__nand2_1 _37434_ (.A(net1146),
    .B(net2859),
    .Y(_16175_));
 sky130_fd_sc_hd__o21ai_0 _37435_ (.A1(net2859),
    .A2(net1296),
    .B1(_16175_),
    .Y(_16176_));
 sky130_fd_sc_hd__mux2i_1 _37436_ (.A0(_16174_),
    .A1(_16176_),
    .S(net1688),
    .Y(_16177_));
 sky130_fd_sc_hd__nand2_1 _37437_ (.A(net1151),
    .B(net2859),
    .Y(_16178_));
 sky130_fd_sc_hd__o21ai_0 _37438_ (.A1(net2859),
    .A2(net1287),
    .B1(_16178_),
    .Y(_16179_));
 sky130_fd_sc_hd__nand2_1 _37439_ (.A(_16179_),
    .B(net1688),
    .Y(_16180_));
 sky130_fd_sc_hd__nand2_1 _37440_ (.A(net1148),
    .B(net2859),
    .Y(_16181_));
 sky130_fd_sc_hd__o21ai_0 _37441_ (.A1(net2859),
    .A2(net1292),
    .B1(_16181_),
    .Y(_16182_));
 sky130_fd_sc_hd__nand2_1 _37442_ (.A(_16182_),
    .B(net1250),
    .Y(_16183_));
 sky130_fd_sc_hd__nand2_1 _37443_ (.A(_16180_),
    .B(_16183_),
    .Y(_16184_));
 sky130_fd_sc_hd__nand2_1 _37444_ (.A(_16184_),
    .B(net1703),
    .Y(_16185_));
 sky130_fd_sc_hd__o21ai_0 _37445_ (.A1(net1703),
    .A2(_16177_),
    .B1(_16185_),
    .Y(_16186_));
 sky130_fd_sc_hd__nand2_1 _37446_ (.A(_16186_),
    .B(net1387),
    .Y(_16187_));
 sky130_fd_sc_hd__o21ai_0 _37447_ (.A1(net1387),
    .A2(_16172_),
    .B1(_16187_),
    .Y(_16188_));
 sky130_fd_sc_hd__nand2_1 _37448_ (.A(_16188_),
    .B(net1391),
    .Y(_16189_));
 sky130_fd_sc_hd__nand3_1 _37449_ (.A(_16158_),
    .B(net1200),
    .C(_16189_),
    .Y(_16190_));
 sky130_fd_sc_hd__nand3_1 _37450_ (.A(_16127_),
    .B(net2297),
    .C(_16190_),
    .Y(_16191_));
 sky130_fd_sc_hd__o211ai_1 _37451_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[0] ),
    .A2(net2297),
    .B1(net2183),
    .C1(_16191_),
    .Y(_16192_));
 sky130_fd_sc_hd__inv_2 _37452_ (.A(_16192_),
    .Y(_04453_));
 sky130_fd_sc_hd__nand2_1 _37453_ (.A(_16115_),
    .B(net1383),
    .Y(_16193_));
 sky130_fd_sc_hd__o21ai_0 _37454_ (.A1(net1383),
    .A2(_16106_),
    .B1(_16193_),
    .Y(_16194_));
 sky130_fd_sc_hd__nand2_1 _37455_ (.A(_16120_),
    .B(net1700),
    .Y(_16195_));
 sky130_fd_sc_hd__o21ai_0 _37456_ (.A1(net1700),
    .A2(_16091_),
    .B1(_16195_),
    .Y(_16196_));
 sky130_fd_sc_hd__nand2_1 _37457_ (.A(_16196_),
    .B(net1388),
    .Y(_16197_));
 sky130_fd_sc_hd__o21ai_0 _37458_ (.A1(net1388),
    .A2(_16194_),
    .B1(_16197_),
    .Y(_16198_));
 sky130_fd_sc_hd__nor2_1 _37459_ (.A(net1177),
    .B(_16198_),
    .Y(_16199_));
 sky130_fd_sc_hd__mux2i_1 _37460_ (.A0(_16101_),
    .A1(_16177_),
    .S(net1703),
    .Y(_16200_));
 sky130_fd_sc_hd__nand2_1 _37461_ (.A(_16170_),
    .B(net1702),
    .Y(_16201_));
 sky130_fd_sc_hd__o21ai_0 _37462_ (.A1(net1703),
    .A2(_16184_),
    .B1(_16201_),
    .Y(_16202_));
 sky130_fd_sc_hd__nand2_1 _37463_ (.A(_16202_),
    .B(net1186),
    .Y(_16203_));
 sky130_fd_sc_hd__o21ai_0 _37464_ (.A1(net1186),
    .A2(_16200_),
    .B1(_16203_),
    .Y(_16204_));
 sky130_fd_sc_hd__o21ai_0 _37465_ (.A1(net1390),
    .A2(_16204_),
    .B1(net1199),
    .Y(_16205_));
 sky130_fd_sc_hd__nand2_1 _37468_ (.A(net2857),
    .B(\inst$top.soc.cpu.d.sink__payload.sext ),
    .Y(_16208_));
 sky130_fd_sc_hd__nor2_1 _37469_ (.A(_16208_),
    .B(net1221),
    .Y(_16209_));
 sky130_fd_sc_hd__nand2_1 _37470_ (.A(_16209_),
    .B(net1382),
    .Y(_16210_));
 sky130_fd_sc_hd__o21ai_0 _37471_ (.A1(net1382),
    .A2(_16077_),
    .B1(_16210_),
    .Y(_16211_));
 sky130_fd_sc_hd__nand2_1 _37472_ (.A(_16068_),
    .B(net1382),
    .Y(_16212_));
 sky130_fd_sc_hd__o21ai_0 _37473_ (.A1(net1382),
    .A2(_16085_),
    .B1(_16212_),
    .Y(_16213_));
 sky130_fd_sc_hd__nand2_1 _37474_ (.A(_16213_),
    .B(net1185),
    .Y(_16214_));
 sky130_fd_sc_hd__o21ai_0 _37475_ (.A1(net1185),
    .A2(_16211_),
    .B1(_16214_),
    .Y(_16215_));
 sky130_fd_sc_hd__inv_1 _37476_ (.A(_16209_),
    .Y(_16216_));
 sky130_fd_sc_hd__nor2_1 _37477_ (.A(net1177),
    .B(_16216_),
    .Y(_16217_));
 sky130_fd_sc_hd__inv_1 _37478_ (.A(_16217_),
    .Y(_16218_));
 sky130_fd_sc_hd__o21ai_0 _37479_ (.A1(net1390),
    .A2(_16215_),
    .B1(_16218_),
    .Y(_16219_));
 sky130_fd_sc_hd__nand2_1 _37481_ (.A(_16219_),
    .B(net1072),
    .Y(_16221_));
 sky130_fd_sc_hd__o211ai_1 _37482_ (.A1(_16199_),
    .A2(_16205_),
    .B1(net2296),
    .C1(_16221_),
    .Y(_16222_));
 sky130_fd_sc_hd__o211ai_1 _37483_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[10] ),
    .A2(net2293),
    .B1(net2181),
    .C1(_16222_),
    .Y(_16223_));
 sky130_fd_sc_hd__inv_2 _37484_ (.A(_16223_),
    .Y(_04454_));
 sky130_fd_sc_hd__nand2_1 _37485_ (.A(_16089_),
    .B(net1685),
    .Y(_16224_));
 sky130_fd_sc_hd__o21ai_0 _37486_ (.A1(net1685),
    .A2(_16083_),
    .B1(_16224_),
    .Y(_16225_));
 sky130_fd_sc_hd__nand2_1 _37487_ (.A(_16225_),
    .B(net1383),
    .Y(_16226_));
 sky130_fd_sc_hd__nand2_1 _37488_ (.A(_16117_),
    .B(net1685),
    .Y(_16227_));
 sky130_fd_sc_hd__o21ai_0 _37489_ (.A1(net1685),
    .A2(_16087_),
    .B1(_16227_),
    .Y(_16228_));
 sky130_fd_sc_hd__nand2_1 _37490_ (.A(_16228_),
    .B(net1700),
    .Y(_16229_));
 sky130_fd_sc_hd__nand2_1 _37491_ (.A(_16226_),
    .B(_16229_),
    .Y(_16230_));
 sky130_fd_sc_hd__or2_2 _37492_ (.A(net1685),
    .B(_16119_),
    .X(_16231_));
 sky130_fd_sc_hd__o21ai_0 _37493_ (.A1(net1250),
    .A2(_16113_),
    .B1(_16231_),
    .Y(_16232_));
 sky130_fd_sc_hd__nand2_1 _37494_ (.A(_16232_),
    .B(net1383),
    .Y(_16233_));
 sky130_fd_sc_hd__mux2i_1 _37495_ (.A0(_16103_),
    .A1(_16110_),
    .S(net1250),
    .Y(_16234_));
 sky130_fd_sc_hd__nand2_1 _37496_ (.A(_16234_),
    .B(net1700),
    .Y(_16235_));
 sky130_fd_sc_hd__nand2_1 _37497_ (.A(_16233_),
    .B(_16235_),
    .Y(_16236_));
 sky130_fd_sc_hd__nand2_1 _37498_ (.A(_16236_),
    .B(net1184),
    .Y(_16237_));
 sky130_fd_sc_hd__o21ai_0 _37499_ (.A1(net1184),
    .A2(_16230_),
    .B1(_16237_),
    .Y(_16238_));
 sky130_fd_sc_hd__nor2_1 _37500_ (.A(net1175),
    .B(_16238_),
    .Y(_16239_));
 sky130_fd_sc_hd__mux2i_1 _37501_ (.A0(_16105_),
    .A1(_16098_),
    .S(net1688),
    .Y(_16240_));
 sky130_fd_sc_hd__mux2i_1 _37502_ (.A0(_16100_),
    .A1(_16174_),
    .S(net1688),
    .Y(_16241_));
 sky130_fd_sc_hd__inv_1 _37503_ (.A(_16241_),
    .Y(_16242_));
 sky130_fd_sc_hd__nand2_1 _37504_ (.A(_16242_),
    .B(net1703),
    .Y(_16243_));
 sky130_fd_sc_hd__o21ai_0 _37505_ (.A1(net1700),
    .A2(_16240_),
    .B1(_16243_),
    .Y(_16244_));
 sky130_fd_sc_hd__mux2i_1 _37506_ (.A0(_16176_),
    .A1(_16182_),
    .S(net1688),
    .Y(_16245_));
 sky130_fd_sc_hd__nand2_1 _37507_ (.A(_16245_),
    .B(net1384),
    .Y(_16246_));
 sky130_fd_sc_hd__mux2i_1 _37508_ (.A0(_16179_),
    .A1(_16167_),
    .S(net1688),
    .Y(_16247_));
 sky130_fd_sc_hd__nand2_1 _37509_ (.A(_16247_),
    .B(net1702),
    .Y(_16248_));
 sky130_fd_sc_hd__nand2_1 _37510_ (.A(_16246_),
    .B(_16248_),
    .Y(_16249_));
 sky130_fd_sc_hd__nand2_1 _37511_ (.A(_16249_),
    .B(net1186),
    .Y(_16250_));
 sky130_fd_sc_hd__o21ai_0 _37512_ (.A1(net1186),
    .A2(_16244_),
    .B1(_16250_),
    .Y(_16251_));
 sky130_fd_sc_hd__o21ai_0 _37513_ (.A1(net1391),
    .A2(_16251_),
    .B1(net1200),
    .Y(_16252_));
 sky130_fd_sc_hd__o21ai_0 _37514_ (.A1(net1686),
    .A2(_16209_),
    .B1(_16073_),
    .Y(_16253_));
 sky130_fd_sc_hd__o21ai_0 _37515_ (.A1(net1382),
    .A2(_16253_),
    .B1(_16210_),
    .Y(_16254_));
 sky130_fd_sc_hd__mux2i_1 _37516_ (.A0(_16066_),
    .A1(_16081_),
    .S(net1686),
    .Y(_16255_));
 sky130_fd_sc_hd__nand2_1 _37517_ (.A(_16075_),
    .B(net1250),
    .Y(_16256_));
 sky130_fd_sc_hd__o21ai_0 _37518_ (.A1(net1250),
    .A2(_16064_),
    .B1(_16256_),
    .Y(_16257_));
 sky130_fd_sc_hd__nand2_1 _37519_ (.A(_16257_),
    .B(net1382),
    .Y(_16258_));
 sky130_fd_sc_hd__o21ai_0 _37520_ (.A1(net1382),
    .A2(_16255_),
    .B1(_16258_),
    .Y(_16259_));
 sky130_fd_sc_hd__nand2_1 _37521_ (.A(_16259_),
    .B(net1184),
    .Y(_16260_));
 sky130_fd_sc_hd__o21ai_0 _37522_ (.A1(net1184),
    .A2(_16254_),
    .B1(_16260_),
    .Y(_16261_));
 sky130_fd_sc_hd__o21ai_0 _37523_ (.A1(net1392),
    .A2(_16261_),
    .B1(_16218_),
    .Y(_16262_));
 sky130_fd_sc_hd__nand2_1 _37524_ (.A(_16262_),
    .B(net1074),
    .Y(_16263_));
 sky130_fd_sc_hd__o211ai_1 _37525_ (.A1(_16239_),
    .A2(_16252_),
    .B1(net2296),
    .C1(_16263_),
    .Y(_16264_));
 sky130_fd_sc_hd__o211ai_1 _37526_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[11] ),
    .A2(net2295),
    .B1(net2181),
    .C1(_16264_),
    .Y(_16265_));
 sky130_fd_sc_hd__inv_2 _37527_ (.A(_16265_),
    .Y(_04455_));
 sky130_fd_sc_hd__nand2_1 _37529_ (.A(_16122_),
    .B(net1185),
    .Y(_16267_));
 sky130_fd_sc_hd__o21ai_0 _37530_ (.A1(net1185),
    .A2(_16093_),
    .B1(_16267_),
    .Y(_16268_));
 sky130_fd_sc_hd__mux2i_1 _37531_ (.A0(_16108_),
    .A1(_16186_),
    .S(net1185),
    .Y(_16269_));
 sky130_fd_sc_hd__o21ai_0 _37532_ (.A1(net1391),
    .A2(_16269_),
    .B1(net1198),
    .Y(_16270_));
 sky130_fd_sc_hd__o21bai_1 _37533_ (.A1(net1175),
    .A2(_16268_),
    .B1_N(_16270_),
    .Y(_16271_));
 sky130_fd_sc_hd__nand3_1 _37534_ (.A(_16069_),
    .B(_16079_),
    .C(net1185),
    .Y(_16272_));
 sky130_fd_sc_hd__nor2_1 _37535_ (.A(net1185),
    .B(_16216_),
    .Y(_16273_));
 sky130_fd_sc_hd__inv_1 _37536_ (.A(_16273_),
    .Y(_16274_));
 sky130_fd_sc_hd__nand2_1 _37537_ (.A(_16272_),
    .B(_16274_),
    .Y(_16275_));
 sky130_fd_sc_hd__inv_1 _37538_ (.A(_16275_),
    .Y(_16276_));
 sky130_fd_sc_hd__o21ai_0 _37539_ (.A1(net1390),
    .A2(_16276_),
    .B1(_16218_),
    .Y(_16277_));
 sky130_fd_sc_hd__nand2_1 _37540_ (.A(_16277_),
    .B(net1074),
    .Y(_16278_));
 sky130_fd_sc_hd__o21ai_0 _37541_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[12] ),
    .A2(net2295),
    .B1(net2183),
    .Y(_16279_));
 sky130_fd_sc_hd__a31oi_1 _37542_ (.A1(_16271_),
    .A2(_16278_),
    .A3(net2295),
    .B1(_16279_),
    .Y(_04456_));
 sky130_fd_sc_hd__nand2_1 _37543_ (.A(_16228_),
    .B(net1383),
    .Y(_16280_));
 sky130_fd_sc_hd__o21a_1 _37544_ (.A1(net1383),
    .A2(_16232_),
    .B1(_16280_),
    .X(_16281_));
 sky130_fd_sc_hd__nand2_1 _37545_ (.A(_16281_),
    .B(net1184),
    .Y(_16282_));
 sky130_fd_sc_hd__nand2_1 _37546_ (.A(_16255_),
    .B(net1383),
    .Y(_16283_));
 sky130_fd_sc_hd__o21ai_0 _37547_ (.A1(net1383),
    .A2(_16225_),
    .B1(_16283_),
    .Y(_16284_));
 sky130_fd_sc_hd__nand2_1 _37548_ (.A(_16284_),
    .B(net1386),
    .Y(_16285_));
 sky130_fd_sc_hd__nand2_1 _37549_ (.A(_16282_),
    .B(_16285_),
    .Y(_16286_));
 sky130_fd_sc_hd__nand2_1 _37550_ (.A(_16242_),
    .B(net1384),
    .Y(_16287_));
 sky130_fd_sc_hd__o21ai_0 _37551_ (.A1(net1384),
    .A2(_16245_),
    .B1(_16287_),
    .Y(_16288_));
 sky130_fd_sc_hd__nand2_1 _37552_ (.A(_16288_),
    .B(net1186),
    .Y(_16289_));
 sky130_fd_sc_hd__mux2i_1 _37553_ (.A0(_16240_),
    .A1(_16234_),
    .S(net1384),
    .Y(_16290_));
 sky130_fd_sc_hd__nand2_1 _37554_ (.A(_16290_),
    .B(net1387),
    .Y(_16291_));
 sky130_fd_sc_hd__nand2_1 _37555_ (.A(_16289_),
    .B(_16291_),
    .Y(_16292_));
 sky130_fd_sc_hd__nand2_1 _37556_ (.A(_16292_),
    .B(net1178),
    .Y(_16293_));
 sky130_fd_sc_hd__o211ai_1 _37557_ (.A1(net1178),
    .A2(_16286_),
    .B1(net1200),
    .C1(_16293_),
    .Y(_16294_));
 sky130_fd_sc_hd__nand2_1 _37558_ (.A(_16257_),
    .B(net1701),
    .Y(_16295_));
 sky130_fd_sc_hd__nand2_1 _37559_ (.A(_16253_),
    .B(net1382),
    .Y(_16296_));
 sky130_fd_sc_hd__nand2_1 _37560_ (.A(_16295_),
    .B(_16296_),
    .Y(_16297_));
 sky130_fd_sc_hd__o21ai_0 _37561_ (.A1(net1388),
    .A2(_16297_),
    .B1(_16274_),
    .Y(_16298_));
 sky130_fd_sc_hd__nand2_1 _37562_ (.A(_16298_),
    .B(net1175),
    .Y(_16299_));
 sky130_fd_sc_hd__nand2_1 _37563_ (.A(_16299_),
    .B(_16218_),
    .Y(_16300_));
 sky130_fd_sc_hd__nand2_1 _37564_ (.A(_16300_),
    .B(net1073),
    .Y(_16301_));
 sky130_fd_sc_hd__nand3_1 _37565_ (.A(_16294_),
    .B(net2297),
    .C(_16301_),
    .Y(_16302_));
 sky130_fd_sc_hd__o211ai_1 _37566_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[13] ),
    .A2(net2293),
    .B1(net2181),
    .C1(_16302_),
    .Y(_16303_));
 sky130_fd_sc_hd__inv_2 _37567_ (.A(_16303_),
    .Y(_04457_));
 sky130_fd_sc_hd__a21oi_1 _37568_ (.A1(_16211_),
    .A2(net1185),
    .B1(_16273_),
    .Y(_16304_));
 sky130_fd_sc_hd__inv_1 _37569_ (.A(_16304_),
    .Y(_16305_));
 sky130_fd_sc_hd__a21oi_1 _37570_ (.A1(_16305_),
    .A2(net1177),
    .B1(_16217_),
    .Y(_16306_));
 sky130_fd_sc_hd__nand2_1 _37571_ (.A(_16213_),
    .B(net1388),
    .Y(_16307_));
 sky130_fd_sc_hd__o21ai_0 _37572_ (.A1(net1388),
    .A2(_16196_),
    .B1(_16307_),
    .Y(_16308_));
 sky130_fd_sc_hd__nand2_1 _37573_ (.A(_16308_),
    .B(net1390),
    .Y(_16309_));
 sky130_fd_sc_hd__nand2_1 _37574_ (.A(_16200_),
    .B(net1184),
    .Y(_16310_));
 sky130_fd_sc_hd__nand2_1 _37575_ (.A(_16194_),
    .B(net1386),
    .Y(_16311_));
 sky130_fd_sc_hd__nand2_1 _37576_ (.A(_16310_),
    .B(_16311_),
    .Y(_16312_));
 sky130_fd_sc_hd__nand2_1 _37577_ (.A(_16312_),
    .B(net1176),
    .Y(_16313_));
 sky130_fd_sc_hd__nand3_1 _37578_ (.A(_16309_),
    .B(net1198),
    .C(_16313_),
    .Y(_16314_));
 sky130_fd_sc_hd__o21ai_0 _37579_ (.A1(net1198),
    .A2(_16306_),
    .B1(_16314_),
    .Y(_16315_));
 sky130_fd_sc_hd__nor2_1 _37580_ (.A(\inst$top.soc.cpu.shifter.m_result$7[14] ),
    .B(net2295),
    .Y(_16316_));
 sky130_fd_sc_hd__nor2_1 _37581_ (.A(net3011),
    .B(_16316_),
    .Y(_16317_));
 sky130_fd_sc_hd__o21ai_0 _37582_ (.A1(net1926),
    .A2(_16315_),
    .B1(_16317_),
    .Y(_16318_));
 sky130_fd_sc_hd__inv_2 _37583_ (.A(_16318_),
    .Y(_04458_));
 sky130_fd_sc_hd__nand2_1 _37584_ (.A(_16244_),
    .B(net1184),
    .Y(_16319_));
 sky130_fd_sc_hd__o21ai_0 _37585_ (.A1(net1184),
    .A2(_16236_),
    .B1(_16319_),
    .Y(_16320_));
 sky130_fd_sc_hd__nand2_1 _37586_ (.A(_16320_),
    .B(net1176),
    .Y(_16321_));
 sky130_fd_sc_hd__nor2_1 _37587_ (.A(net1184),
    .B(_16259_),
    .Y(_16322_));
 sky130_fd_sc_hd__a31oi_1 _37588_ (.A1(net1184),
    .A2(_16229_),
    .A3(_16226_),
    .B1(_16322_),
    .Y(_16323_));
 sky130_fd_sc_hd__nand2_1 _37589_ (.A(_16323_),
    .B(net1390),
    .Y(_16324_));
 sky130_fd_sc_hd__nand3_1 _37590_ (.A(_16321_),
    .B(net1198),
    .C(_16324_),
    .Y(_16325_));
 sky130_fd_sc_hd__a21oi_1 _37591_ (.A1(_16254_),
    .A2(net1185),
    .B1(_16273_),
    .Y(_16326_));
 sky130_fd_sc_hd__o21ai_0 _37592_ (.A1(net1390),
    .A2(_16326_),
    .B1(_16218_),
    .Y(_16327_));
 sky130_fd_sc_hd__nand2_1 _37593_ (.A(_16327_),
    .B(net1072),
    .Y(_16328_));
 sky130_fd_sc_hd__nand3_1 _37594_ (.A(_16325_),
    .B(net2296),
    .C(_16328_),
    .Y(_16329_));
 sky130_fd_sc_hd__o211ai_1 _37595_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[15] ),
    .A2(net2296),
    .B1(net2183),
    .C1(_16329_),
    .Y(_16330_));
 sky130_fd_sc_hd__inv_2 _37596_ (.A(_16330_),
    .Y(_04459_));
 sky130_fd_sc_hd__nand2_1 _37598_ (.A(_16126_),
    .B(net1200),
    .Y(_16332_));
 sky130_fd_sc_hd__o21ai_1 _37599_ (.A1(net1198),
    .A2(_16216_),
    .B1(net2296),
    .Y(_16333_));
 sky130_fd_sc_hd__inv_2 _37600_ (.A(_16333_),
    .Y(_16334_));
 sky130_fd_sc_hd__a221oi_2 _37602_ (.A1(_13404_),
    .A2(net1918),
    .B1(_16332_),
    .B2(_16334_),
    .C1(net3006),
    .Y(_04460_));
 sky130_fd_sc_hd__nand2_1 _37603_ (.A(_16297_),
    .B(net1386),
    .Y(_16336_));
 sky130_fd_sc_hd__o21ai_0 _37604_ (.A1(net1386),
    .A2(_16284_),
    .B1(_16336_),
    .Y(_16337_));
 sky130_fd_sc_hd__nand2_1 _37605_ (.A(_16281_),
    .B(net1386),
    .Y(_16338_));
 sky130_fd_sc_hd__o21ai_0 _37606_ (.A1(net1386),
    .A2(_16290_),
    .B1(_16338_),
    .Y(_16339_));
 sky130_fd_sc_hd__nand2_1 _37607_ (.A(_16339_),
    .B(net1176),
    .Y(_16340_));
 sky130_fd_sc_hd__o21ai_0 _37608_ (.A1(net1175),
    .A2(_16337_),
    .B1(_16340_),
    .Y(_16341_));
 sky130_fd_sc_hd__nand2_1 _37609_ (.A(_16341_),
    .B(net1199),
    .Y(_16342_));
 sky130_fd_sc_hd__o21ai_0 _37610_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[17] ),
    .A2(net2295),
    .B1(net2183),
    .Y(_16343_));
 sky130_fd_sc_hd__a21oi_1 _37611_ (.A1(_16342_),
    .A2(_16334_),
    .B1(_16343_),
    .Y(_04461_));
 sky130_fd_sc_hd__nand2_1 _37612_ (.A(_16198_),
    .B(net1177),
    .Y(_16344_));
 sky130_fd_sc_hd__o21ai_0 _37613_ (.A1(net1177),
    .A2(_16215_),
    .B1(_16344_),
    .Y(_16345_));
 sky130_fd_sc_hd__nand2_1 _37614_ (.A(_16345_),
    .B(net1202),
    .Y(_16346_));
 sky130_fd_sc_hd__a221oi_2 _37615_ (.A1(_13578_),
    .A2(net1924),
    .B1(_16346_),
    .B2(_16334_),
    .C1(net3005),
    .Y(_04462_));
 sky130_fd_sc_hd__nand2_1 _37616_ (.A(_16238_),
    .B(net1175),
    .Y(_16347_));
 sky130_fd_sc_hd__o21ai_0 _37617_ (.A1(net1175),
    .A2(_16261_),
    .B1(_16347_),
    .Y(_16348_));
 sky130_fd_sc_hd__nand2_1 _37618_ (.A(_16348_),
    .B(net1202),
    .Y(_16349_));
 sky130_fd_sc_hd__a221oi_2 _37619_ (.A1(_13596_),
    .A2(net1924),
    .B1(_16349_),
    .B2(_16334_),
    .C1(net3010),
    .Y(_04463_));
 sky130_fd_sc_hd__nand2_1 _37620_ (.A(_16341_),
    .B(net1073),
    .Y(_16350_));
 sky130_fd_sc_hd__mux2i_1 _37621_ (.A0(_16160_),
    .A1(_16169_),
    .S(net1250),
    .Y(_16351_));
 sky130_fd_sc_hd__nand2_1 _37622_ (.A(_16351_),
    .B(net1702),
    .Y(_16352_));
 sky130_fd_sc_hd__nand2_1 _37623_ (.A(_16247_),
    .B(net1384),
    .Y(_16353_));
 sky130_fd_sc_hd__nand2_1 _37624_ (.A(_16352_),
    .B(_16353_),
    .Y(_16354_));
 sky130_fd_sc_hd__nand2_1 _37625_ (.A(_16288_),
    .B(net1387),
    .Y(_16355_));
 sky130_fd_sc_hd__o21ai_0 _37626_ (.A1(net1386),
    .A2(_16354_),
    .B1(_16355_),
    .Y(_16356_));
 sky130_fd_sc_hd__nand2_1 _37627_ (.A(_16356_),
    .B(net1391),
    .Y(_16357_));
 sky130_fd_sc_hd__nand2_1 _37628_ (.A(_16130_),
    .B(net1687),
    .Y(_16358_));
 sky130_fd_sc_hd__o21ai_0 _37629_ (.A1(net1687),
    .A2(_16162_),
    .B1(_16358_),
    .Y(_16359_));
 sky130_fd_sc_hd__mux2i_1 _37630_ (.A0(_16133_),
    .A1(_16139_),
    .S(net1687),
    .Y(_16360_));
 sky130_fd_sc_hd__nand2_1 _37631_ (.A(_16360_),
    .B(net1704),
    .Y(_16361_));
 sky130_fd_sc_hd__o21ai_0 _37632_ (.A1(net1704),
    .A2(_16359_),
    .B1(_16361_),
    .Y(_16362_));
 sky130_fd_sc_hd__inv_1 _37633_ (.A(_16362_),
    .Y(_16363_));
 sky130_fd_sc_hd__nand2_1 _37634_ (.A(_16152_),
    .B(net1687),
    .Y(_16364_));
 sky130_fd_sc_hd__nand2_1 _37635_ (.A(_16137_),
    .B(net1250),
    .Y(_16365_));
 sky130_fd_sc_hd__nand2_1 _37636_ (.A(_16364_),
    .B(_16365_),
    .Y(_16366_));
 sky130_fd_sc_hd__nor2_1 _37637_ (.A(net1704),
    .B(_16366_),
    .Y(_16367_));
 sky130_fd_sc_hd__o21ai_0 _37638_ (.A1(net1687),
    .A2(_16150_),
    .B1(net1704),
    .Y(_16368_));
 sky130_fd_sc_hd__a21oi_1 _37639_ (.A1(net1687),
    .A2(_16144_),
    .B1(_16368_),
    .Y(_16369_));
 sky130_fd_sc_hd__o21ai_0 _37640_ (.A1(_16367_),
    .A2(_16369_),
    .B1(net1188),
    .Y(_16370_));
 sky130_fd_sc_hd__o211ai_1 _37641_ (.A1(net1188),
    .A2(_16363_),
    .B1(net1179),
    .C1(_16370_),
    .Y(_16371_));
 sky130_fd_sc_hd__nand3_1 _37642_ (.A(_16357_),
    .B(net1200),
    .C(_16371_),
    .Y(_16372_));
 sky130_fd_sc_hd__nand3_1 _37643_ (.A(_16350_),
    .B(net2298),
    .C(_16372_),
    .Y(_16373_));
 sky130_fd_sc_hd__o211ai_1 _37644_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[1] ),
    .A2(net2297),
    .B1(net2183),
    .C1(_16373_),
    .Y(_16374_));
 sky130_fd_sc_hd__inv_2 _37645_ (.A(_16374_),
    .Y(_04464_));
 sky130_fd_sc_hd__nand2_1 _37648_ (.A(_16276_),
    .B(net1390),
    .Y(_16377_));
 sky130_fd_sc_hd__o21ai_0 _37649_ (.A1(net1390),
    .A2(_16268_),
    .B1(_16377_),
    .Y(_16378_));
 sky130_fd_sc_hd__o21ai_0 _37650_ (.A1(net1076),
    .A2(_16378_),
    .B1(_16334_),
    .Y(_16379_));
 sky130_fd_sc_hd__o211a_1 _37651_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[20] ),
    .A2(net2294),
    .B1(net2182),
    .C1(_16379_),
    .X(_16380_));
 sky130_fd_sc_hd__nand3_1 _37653_ (.A(_16282_),
    .B(net1176),
    .C(_16285_),
    .Y(_16381_));
 sky130_fd_sc_hd__o21ai_0 _37654_ (.A1(net1176),
    .A2(_16298_),
    .B1(_16381_),
    .Y(_16382_));
 sky130_fd_sc_hd__nor2_1 _37655_ (.A(net1073),
    .B(_16382_),
    .Y(_16383_));
 sky130_fd_sc_hd__o221a_2 _37656_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[21] ),
    .A2(net2297),
    .B1(_16333_),
    .B2(_16383_),
    .C1(net2183),
    .X(_16384_));
 sky130_fd_sc_hd__nand2_1 _37658_ (.A(_16308_),
    .B(net1177),
    .Y(_16385_));
 sky130_fd_sc_hd__o21ai_0 _37659_ (.A1(net1177),
    .A2(_16305_),
    .B1(_16385_),
    .Y(_16386_));
 sky130_fd_sc_hd__o21ai_0 _37660_ (.A1(net1076),
    .A2(_16386_),
    .B1(_16334_),
    .Y(_16387_));
 sky130_fd_sc_hd__o211a_1 _37661_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[22] ),
    .A2(net2294),
    .B1(net2181),
    .C1(_16387_),
    .X(_16388_));
 sky130_fd_sc_hd__nand2_1 _37663_ (.A(_16323_),
    .B(net1175),
    .Y(_16389_));
 sky130_fd_sc_hd__nand2_1 _37664_ (.A(_16326_),
    .B(net1390),
    .Y(_16390_));
 sky130_fd_sc_hd__nand3_1 _37665_ (.A(_16389_),
    .B(net1198),
    .C(_16390_),
    .Y(_16391_));
 sky130_fd_sc_hd__a221oi_2 _37666_ (.A1(_13903_),
    .A2(net1926),
    .B1(_16391_),
    .B2(_16334_),
    .C1(net3011),
    .Y(_04468_));
 sky130_fd_sc_hd__o21ai_0 _37668_ (.A1(net1391),
    .A2(_16095_),
    .B1(_16218_),
    .Y(_16393_));
 sky130_fd_sc_hd__a21oi_1 _37669_ (.A1(_16393_),
    .A2(net1200),
    .B1(_16333_),
    .Y(_16394_));
 sky130_fd_sc_hd__a211oi_2 _37670_ (.A1(_13952_),
    .A2(net1927),
    .B1(net3011),
    .C1(_16394_),
    .Y(_04469_));
 sky130_fd_sc_hd__o21ai_0 _37671_ (.A1(net1390),
    .A2(_16337_),
    .B1(_16218_),
    .Y(_16395_));
 sky130_fd_sc_hd__a21oi_1 _37672_ (.A1(_16395_),
    .A2(net1199),
    .B1(_16333_),
    .Y(_16396_));
 sky130_fd_sc_hd__a211oi_2 _37673_ (.A1(_14002_),
    .A2(net1925),
    .B1(net3010),
    .C1(_16396_),
    .Y(_04470_));
 sky130_fd_sc_hd__a21oi_1 _37674_ (.A1(_16219_),
    .A2(net1198),
    .B1(_16333_),
    .Y(_16397_));
 sky130_fd_sc_hd__a211oi_2 _37675_ (.A1(_14014_),
    .A2(net1925),
    .B1(net3010),
    .C1(_16397_),
    .Y(_04471_));
 sky130_fd_sc_hd__a21oi_1 _37676_ (.A1(_16262_),
    .A2(net1199),
    .B1(_16333_),
    .Y(_16398_));
 sky130_fd_sc_hd__a211oi_2 _37677_ (.A1(_14068_),
    .A2(net1927),
    .B1(net3011),
    .C1(_16398_),
    .Y(_04472_));
 sky130_fd_sc_hd__a21oi_1 _37679_ (.A1(_16277_),
    .A2(net1198),
    .B1(_16333_),
    .Y(_16400_));
 sky130_fd_sc_hd__a211oi_2 _37680_ (.A1(_14166_),
    .A2(net1926),
    .B1(net3011),
    .C1(_16400_),
    .Y(_04473_));
 sky130_fd_sc_hd__a21oi_1 _37681_ (.A1(_16300_),
    .A2(net1200),
    .B1(_16333_),
    .Y(_16401_));
 sky130_fd_sc_hd__a211oi_2 _37682_ (.A1(_14230_),
    .A2(net1926),
    .B1(net3004),
    .C1(_16401_),
    .Y(_04474_));
 sky130_fd_sc_hd__o21ai_0 _37683_ (.A1(net1702),
    .A2(_16140_),
    .B1(net1188),
    .Y(_16402_));
 sky130_fd_sc_hd__a21oi_1 _37684_ (.A1(net1702),
    .A2(_16154_),
    .B1(_16402_),
    .Y(_16403_));
 sky130_fd_sc_hd__mux2i_1 _37685_ (.A0(_16164_),
    .A1(_16135_),
    .S(net1702),
    .Y(_16404_));
 sky130_fd_sc_hd__o21ai_0 _37686_ (.A1(net1186),
    .A2(_16404_),
    .B1(net1179),
    .Y(_16405_));
 sky130_fd_sc_hd__o221ai_1 _37687_ (.A1(net1179),
    .A2(_16204_),
    .B1(_16403_),
    .B2(_16405_),
    .C1(net1201),
    .Y(_16406_));
 sky130_fd_sc_hd__nand2_1 _37688_ (.A(_16345_),
    .B(net1072),
    .Y(_16407_));
 sky130_fd_sc_hd__nand3_1 _37689_ (.A(_16406_),
    .B(net2296),
    .C(_16407_),
    .Y(_16408_));
 sky130_fd_sc_hd__o211ai_1 _37690_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[2] ),
    .A2(net2295),
    .B1(net2181),
    .C1(_16408_),
    .Y(_16409_));
 sky130_fd_sc_hd__inv_2 _37691_ (.A(_16409_),
    .Y(_04475_));
 sky130_fd_sc_hd__o21ai_0 _37692_ (.A1(net1072),
    .A2(_16306_),
    .B1(_16334_),
    .Y(_16410_));
 sky130_fd_sc_hd__o211a_1 _37693_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[30] ),
    .A2(net2295),
    .B1(net2181),
    .C1(_16410_),
    .X(_16411_));
 sky130_fd_sc_hd__a21oi_1 _37695_ (.A1(_16327_),
    .A2(net1198),
    .B1(_16333_),
    .Y(_16412_));
 sky130_fd_sc_hd__a211oi_2 _37696_ (.A1(_12990_),
    .A2(net1926),
    .B1(net3004),
    .C1(_16412_),
    .Y(_04477_));
 sky130_fd_sc_hd__a21oi_1 _37697_ (.A1(_16364_),
    .A2(_16365_),
    .B1(net1384),
    .Y(_16413_));
 sky130_fd_sc_hd__o21ai_0 _37698_ (.A1(net1704),
    .A2(_16360_),
    .B1(net1188),
    .Y(_16414_));
 sky130_fd_sc_hd__nand2_1 _37699_ (.A(_16359_),
    .B(net1702),
    .Y(_16415_));
 sky130_fd_sc_hd__o21ai_0 _37700_ (.A1(net1702),
    .A2(_16351_),
    .B1(_16415_),
    .Y(_16416_));
 sky130_fd_sc_hd__o221ai_1 _37701_ (.A1(_16413_),
    .A2(_16414_),
    .B1(net1188),
    .B2(_16416_),
    .C1(net1179),
    .Y(_16417_));
 sky130_fd_sc_hd__o211ai_1 _37702_ (.A1(net1178),
    .A2(_16251_),
    .B1(net1200),
    .C1(_16417_),
    .Y(_16418_));
 sky130_fd_sc_hd__nand2_1 _37703_ (.A(_16348_),
    .B(net1072),
    .Y(_16419_));
 sky130_fd_sc_hd__nand3_1 _37704_ (.A(_16418_),
    .B(net2295),
    .C(_16419_),
    .Y(_16420_));
 sky130_fd_sc_hd__o211ai_1 _37705_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[3] ),
    .A2(net2295),
    .B1(net2183),
    .C1(_16420_),
    .Y(_16421_));
 sky130_fd_sc_hd__inv_2 _37706_ (.A(_16421_),
    .Y(_04478_));
 sky130_fd_sc_hd__nand2_1 _37707_ (.A(_16269_),
    .B(net1391),
    .Y(_16422_));
 sky130_fd_sc_hd__a21oi_1 _37708_ (.A1(_16142_),
    .A2(net1187),
    .B1(net1391),
    .Y(_16423_));
 sky130_fd_sc_hd__o21ai_0 _37709_ (.A1(net1187),
    .A2(_16172_),
    .B1(_16423_),
    .Y(_16424_));
 sky130_fd_sc_hd__nand3_1 _37710_ (.A(_16422_),
    .B(net1200),
    .C(_16424_),
    .Y(_16425_));
 sky130_fd_sc_hd__nand2_1 _37711_ (.A(_16378_),
    .B(net1072),
    .Y(_16426_));
 sky130_fd_sc_hd__nand3_1 _37712_ (.A(_16425_),
    .B(_16426_),
    .C(net2295),
    .Y(_16427_));
 sky130_fd_sc_hd__nand2_1 _37713_ (.A(net1926),
    .B(\inst$top.soc.cpu.shifter.m_result$7[4] ),
    .Y(_16428_));
 sky130_fd_sc_hd__a21oi_1 _37714_ (.A1(_16427_),
    .A2(_16428_),
    .B1(net3010),
    .Y(_04479_));
 sky130_fd_sc_hd__nor2_1 _37715_ (.A(net1388),
    .B(_16362_),
    .Y(_16429_));
 sky130_fd_sc_hd__o21ai_0 _37716_ (.A1(net1186),
    .A2(_16354_),
    .B1(net1178),
    .Y(_16430_));
 sky130_fd_sc_hd__o22ai_1 _37717_ (.A1(_16429_),
    .A2(_16430_),
    .B1(net1178),
    .B2(_16292_),
    .Y(_16431_));
 sky130_fd_sc_hd__a21oi_1 _37719_ (.A1(_16382_),
    .A2(net1073),
    .B1(net1927),
    .Y(_16433_));
 sky130_fd_sc_hd__o21ai_0 _37720_ (.A1(net1073),
    .A2(_16431_),
    .B1(_16433_),
    .Y(_16434_));
 sky130_fd_sc_hd__nand2_1 _37722_ (.A(net1927),
    .B(\inst$top.soc.cpu.shifter.m_result$7[5] ),
    .Y(_16436_));
 sky130_fd_sc_hd__a21oi_1 _37723_ (.A1(_16434_),
    .A2(_16436_),
    .B1(net3011),
    .Y(_04480_));
 sky130_fd_sc_hd__a21oi_1 _37724_ (.A1(_16404_),
    .A2(net1186),
    .B1(net1391),
    .Y(_16437_));
 sky130_fd_sc_hd__o21ai_0 _37725_ (.A1(net1186),
    .A2(_16202_),
    .B1(_16437_),
    .Y(_16438_));
 sky130_fd_sc_hd__o21ai_0 _37726_ (.A1(net1175),
    .A2(_16312_),
    .B1(_16438_),
    .Y(_16439_));
 sky130_fd_sc_hd__a21oi_1 _37727_ (.A1(_16386_),
    .A2(net1072),
    .B1(net1926),
    .Y(_16440_));
 sky130_fd_sc_hd__o21ai_0 _37728_ (.A1(net1072),
    .A2(_16439_),
    .B1(_16440_),
    .Y(_16441_));
 sky130_fd_sc_hd__nand2_1 _37729_ (.A(net1926),
    .B(\inst$top.soc.cpu.shifter.m_result$7[6] ),
    .Y(_16442_));
 sky130_fd_sc_hd__a21oi_1 _37730_ (.A1(_16441_),
    .A2(_16442_),
    .B1(net3010),
    .Y(_04481_));
 sky130_fd_sc_hd__a21oi_1 _37731_ (.A1(_16416_),
    .A2(net1186),
    .B1(net1391),
    .Y(_16443_));
 sky130_fd_sc_hd__o21ai_0 _37732_ (.A1(net1187),
    .A2(_16249_),
    .B1(_16443_),
    .Y(_16444_));
 sky130_fd_sc_hd__o21ai_0 _37733_ (.A1(net1175),
    .A2(_16320_),
    .B1(_16444_),
    .Y(_16445_));
 sky130_fd_sc_hd__nand2_1 _37734_ (.A(_16389_),
    .B(_16390_),
    .Y(_16446_));
 sky130_fd_sc_hd__a21oi_1 _37735_ (.A1(_16446_),
    .A2(net1072),
    .B1(net1926),
    .Y(_16447_));
 sky130_fd_sc_hd__o21ai_0 _37736_ (.A1(net1072),
    .A2(_16445_),
    .B1(_16447_),
    .Y(_16448_));
 sky130_fd_sc_hd__nand2_1 _37737_ (.A(net1926),
    .B(\inst$top.soc.cpu.shifter.m_result$7[7] ),
    .Y(_16449_));
 sky130_fd_sc_hd__a21oi_1 _37738_ (.A1(_16448_),
    .A2(_16449_),
    .B1(net3011),
    .Y(_04482_));
 sky130_fd_sc_hd__nand2_1 _37739_ (.A(_16393_),
    .B(net1073),
    .Y(_16450_));
 sky130_fd_sc_hd__nand2_1 _37740_ (.A(_16188_),
    .B(net1178),
    .Y(_16451_));
 sky130_fd_sc_hd__o211ai_1 _37741_ (.A1(net1178),
    .A2(_16124_),
    .B1(net1200),
    .C1(_16451_),
    .Y(_16452_));
 sky130_fd_sc_hd__nand3_1 _37742_ (.A(_16450_),
    .B(net2297),
    .C(_16452_),
    .Y(_16453_));
 sky130_fd_sc_hd__o211ai_1 _37743_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[8] ),
    .A2(net2297),
    .B1(net2183),
    .C1(_16453_),
    .Y(_16454_));
 sky130_fd_sc_hd__inv_2 _37744_ (.A(_16454_),
    .Y(_04483_));
 sky130_fd_sc_hd__nand2_1 _37745_ (.A(_16356_),
    .B(net1178),
    .Y(_16455_));
 sky130_fd_sc_hd__o211ai_1 _37746_ (.A1(net1175),
    .A2(_16339_),
    .B1(net1198),
    .C1(_16455_),
    .Y(_16456_));
 sky130_fd_sc_hd__nand2_1 _37747_ (.A(_16395_),
    .B(net1073),
    .Y(_16457_));
 sky130_fd_sc_hd__nand3_1 _37748_ (.A(_16456_),
    .B(net2297),
    .C(_16457_),
    .Y(_16458_));
 sky130_fd_sc_hd__o211ai_1 _37749_ (.A1(\inst$top.soc.cpu.shifter.m_result$7[9] ),
    .A2(net2297),
    .B1(net2183),
    .C1(_16458_),
    .Y(_16459_));
 sky130_fd_sc_hd__inv_2 _37750_ (.A(_16459_),
    .Y(_04484_));
 sky130_fd_sc_hd__nor2_1 _37752_ (.A(\inst$top.soc.cpu.sink__payload$12[100] ),
    .B(net696),
    .Y(_16461_));
 sky130_fd_sc_hd__o21ai_1 _37753_ (.A1(\inst$top.soc.cpu.sink__payload$6[43] ),
    .A2(net650),
    .B1(net2143),
    .Y(_16462_));
 sky130_fd_sc_hd__nor2_4 _37754_ (.A(_16461_),
    .B(_16462_),
    .Y(_04485_));
 sky130_fd_sc_hd__nor2_1 _37755_ (.A(\inst$top.soc.cpu.sink__payload$12[101] ),
    .B(net700),
    .Y(_16463_));
 sky130_fd_sc_hd__o21ai_1 _37756_ (.A1(net2767),
    .A2(net654),
    .B1(net2147),
    .Y(_16464_));
 sky130_fd_sc_hd__nor2_4 _37757_ (.A(_16463_),
    .B(_16464_),
    .Y(_04486_));
 sky130_fd_sc_hd__nor2_1 _37758_ (.A(\inst$top.soc.cpu.sink__payload$12[102] ),
    .B(net700),
    .Y(_16465_));
 sky130_fd_sc_hd__o21ai_1 _37759_ (.A1(net2724),
    .A2(net654),
    .B1(net2147),
    .Y(_16466_));
 sky130_fd_sc_hd__nor2_4 _37760_ (.A(_16465_),
    .B(_16466_),
    .Y(_04487_));
 sky130_fd_sc_hd__nor2_1 _37761_ (.A(\inst$top.soc.cpu.sink__payload$12[103] ),
    .B(net700),
    .Y(_16467_));
 sky130_fd_sc_hd__o21ai_1 _37763_ (.A1(net2703),
    .A2(net654),
    .B1(net2147),
    .Y(_16469_));
 sky130_fd_sc_hd__nor2_4 _37764_ (.A(_16467_),
    .B(_16469_),
    .Y(_04488_));
 sky130_fd_sc_hd__nor2_1 _37765_ (.A(\inst$top.soc.cpu.sink__payload$12[104] ),
    .B(net703),
    .Y(_16470_));
 sky130_fd_sc_hd__o21ai_1 _37767_ (.A1(net2696),
    .A2(net654),
    .B1(net2148),
    .Y(_16472_));
 sky130_fd_sc_hd__nor2_4 _37768_ (.A(_16470_),
    .B(_16472_),
    .Y(_04489_));
 sky130_fd_sc_hd__nor2_1 _37769_ (.A(\inst$top.soc.cpu.sink__payload$12[105] ),
    .B(net702),
    .Y(_16473_));
 sky130_fd_sc_hd__o21ai_1 _37770_ (.A1(net2690),
    .A2(net655),
    .B1(net2148),
    .Y(_16474_));
 sky130_fd_sc_hd__nor2_4 _37771_ (.A(_16473_),
    .B(_16474_),
    .Y(_04490_));
 sky130_fd_sc_hd__nor2_1 _37772_ (.A(\inst$top.soc.cpu.d.sink__payload.rd_we ),
    .B(net693),
    .Y(_16475_));
 sky130_fd_sc_hd__inv_1 _37773_ (.A(\inst$top.soc.cpu.sink__payload$6[45] ),
    .Y(_16476_));
 sky130_fd_sc_hd__nand3_1 _37774_ (.A(_20300_),
    .B(_11908_),
    .C(_16476_),
    .Y(_16477_));
 sky130_fd_sc_hd__nand2_1 _37775_ (.A(_16477_),
    .B(_06040_),
    .Y(_16478_));
 sky130_fd_sc_hd__nand2_1 _37776_ (.A(net693),
    .B(_16478_),
    .Y(_16479_));
 sky130_fd_sc_hd__nand2_1 _37777_ (.A(_16479_),
    .B(net2144),
    .Y(_16480_));
 sky130_fd_sc_hd__nor2_4 _37778_ (.A(_16475_),
    .B(_16480_),
    .Y(_04491_));
 sky130_fd_sc_hd__nor2_1 _37779_ (.A(\inst$top.soc.cpu.d.sink__payload.rs1_re ),
    .B(net690),
    .Y(_16481_));
 sky130_fd_sc_hd__nand2_1 _37781_ (.A(net687),
    .B(net1191),
    .Y(_16483_));
 sky130_fd_sc_hd__nand2_1 _37782_ (.A(_16483_),
    .B(net2074),
    .Y(_16484_));
 sky130_fd_sc_hd__nor2_4 _37783_ (.A(_16481_),
    .B(_16484_),
    .Y(_04492_));
 sky130_fd_sc_hd__nor2_1 _37784_ (.A(\inst$top.soc.cpu.d.sink__payload.rs2_re ),
    .B(net687),
    .Y(_16485_));
 sky130_fd_sc_hd__nand2_1 _37785_ (.A(_20312_),
    .B(_20296_),
    .Y(_16486_));
 sky130_fd_sc_hd__o21ai_1 _37786_ (.A1(_16486_),
    .A2(net643),
    .B1(net2077),
    .Y(_16487_));
 sky130_fd_sc_hd__nor2_4 _37787_ (.A(_16485_),
    .B(_16487_),
    .Y(_04493_));
 sky130_fd_sc_hd__nor2_1 _37788_ (.A(\inst$top.soc.cpu.sink__payload$12[10] ),
    .B(net680),
    .Y(_16488_));
 sky130_fd_sc_hd__o21ai_1 _37789_ (.A1(\inst$top.soc.cpu.sink__payload$6[10] ),
    .A2(net637),
    .B1(net2067),
    .Y(_16489_));
 sky130_fd_sc_hd__nor2_4 _37790_ (.A(_16488_),
    .B(_16489_),
    .Y(_04494_));
 sky130_fd_sc_hd__nor2_1 _37792_ (.A(\inst$top.soc.cpu.sink__payload$12[111] ),
    .B(net695),
    .Y(_16491_));
 sky130_fd_sc_hd__o21ai_1 _37793_ (.A1(_06044_),
    .A2(net648),
    .B1(net2142),
    .Y(_16492_));
 sky130_fd_sc_hd__nor2_4 _37794_ (.A(_16491_),
    .B(_16492_),
    .Y(_04495_));
 sky130_fd_sc_hd__nor2_1 _37795_ (.A(\inst$top.soc.cpu.sink__payload$12[112] ),
    .B(net693),
    .Y(_16493_));
 sky130_fd_sc_hd__o21ai_1 _37796_ (.A1(_06042_),
    .A2(net648),
    .B1(net2144),
    .Y(_16494_));
 sky130_fd_sc_hd__nor2_4 _37797_ (.A(_16493_),
    .B(_16494_),
    .Y(_04496_));
 sky130_fd_sc_hd__nor2_1 _37798_ (.A(\inst$top.soc.cpu.sink__payload$12[113] ),
    .B(net693),
    .Y(_16495_));
 sky130_fd_sc_hd__o21ai_1 _37799_ (.A1(\inst$top.soc.cpu.csrf.d_addr[4] ),
    .A2(net648),
    .B1(net2142),
    .Y(_16496_));
 sky130_fd_sc_hd__nor2_4 _37800_ (.A(_16495_),
    .B(_16496_),
    .Y(_04497_));
 sky130_fd_sc_hd__nor2_1 _37801_ (.A(\inst$top.soc.cpu.sink__payload$12[114] ),
    .B(net694),
    .Y(_16497_));
 sky130_fd_sc_hd__o21ai_1 _37802_ (.A1(\inst$top.soc.cpu.csrf.d_addr[5] ),
    .A2(net647),
    .B1(net2141),
    .Y(_16498_));
 sky130_fd_sc_hd__nor2_4 _37803_ (.A(_16497_),
    .B(_16498_),
    .Y(_04498_));
 sky130_fd_sc_hd__nor2_1 _37804_ (.A(\inst$top.soc.cpu.sink__payload$12[115] ),
    .B(net694),
    .Y(_16499_));
 sky130_fd_sc_hd__o21ai_1 _37805_ (.A1(\inst$top.soc.cpu.csrf.d_addr[6] ),
    .A2(net647),
    .B1(net2141),
    .Y(_16500_));
 sky130_fd_sc_hd__nor2_4 _37806_ (.A(_16499_),
    .B(_16500_),
    .Y(_04499_));
 sky130_fd_sc_hd__nor2_1 _37807_ (.A(\inst$top.soc.cpu.sink__payload$12[116] ),
    .B(net683),
    .Y(_16501_));
 sky130_fd_sc_hd__o21ai_1 _37809_ (.A1(\inst$top.soc.cpu.csrf.d_addr[7] ),
    .A2(net641),
    .B1(net2074),
    .Y(_16503_));
 sky130_fd_sc_hd__nor2_4 _37810_ (.A(_16501_),
    .B(_16503_),
    .Y(_04500_));
 sky130_fd_sc_hd__nor2_1 _37811_ (.A(\inst$top.soc.cpu.sink__payload$12[117] ),
    .B(net687),
    .Y(_16504_));
 sky130_fd_sc_hd__o21ai_1 _37813_ (.A1(\inst$top.soc.cpu.csrf.d_addr[8] ),
    .A2(net643),
    .B1(net2077),
    .Y(_16506_));
 sky130_fd_sc_hd__nor2_4 _37814_ (.A(_16504_),
    .B(_16506_),
    .Y(_04501_));
 sky130_fd_sc_hd__nor2_1 _37815_ (.A(\inst$top.soc.cpu.sink__payload$12[118] ),
    .B(net683),
    .Y(_16507_));
 sky130_fd_sc_hd__o21ai_1 _37816_ (.A1(\inst$top.soc.cpu.csrf.d_addr[9] ),
    .A2(net641),
    .B1(net2074),
    .Y(_16508_));
 sky130_fd_sc_hd__nor2_4 _37817_ (.A(_16507_),
    .B(_16508_),
    .Y(_04502_));
 sky130_fd_sc_hd__nor2_1 _37818_ (.A(\inst$top.soc.cpu.sink__payload$12[119] ),
    .B(net699),
    .Y(_16509_));
 sky130_fd_sc_hd__o21ai_1 _37819_ (.A1(\inst$top.soc.cpu.csrf.d_addr[10] ),
    .A2(net648),
    .B1(net2142),
    .Y(_16510_));
 sky130_fd_sc_hd__nor2_4 _37820_ (.A(_16509_),
    .B(_16510_),
    .Y(_04503_));
 sky130_fd_sc_hd__nor2_1 _37821_ (.A(\inst$top.soc.cpu.sink__payload$12[11] ),
    .B(net680),
    .Y(_16511_));
 sky130_fd_sc_hd__o21ai_1 _37822_ (.A1(\inst$top.soc.cpu.sink__payload$6[11] ),
    .A2(net637),
    .B1(net2065),
    .Y(_16512_));
 sky130_fd_sc_hd__nor2_4 _37823_ (.A(_16511_),
    .B(_16512_),
    .Y(_04504_));
 sky130_fd_sc_hd__nor2_1 _37825_ (.A(\inst$top.soc.cpu.sink__payload$12[120] ),
    .B(net699),
    .Y(_16514_));
 sky130_fd_sc_hd__o21ai_1 _37826_ (.A1(\inst$top.soc.cpu.csrf.d_addr[11] ),
    .A2(net653),
    .B1(net2146),
    .Y(_16515_));
 sky130_fd_sc_hd__nor2_4 _37827_ (.A(_16514_),
    .B(_16515_),
    .Y(_04505_));
 sky130_fd_sc_hd__nor2_1 _37828_ (.A(\inst$top.soc.cpu.sink__payload$12[121] ),
    .B(net694),
    .Y(_16516_));
 sky130_fd_sc_hd__o21ai_1 _37829_ (.A1(\inst$top.soc.cpu.d_offset[12] ),
    .A2(net648),
    .B1(net2142),
    .Y(_16517_));
 sky130_fd_sc_hd__nor2_4 _37830_ (.A(_16516_),
    .B(_16517_),
    .Y(_04506_));
 sky130_fd_sc_hd__nor2_1 _37831_ (.A(\inst$top.soc.cpu.sink__payload$12[122] ),
    .B(net694),
    .Y(_16518_));
 sky130_fd_sc_hd__o21ai_1 _37832_ (.A1(\inst$top.soc.cpu.d_offset[13] ),
    .A2(net647),
    .B1(net2142),
    .Y(_16519_));
 sky130_fd_sc_hd__nor2_4 _37833_ (.A(_16518_),
    .B(_16519_),
    .Y(_04507_));
 sky130_fd_sc_hd__nor2_1 _37834_ (.A(\inst$top.soc.cpu.sink__payload$12[123] ),
    .B(net688),
    .Y(_16520_));
 sky130_fd_sc_hd__o21ai_1 _37835_ (.A1(\inst$top.soc.cpu.d_offset[14] ),
    .A2(net647),
    .B1(net2077),
    .Y(_16521_));
 sky130_fd_sc_hd__nor2_4 _37836_ (.A(_16520_),
    .B(_16521_),
    .Y(_04508_));
 sky130_fd_sc_hd__nor2_1 _37837_ (.A(\inst$top.soc.cpu.sink__payload$12[124] ),
    .B(net693),
    .Y(_16522_));
 sky130_fd_sc_hd__o21ai_1 _37838_ (.A1(\inst$top.soc.cpu.d_offset[15] ),
    .A2(net648),
    .B1(net2144),
    .Y(_16523_));
 sky130_fd_sc_hd__nor2_4 _37839_ (.A(_16522_),
    .B(_16523_),
    .Y(_04509_));
 sky130_fd_sc_hd__nor2_1 _37840_ (.A(\inst$top.soc.cpu.sink__payload$12[125] ),
    .B(net696),
    .Y(_16524_));
 sky130_fd_sc_hd__o21ai_1 _37842_ (.A1(\inst$top.soc.cpu.d_offset[16] ),
    .A2(net650),
    .B1(net2144),
    .Y(_16526_));
 sky130_fd_sc_hd__nor2_4 _37843_ (.A(_16524_),
    .B(_16526_),
    .Y(_04510_));
 sky130_fd_sc_hd__nor2_1 _37844_ (.A(\inst$top.soc.cpu.sink__payload$12[126] ),
    .B(net696),
    .Y(_16527_));
 sky130_fd_sc_hd__o21ai_1 _37846_ (.A1(\inst$top.soc.cpu.d_offset[17] ),
    .A2(net650),
    .B1(net2143),
    .Y(_16529_));
 sky130_fd_sc_hd__nor2_4 _37847_ (.A(_16527_),
    .B(_16529_),
    .Y(_04511_));
 sky130_fd_sc_hd__nor2_1 _37848_ (.A(\inst$top.soc.cpu.sink__payload$12[127] ),
    .B(net693),
    .Y(_16530_));
 sky130_fd_sc_hd__o21ai_1 _37849_ (.A1(\inst$top.soc.cpu.d_offset[18] ),
    .A2(net650),
    .B1(net2143),
    .Y(_16531_));
 sky130_fd_sc_hd__nor2_4 _37850_ (.A(_16530_),
    .B(_16531_),
    .Y(_04512_));
 sky130_fd_sc_hd__nor2_1 _37851_ (.A(\inst$top.soc.cpu.sink__payload$12[128] ),
    .B(net693),
    .Y(_16532_));
 sky130_fd_sc_hd__o21ai_1 _37852_ (.A1(\inst$top.soc.cpu.d_offset[19] ),
    .A2(net650),
    .B1(net2143),
    .Y(_16533_));
 sky130_fd_sc_hd__nor2_4 _37853_ (.A(_16532_),
    .B(_16533_),
    .Y(_04513_));
 sky130_fd_sc_hd__nor2_1 _37854_ (.A(\inst$top.soc.cpu.sink__payload$12[129] ),
    .B(net694),
    .Y(_16534_));
 sky130_fd_sc_hd__o21ai_1 _37855_ (.A1(\inst$top.soc.cpu.d_offset[20] ),
    .A2(net647),
    .B1(net2141),
    .Y(_16535_));
 sky130_fd_sc_hd__nor2_4 _37856_ (.A(_16534_),
    .B(_16535_),
    .Y(_04514_));
 sky130_fd_sc_hd__nor2_1 _37858_ (.A(\inst$top.soc.cpu.sink__payload$12[12] ),
    .B(net680),
    .Y(_16537_));
 sky130_fd_sc_hd__o21ai_1 _37859_ (.A1(\inst$top.soc.cpu.sink__payload$6[12] ),
    .A2(net645),
    .B1(net2071),
    .Y(_16538_));
 sky130_fd_sc_hd__nor2_4 _37860_ (.A(_16537_),
    .B(_16538_),
    .Y(_04515_));
 sky130_fd_sc_hd__nor2_1 _37861_ (.A(\inst$top.soc.cpu.sink__payload$12[130] ),
    .B(net693),
    .Y(_16539_));
 sky130_fd_sc_hd__o21ai_1 _37862_ (.A1(\inst$top.soc.cpu.d_offset[21] ),
    .A2(net648),
    .B1(net2141),
    .Y(_16540_));
 sky130_fd_sc_hd__nor2_4 _37863_ (.A(_16539_),
    .B(_16540_),
    .Y(_04516_));
 sky130_fd_sc_hd__nor2_1 _37864_ (.A(\inst$top.soc.cpu.sink__payload$12[131] ),
    .B(net693),
    .Y(_16541_));
 sky130_fd_sc_hd__o21ai_1 _37865_ (.A1(\inst$top.soc.cpu.d_offset[22] ),
    .A2(net648),
    .B1(net2141),
    .Y(_16542_));
 sky130_fd_sc_hd__nor2_4 _37866_ (.A(_16541_),
    .B(_16542_),
    .Y(_04517_));
 sky130_fd_sc_hd__nor2_1 _37867_ (.A(\inst$top.soc.cpu.sink__payload$12[132] ),
    .B(net694),
    .Y(_16543_));
 sky130_fd_sc_hd__o21ai_1 _37868_ (.A1(\inst$top.soc.cpu.d_offset[23] ),
    .A2(net647),
    .B1(net2141),
    .Y(_16544_));
 sky130_fd_sc_hd__nor2_4 _37869_ (.A(_16543_),
    .B(_16544_),
    .Y(_04518_));
 sky130_fd_sc_hd__nor2_1 _37870_ (.A(\inst$top.soc.cpu.sink__payload$12[133] ),
    .B(net688),
    .Y(_16545_));
 sky130_fd_sc_hd__o21ai_1 _37871_ (.A1(\inst$top.soc.cpu.d_offset[24] ),
    .A2(net647),
    .B1(net2076),
    .Y(_16546_));
 sky130_fd_sc_hd__nor2_4 _37872_ (.A(_16545_),
    .B(_16546_),
    .Y(_04519_));
 sky130_fd_sc_hd__nor2_1 _37873_ (.A(\inst$top.soc.cpu.sink__payload$12[134] ),
    .B(net694),
    .Y(_16547_));
 sky130_fd_sc_hd__o21ai_1 _37876_ (.A1(\inst$top.soc.cpu.d_offset[25] ),
    .A2(net648),
    .B1(net2141),
    .Y(_16550_));
 sky130_fd_sc_hd__nor2_4 _37877_ (.A(_16547_),
    .B(_16550_),
    .Y(_04520_));
 sky130_fd_sc_hd__nor2_1 _37878_ (.A(\inst$top.soc.cpu.sink__payload$12[135] ),
    .B(net687),
    .Y(_16551_));
 sky130_fd_sc_hd__o21ai_1 _37880_ (.A1(\inst$top.soc.cpu.d_offset[26] ),
    .A2(net643),
    .B1(net2076),
    .Y(_16553_));
 sky130_fd_sc_hd__nor2_4 _37881_ (.A(_16551_),
    .B(_16553_),
    .Y(_04521_));
 sky130_fd_sc_hd__nor2_1 _37882_ (.A(\inst$top.soc.cpu.sink__payload$12[136] ),
    .B(net688),
    .Y(_16554_));
 sky130_fd_sc_hd__o21ai_1 _37883_ (.A1(\inst$top.soc.cpu.d_offset[27] ),
    .A2(net643),
    .B1(net2076),
    .Y(_16555_));
 sky130_fd_sc_hd__nor2_4 _37884_ (.A(_16554_),
    .B(_16555_),
    .Y(_04522_));
 sky130_fd_sc_hd__nor2_1 _37885_ (.A(\inst$top.soc.cpu.sink__payload$12[137] ),
    .B(net688),
    .Y(_16556_));
 sky130_fd_sc_hd__o21ai_1 _37886_ (.A1(\inst$top.soc.cpu.d_offset[28] ),
    .A2(net643),
    .B1(net2076),
    .Y(_16557_));
 sky130_fd_sc_hd__nor2_4 _37887_ (.A(_16556_),
    .B(_16557_),
    .Y(_04523_));
 sky130_fd_sc_hd__nor2_1 _37888_ (.A(\inst$top.soc.cpu.sink__payload$12[138] ),
    .B(net687),
    .Y(_16558_));
 sky130_fd_sc_hd__o21ai_1 _37889_ (.A1(\inst$top.soc.cpu.d_offset[29] ),
    .A2(net643),
    .B1(net2076),
    .Y(_16559_));
 sky130_fd_sc_hd__nor2_4 _37890_ (.A(_16558_),
    .B(_16559_),
    .Y(_04524_));
 sky130_fd_sc_hd__nor2_1 _37892_ (.A(\inst$top.soc.cpu.sink__payload$12[139] ),
    .B(net687),
    .Y(_16561_));
 sky130_fd_sc_hd__o21ai_1 _37893_ (.A1(\inst$top.soc.cpu.d_offset[30] ),
    .A2(net643),
    .B1(net2076),
    .Y(_16562_));
 sky130_fd_sc_hd__nor2_4 _37894_ (.A(_16561_),
    .B(_16562_),
    .Y(_04525_));
 sky130_fd_sc_hd__nor2_1 _37895_ (.A(\inst$top.soc.cpu.sink__payload$12[13] ),
    .B(net684),
    .Y(_16563_));
 sky130_fd_sc_hd__o21ai_1 _37896_ (.A1(\inst$top.soc.cpu.sink__payload$6[13] ),
    .A2(net641),
    .B1(net2074),
    .Y(_16564_));
 sky130_fd_sc_hd__nor2_4 _37897_ (.A(_16563_),
    .B(_16564_),
    .Y(_04526_));
 sky130_fd_sc_hd__nor2_1 _37898_ (.A(\inst$top.soc.cpu.sink__payload$12[140] ),
    .B(net700),
    .Y(_16565_));
 sky130_fd_sc_hd__nand2_1 _37899_ (.A(net700),
    .B(_11911_),
    .Y(_16566_));
 sky130_fd_sc_hd__nand2_1 _37900_ (.A(_16566_),
    .B(net2147),
    .Y(_16567_));
 sky130_fd_sc_hd__nor2_4 _37901_ (.A(_16565_),
    .B(_16567_),
    .Y(_04527_));
 sky130_fd_sc_hd__nor2_1 _37902_ (.A(\inst$top.soc.cpu.sink__payload$6[61] ),
    .B(\inst$top.soc.cpu.sink__payload$6[63] ),
    .Y(_16568_));
 sky130_fd_sc_hd__inv_1 _37903_ (.A(_16568_),
    .Y(_16569_));
 sky130_fd_sc_hd__nor2_1 _37904_ (.A(\inst$top.soc.cpu.sink__payload$6[62] ),
    .B(_16569_),
    .Y(_16570_));
 sky130_fd_sc_hd__inv_1 _37905_ (.A(_16570_),
    .Y(_16571_));
 sky130_fd_sc_hd__nor4_1 _37906_ (.A(\inst$top.soc.cpu.sink__payload$6[58] ),
    .B(\inst$top.soc.cpu.sink__payload$6[60] ),
    .C(\inst$top.soc.cpu.sink__payload$6[57] ),
    .D(\inst$top.soc.cpu.sink__payload$6[59] ),
    .Y(_16572_));
 sky130_fd_sc_hd__inv_1 _37907_ (.A(_16572_),
    .Y(_16573_));
 sky130_fd_sc_hd__nor2_1 _37908_ (.A(_16571_),
    .B(_16573_),
    .Y(_16574_));
 sky130_fd_sc_hd__o21ai_0 _37909_ (.A1(_20282_),
    .A2(_16574_),
    .B1(_20306_),
    .Y(_16575_));
 sky130_fd_sc_hd__nand3b_1 _37910_ (.A_N(_16575_),
    .B(net2820),
    .C(_16052_),
    .Y(_16576_));
 sky130_fd_sc_hd__nand2_1 _37911_ (.A(_16572_),
    .B(_16568_),
    .Y(_16577_));
 sky130_fd_sc_hd__inv_1 _37912_ (.A(_16577_),
    .Y(_16578_));
 sky130_fd_sc_hd__o211ai_1 _37913_ (.A1(_20282_),
    .A2(_16578_),
    .B1(_20306_),
    .C1(_16042_),
    .Y(_16579_));
 sky130_fd_sc_hd__inv_1 _37914_ (.A(_20354_),
    .Y(_16580_));
 sky130_fd_sc_hd__nand2_1 _37915_ (.A(_16580_),
    .B(_20311_),
    .Y(_16581_));
 sky130_fd_sc_hd__inv_1 _37916_ (.A(_16581_),
    .Y(_16582_));
 sky130_fd_sc_hd__nand3_1 _37917_ (.A(_16576_),
    .B(_16579_),
    .C(_16582_),
    .Y(_16583_));
 sky130_fd_sc_hd__nand2_1 _37918_ (.A(net700),
    .B(_16583_),
    .Y(_16584_));
 sky130_fd_sc_hd__nand2_1 _37919_ (.A(net650),
    .B(\inst$top.soc.cpu.d.sink__payload.bypass_x ),
    .Y(_16585_));
 sky130_fd_sc_hd__a21oi_4 _37920_ (.A1(_16584_),
    .A2(_16585_),
    .B1(net2993),
    .Y(_04528_));
 sky130_fd_sc_hd__a2111oi_0 _37921_ (.A1(_11908_),
    .A2(\inst$top.soc.cpu.sink__payload$6[62] ),
    .B1(_16052_),
    .C1(_16569_),
    .D1(_16573_),
    .Y(_16586_));
 sky130_fd_sc_hd__nand2_1 _37922_ (.A(_16586_),
    .B(_20306_),
    .Y(_16587_));
 sky130_fd_sc_hd__nor3_1 _37923_ (.A(net2820),
    .B(_16476_),
    .C(_16575_),
    .Y(_16588_));
 sky130_fd_sc_hd__inv_1 _37924_ (.A(_16588_),
    .Y(_16589_));
 sky130_fd_sc_hd__nor2_1 _37925_ (.A(\inst$top.soc.cpu.sink__payload$6[58] ),
    .B(\inst$top.soc.cpu.sink__payload$6[59] ),
    .Y(_16590_));
 sky130_fd_sc_hd__inv_1 _37926_ (.A(_16590_),
    .Y(_16591_));
 sky130_fd_sc_hd__nor2_1 _37927_ (.A(\inst$top.soc.cpu.sink__payload$6[60] ),
    .B(_16571_),
    .Y(_16592_));
 sky130_fd_sc_hd__inv_1 _37928_ (.A(_16592_),
    .Y(_16593_));
 sky130_fd_sc_hd__nor3_1 _37929_ (.A(_06045_),
    .B(_16591_),
    .C(_16593_),
    .Y(_16594_));
 sky130_fd_sc_hd__nor2_1 _37930_ (.A(_20292_),
    .B(_20305_),
    .Y(_16595_));
 sky130_fd_sc_hd__nand3_1 _37931_ (.A(_16594_),
    .B(net2820),
    .C(_16595_),
    .Y(_16596_));
 sky130_fd_sc_hd__nand3_1 _37932_ (.A(_16587_),
    .B(_16589_),
    .C(_16596_),
    .Y(_16597_));
 sky130_fd_sc_hd__nand2_1 _37933_ (.A(net700),
    .B(_16597_),
    .Y(_16598_));
 sky130_fd_sc_hd__nand2_1 _37934_ (.A(net654),
    .B(\inst$top.soc.cpu.d.sink__payload.bypass_m ),
    .Y(_16599_));
 sky130_fd_sc_hd__a21oi_4 _37935_ (.A1(_16598_),
    .A2(_16599_),
    .B1(net2993),
    .Y(_04529_));
 sky130_fd_sc_hd__nor2_1 _37936_ (.A(\inst$top.soc.cpu.sink__payload$12[143] ),
    .B(net694),
    .Y(_16600_));
 sky130_fd_sc_hd__o21ai_1 _37937_ (.A1(\inst$top.soc.cpu.sink__payload$6[44] ),
    .A2(net647),
    .B1(net2141),
    .Y(_16601_));
 sky130_fd_sc_hd__nor2_4 _37938_ (.A(_16600_),
    .B(_16601_),
    .Y(_04530_));
 sky130_fd_sc_hd__nor2_1 _37939_ (.A(\inst$top.soc.cpu.sink__payload$12[144] ),
    .B(net694),
    .Y(_16602_));
 sky130_fd_sc_hd__o21ai_1 _37940_ (.A1(\inst$top.soc.cpu.sink__payload$6[45] ),
    .A2(net647),
    .B1(net2141),
    .Y(_16603_));
 sky130_fd_sc_hd__nor2_4 _37941_ (.A(_16602_),
    .B(_16603_),
    .Y(_04531_));
 sky130_fd_sc_hd__nor2_1 _37942_ (.A(\inst$top.soc.cpu.d.sink__payload.lui ),
    .B(net699),
    .Y(_16604_));
 sky130_fd_sc_hd__o21ai_1 _37943_ (.A1(_20309_),
    .A2(net653),
    .B1(net2147),
    .Y(_16605_));
 sky130_fd_sc_hd__nor2_4 _37944_ (.A(_16604_),
    .B(_16605_),
    .Y(_04532_));
 sky130_fd_sc_hd__nor2_1 _37945_ (.A(\inst$top.soc.cpu.d.sink__payload.auipc ),
    .B(net699),
    .Y(_16606_));
 sky130_fd_sc_hd__o21ai_1 _37947_ (.A1(_20310_),
    .A2(net653),
    .B1(net2146),
    .Y(_16608_));
 sky130_fd_sc_hd__nor2_4 _37948_ (.A(_16606_),
    .B(_16608_),
    .Y(_04533_));
 sky130_fd_sc_hd__nor2_1 _37949_ (.A(\inst$top.soc.cpu.d.sink__payload.load ),
    .B(net687),
    .Y(_16609_));
 sky130_fd_sc_hd__o211ai_1 _37950_ (.A1(_11908_),
    .A2(_16476_),
    .B1(_16045_),
    .C1(_20290_),
    .Y(_16610_));
 sky130_fd_sc_hd__nand2_1 _37951_ (.A(net687),
    .B(_16610_),
    .Y(_16611_));
 sky130_fd_sc_hd__nand2_1 _37952_ (.A(_16611_),
    .B(net2077),
    .Y(_16612_));
 sky130_fd_sc_hd__nor2_4 _37953_ (.A(_16609_),
    .B(_16612_),
    .Y(_04534_));
 sky130_fd_sc_hd__nor2_1 _37954_ (.A(\inst$top.soc.cpu.d.sink__payload.store ),
    .B(net688),
    .Y(_16613_));
 sky130_fd_sc_hd__nor3_1 _37955_ (.A(net2820),
    .B(_16046_),
    .C(_09364_),
    .Y(_16614_));
 sky130_fd_sc_hd__o21ai_1 _37957_ (.A1(_16614_),
    .A2(net647),
    .B1(net2077),
    .Y(_16616_));
 sky130_fd_sc_hd__nor2_4 _37958_ (.A(_16613_),
    .B(_16616_),
    .Y(_04535_));
 sky130_fd_sc_hd__nor2_1 _37959_ (.A(\inst$top.soc.cpu.sink__payload$12[14] ),
    .B(net679),
    .Y(_16617_));
 sky130_fd_sc_hd__o21ai_1 _37960_ (.A1(\inst$top.soc.cpu.sink__payload$6[14] ),
    .A2(net634),
    .B1(net2068),
    .Y(_16618_));
 sky130_fd_sc_hd__nor2_4 _37961_ (.A(_16617_),
    .B(_16618_),
    .Y(_04536_));
 sky130_fd_sc_hd__nor4_1 _37962_ (.A(\inst$top.soc.cpu.sink__payload$6[61] ),
    .B(\inst$top.soc.cpu.sink__payload$6[63] ),
    .C(_06051_),
    .D(_16573_),
    .Y(_16619_));
 sky130_fd_sc_hd__nand3_1 _37963_ (.A(_16619_),
    .B(_16042_),
    .C(_16595_),
    .Y(_16620_));
 sky130_fd_sc_hd__nand3_1 _37964_ (.A(_16589_),
    .B(_11910_),
    .C(_16620_),
    .Y(_16621_));
 sky130_fd_sc_hd__nand2_1 _37965_ (.A(net699),
    .B(_16621_),
    .Y(_16622_));
 sky130_fd_sc_hd__nand2_1 _37967_ (.A(net655),
    .B(net2865),
    .Y(_16624_));
 sky130_fd_sc_hd__a21oi_4 _37968_ (.A1(_16622_),
    .A2(_16624_),
    .B1(net3005),
    .Y(_04537_));
 sky130_fd_sc_hd__nor2_1 _37970_ (.A(net2864),
    .B(net692),
    .Y(_16626_));
 sky130_fd_sc_hd__nand2_1 _37971_ (.A(net692),
    .B(_16576_),
    .Y(_16627_));
 sky130_fd_sc_hd__nand2_1 _37972_ (.A(_16627_),
    .B(net2080),
    .Y(_16628_));
 sky130_fd_sc_hd__nor2_4 _37973_ (.A(_16626_),
    .B(_16628_),
    .Y(_04538_));
 sky130_fd_sc_hd__nor2_1 _37974_ (.A(\inst$top.soc.cpu.d.sink__payload.multiply ),
    .B(net699),
    .Y(_16629_));
 sky130_fd_sc_hd__nand3_1 _37975_ (.A(_16594_),
    .B(_11908_),
    .C(_16595_),
    .Y(_16630_));
 sky130_fd_sc_hd__inv_1 _37976_ (.A(_16630_),
    .Y(_16631_));
 sky130_fd_sc_hd__o21ai_1 _37977_ (.A1(_16631_),
    .A2(net653),
    .B1(net2147),
    .Y(_16632_));
 sky130_fd_sc_hd__nor2_4 _37978_ (.A(_16629_),
    .B(_16632_),
    .Y(_04539_));
 sky130_fd_sc_hd__nor2_1 _37979_ (.A(\inst$top.soc.cpu.d.sink__payload.divide ),
    .B(net692),
    .Y(_16633_));
 sky130_fd_sc_hd__nand2_1 _37980_ (.A(net692),
    .B(_16596_),
    .Y(_16634_));
 sky130_fd_sc_hd__nand2_1 _37981_ (.A(_16634_),
    .B(net2146),
    .Y(_16635_));
 sky130_fd_sc_hd__nor2_4 _37982_ (.A(_16633_),
    .B(_16635_),
    .Y(_04540_));
 sky130_fd_sc_hd__nor2_1 _37983_ (.A(\inst$top.soc.cpu.d.sink__payload.shift ),
    .B(net699),
    .Y(_16636_));
 sky130_fd_sc_hd__o2111ai_1 _37984_ (.A1(net2820),
    .A2(_06051_),
    .B1(_20306_),
    .C1(_16051_),
    .D1(_16578_),
    .Y(_16637_));
 sky130_fd_sc_hd__inv_1 _37985_ (.A(_16637_),
    .Y(_16638_));
 sky130_fd_sc_hd__o21ai_1 _37986_ (.A1(_16638_),
    .A2(net653),
    .B1(net2080),
    .Y(_16639_));
 sky130_fd_sc_hd__nor2_4 _37987_ (.A(_16636_),
    .B(_16639_),
    .Y(_04541_));
 sky130_fd_sc_hd__nor2_2 _37988_ (.A(_11908_),
    .B(_16052_),
    .Y(_16640_));
 sky130_fd_sc_hd__nand2_1 _37989_ (.A(net658),
    .B(net2000),
    .Y(_16641_));
 sky130_fd_sc_hd__o21ai_1 _37990_ (.A1(_16640_),
    .A2(net659),
    .B1(_16641_),
    .Y(_16642_));
 sky130_fd_sc_hd__nor2_2 _37991_ (.A(net3010),
    .B(_16642_),
    .Y(_04542_));
 sky130_fd_sc_hd__nand2_1 _37992_ (.A(net700),
    .B(_16619_),
    .Y(_16643_));
 sky130_fd_sc_hd__nand2_1 _37993_ (.A(net655),
    .B(\inst$top.soc.cpu.d.sink__payload.sext ),
    .Y(_16644_));
 sky130_fd_sc_hd__a21oi_4 _37994_ (.A1(_16643_),
    .A2(_16644_),
    .B1(net3005),
    .Y(_04543_));
 sky130_fd_sc_hd__nor2_1 _37995_ (.A(net2852),
    .B(net692),
    .Y(_16645_));
 sky130_fd_sc_hd__a21oi_1 _37996_ (.A1(_20303_),
    .A2(_16042_),
    .B1(_20285_),
    .Y(_16646_));
 sky130_fd_sc_hd__inv_1 _37997_ (.A(_16646_),
    .Y(_16647_));
 sky130_fd_sc_hd__o21ai_1 _37998_ (.A1(_16647_),
    .A2(net644),
    .B1(net2080),
    .Y(_16648_));
 sky130_fd_sc_hd__nor2_4 _37999_ (.A(_16645_),
    .B(_16648_),
    .Y(_04544_));
 sky130_fd_sc_hd__nor2_1 _38000_ (.A(\inst$top.soc.cpu.d.sink__payload.compare ),
    .B(net699),
    .Y(_16649_));
 sky130_fd_sc_hd__o21ai_1 _38001_ (.A1(_16588_),
    .A2(net653),
    .B1(net2146),
    .Y(_16650_));
 sky130_fd_sc_hd__nor2_4 _38002_ (.A(_16649_),
    .B(_16650_),
    .Y(_04545_));
 sky130_fd_sc_hd__nor2_1 _38003_ (.A(\inst$top.soc.cpu.d.sink__payload.branch ),
    .B(net699),
    .Y(_16651_));
 sky130_fd_sc_hd__o21ai_1 _38004_ (.A1(_11909_),
    .A2(net653),
    .B1(net2146),
    .Y(_16652_));
 sky130_fd_sc_hd__nor2_4 _38005_ (.A(_16651_),
    .B(_16652_),
    .Y(_04546_));
 sky130_fd_sc_hd__nor2_1 _38006_ (.A(\inst$top.soc.cpu.sink__payload$12[15] ),
    .B(net683),
    .Y(_16653_));
 sky130_fd_sc_hd__o21ai_1 _38007_ (.A1(\inst$top.soc.cpu.sink__payload$6[15] ),
    .A2(net641),
    .B1(net2074),
    .Y(_16654_));
 sky130_fd_sc_hd__nor2_4 _38008_ (.A(_16653_),
    .B(_16654_),
    .Y(_04547_));
 sky130_fd_sc_hd__nor2_1 _38009_ (.A(\inst$top.soc.cpu.sink__payload$12[109] ),
    .B(net672),
    .Y(_16655_));
 sky130_fd_sc_hd__o21ai_1 _38011_ (.A1(_11017_),
    .A2(net633),
    .B1(net2033),
    .Y(_16657_));
 sky130_fd_sc_hd__nor2_4 _38012_ (.A(_16655_),
    .B(_16657_),
    .Y(_04548_));
 sky130_fd_sc_hd__nand2_1 _38013_ (.A(net644),
    .B(\inst$top.soc.cpu.sink__payload$12[110] ),
    .Y(_16658_));
 sky130_fd_sc_hd__nand3_1 _38014_ (.A(net665),
    .B(net755),
    .C(_11014_),
    .Y(_16659_));
 sky130_fd_sc_hd__a21oi_4 _38015_ (.A1(_16658_),
    .A2(_16659_),
    .B1(net2955),
    .Y(_04549_));
 sky130_fd_sc_hd__nor2_1 _38016_ (.A(\inst$top.soc.cpu.sink__payload$12[162] ),
    .B(net672),
    .Y(_16660_));
 sky130_fd_sc_hd__o21ai_1 _38017_ (.A1(\inst$top.soc.cpu.d_branch_target[2] ),
    .A2(net623),
    .B1(net2029),
    .Y(_16661_));
 sky130_fd_sc_hd__nor2_4 _38018_ (.A(_16660_),
    .B(_16661_),
    .Y(_04550_));
 sky130_fd_sc_hd__nor2_1 _38020_ (.A(\inst$top.soc.cpu.sink__payload$12[163] ),
    .B(net673),
    .Y(_16663_));
 sky130_fd_sc_hd__o21ai_1 _38022_ (.A1(\inst$top.soc.cpu.d_branch_target[3] ),
    .A2(net623),
    .B1(net2036),
    .Y(_16665_));
 sky130_fd_sc_hd__nor2_4 _38023_ (.A(_16663_),
    .B(_16665_),
    .Y(_04551_));
 sky130_fd_sc_hd__nor2_1 _38024_ (.A(\inst$top.soc.cpu.sink__payload$12[164] ),
    .B(net672),
    .Y(_16666_));
 sky130_fd_sc_hd__o21ai_1 _38025_ (.A1(_12573_),
    .A2(net623),
    .B1(net2029),
    .Y(_16667_));
 sky130_fd_sc_hd__nor2_4 _38026_ (.A(_16666_),
    .B(_16667_),
    .Y(_04552_));
 sky130_fd_sc_hd__nor2_1 _38027_ (.A(\inst$top.soc.cpu.sink__payload$12[165] ),
    .B(net673),
    .Y(_16668_));
 sky130_fd_sc_hd__nand2_1 _38028_ (.A(net669),
    .B(_12588_),
    .Y(_16669_));
 sky130_fd_sc_hd__nand2_1 _38029_ (.A(_16669_),
    .B(net2038),
    .Y(_16670_));
 sky130_fd_sc_hd__nor2_4 _38030_ (.A(_16668_),
    .B(_16670_),
    .Y(_04553_));
 sky130_fd_sc_hd__nor2_1 _38031_ (.A(\inst$top.soc.cpu.sink__payload$12[166] ),
    .B(net668),
    .Y(_16671_));
 sky130_fd_sc_hd__nand2_1 _38032_ (.A(net668),
    .B(_12602_),
    .Y(_16672_));
 sky130_fd_sc_hd__nand2_1 _38033_ (.A(_16672_),
    .B(net2038),
    .Y(_16673_));
 sky130_fd_sc_hd__nor2_4 _38034_ (.A(_16671_),
    .B(_16673_),
    .Y(_04554_));
 sky130_fd_sc_hd__nor2_1 _38035_ (.A(\inst$top.soc.cpu.sink__payload$12[167] ),
    .B(net666),
    .Y(_16674_));
 sky130_fd_sc_hd__nand2_1 _38036_ (.A(net666),
    .B(_12616_),
    .Y(_16675_));
 sky130_fd_sc_hd__nand2_1 _38037_ (.A(_16675_),
    .B(net2029),
    .Y(_16676_));
 sky130_fd_sc_hd__nor2_4 _38038_ (.A(_16674_),
    .B(_16676_),
    .Y(_04555_));
 sky130_fd_sc_hd__nor2_1 _38039_ (.A(\inst$top.soc.cpu.sink__payload$12[168] ),
    .B(net679),
    .Y(_16677_));
 sky130_fd_sc_hd__nand2_1 _38040_ (.A(net675),
    .B(_12631_),
    .Y(_16678_));
 sky130_fd_sc_hd__nand2_1 _38042_ (.A(_16678_),
    .B(net2040),
    .Y(_16680_));
 sky130_fd_sc_hd__nor2_4 _38043_ (.A(_16677_),
    .B(_16680_),
    .Y(_04556_));
 sky130_fd_sc_hd__nor2_1 _38044_ (.A(\inst$top.soc.cpu.sink__payload$12[169] ),
    .B(net679),
    .Y(_16681_));
 sky130_fd_sc_hd__nand2_1 _38045_ (.A(net675),
    .B(_12645_),
    .Y(_16682_));
 sky130_fd_sc_hd__nand2_1 _38046_ (.A(_16682_),
    .B(net2040),
    .Y(_16683_));
 sky130_fd_sc_hd__nor2_4 _38047_ (.A(_16681_),
    .B(_16683_),
    .Y(_04557_));
 sky130_fd_sc_hd__nor2_1 _38048_ (.A(\inst$top.soc.cpu.sink__payload$12[16] ),
    .B(net687),
    .Y(_16684_));
 sky130_fd_sc_hd__o21ai_1 _38049_ (.A1(\inst$top.soc.cpu.sink__payload$6[16] ),
    .A2(net643),
    .B1(net2073),
    .Y(_16685_));
 sky130_fd_sc_hd__nor2_4 _38050_ (.A(_16684_),
    .B(_16685_),
    .Y(_04558_));
 sky130_fd_sc_hd__nor2_1 _38051_ (.A(\inst$top.soc.cpu.sink__payload$12[170] ),
    .B(net680),
    .Y(_16686_));
 sky130_fd_sc_hd__o21ai_1 _38052_ (.A1(_12661_),
    .A2(net630),
    .B1(net2067),
    .Y(_16687_));
 sky130_fd_sc_hd__nor2_4 _38053_ (.A(_16686_),
    .B(_16687_),
    .Y(_04559_));
 sky130_fd_sc_hd__nor2_1 _38054_ (.A(\inst$top.soc.cpu.sink__payload$12[171] ),
    .B(net669),
    .Y(_16688_));
 sky130_fd_sc_hd__o21ai_1 _38055_ (.A1(_12677_),
    .A2(net625),
    .B1(net2038),
    .Y(_16689_));
 sky130_fd_sc_hd__nor2_4 _38056_ (.A(_16688_),
    .B(_16689_),
    .Y(_04560_));
 sky130_fd_sc_hd__nor2_1 _38058_ (.A(\inst$top.soc.cpu.sink__payload$12[172] ),
    .B(net679),
    .Y(_16691_));
 sky130_fd_sc_hd__o21ai_1 _38059_ (.A1(_11987_),
    .A2(net629),
    .B1(net2040),
    .Y(_16692_));
 sky130_fd_sc_hd__nor2_4 _38060_ (.A(_16691_),
    .B(_16692_),
    .Y(_04561_));
 sky130_fd_sc_hd__nor2_1 _38061_ (.A(\inst$top.soc.cpu.sink__payload$12[173] ),
    .B(net680),
    .Y(_16693_));
 sky130_fd_sc_hd__o21ai_1 _38062_ (.A1(_12031_),
    .A2(net645),
    .B1(net2068),
    .Y(_16694_));
 sky130_fd_sc_hd__nor2_4 _38063_ (.A(_16693_),
    .B(_16694_),
    .Y(_04562_));
 sky130_fd_sc_hd__nor2_1 _38064_ (.A(\inst$top.soc.cpu.sink__payload$12[174] ),
    .B(net680),
    .Y(_16695_));
 sky130_fd_sc_hd__o21ai_1 _38065_ (.A1(_12054_),
    .A2(net634),
    .B1(net2068),
    .Y(_16696_));
 sky130_fd_sc_hd__nor2_4 _38066_ (.A(_16695_),
    .B(_16696_),
    .Y(_04563_));
 sky130_fd_sc_hd__nor2_1 _38067_ (.A(\inst$top.soc.cpu.sink__payload$12[175] ),
    .B(net680),
    .Y(_16697_));
 sky130_fd_sc_hd__o21ai_1 _38069_ (.A1(_12090_),
    .A2(net637),
    .B1(net2065),
    .Y(_16699_));
 sky130_fd_sc_hd__nor2_4 _38070_ (.A(_16697_),
    .B(_16699_),
    .Y(_04564_));
 sky130_fd_sc_hd__nor2_1 _38071_ (.A(\inst$top.soc.cpu.sink__payload$12[176] ),
    .B(net679),
    .Y(_16700_));
 sky130_fd_sc_hd__nand2_1 _38073_ (.A(net679),
    .B(_12113_),
    .Y(_16702_));
 sky130_fd_sc_hd__nand2_1 _38074_ (.A(_16702_),
    .B(net2044),
    .Y(_16703_));
 sky130_fd_sc_hd__nor2_4 _38075_ (.A(_16700_),
    .B(_16703_),
    .Y(_04565_));
 sky130_fd_sc_hd__nor2_1 _38076_ (.A(\inst$top.soc.cpu.sink__payload$12[177] ),
    .B(net679),
    .Y(_16704_));
 sky130_fd_sc_hd__o21ai_1 _38077_ (.A1(_12144_),
    .A2(net630),
    .B1(net2040),
    .Y(_16705_));
 sky130_fd_sc_hd__nor2_4 _38078_ (.A(_16704_),
    .B(_16705_),
    .Y(_04566_));
 sky130_fd_sc_hd__nor2_1 _38079_ (.A(\inst$top.soc.cpu.sink__payload$12[178] ),
    .B(net668),
    .Y(_16706_));
 sky130_fd_sc_hd__o21ai_1 _38081_ (.A1(_12168_),
    .A2(net623),
    .B1(net2030),
    .Y(_16708_));
 sky130_fd_sc_hd__nor2_4 _38082_ (.A(_16706_),
    .B(_16708_),
    .Y(_04567_));
 sky130_fd_sc_hd__nor2_1 _38083_ (.A(\inst$top.soc.cpu.sink__payload$12[179] ),
    .B(net666),
    .Y(_16709_));
 sky130_fd_sc_hd__nand2_1 _38084_ (.A(net666),
    .B(_12194_),
    .Y(_16710_));
 sky130_fd_sc_hd__nand2_1 _38085_ (.A(_16710_),
    .B(net2036),
    .Y(_16711_));
 sky130_fd_sc_hd__nor2_4 _38086_ (.A(_16709_),
    .B(_16711_),
    .Y(_04568_));
 sky130_fd_sc_hd__nor2_1 _38087_ (.A(\inst$top.soc.cpu.sink__payload$12[17] ),
    .B(net682),
    .Y(_16712_));
 sky130_fd_sc_hd__o21ai_1 _38088_ (.A1(\inst$top.soc.cpu.sink__payload$6[17] ),
    .A2(net638),
    .B1(net2073),
    .Y(_16713_));
 sky130_fd_sc_hd__nor2_4 _38089_ (.A(_16712_),
    .B(_16713_),
    .Y(_04569_));
 sky130_fd_sc_hd__nor2_1 _38090_ (.A(\inst$top.soc.cpu.sink__payload$12[180] ),
    .B(net673),
    .Y(_16714_));
 sky130_fd_sc_hd__o21ai_1 _38091_ (.A1(_12238_),
    .A2(net629),
    .B1(net2037),
    .Y(_16715_));
 sky130_fd_sc_hd__nor2_4 _38092_ (.A(_16714_),
    .B(_16715_),
    .Y(_04570_));
 sky130_fd_sc_hd__nor2_1 _38095_ (.A(\inst$top.soc.cpu.sink__payload$12[181] ),
    .B(net669),
    .Y(_16718_));
 sky130_fd_sc_hd__o21ai_1 _38096_ (.A1(_12261_),
    .A2(net629),
    .B1(net2039),
    .Y(_16719_));
 sky130_fd_sc_hd__nor2_4 _38097_ (.A(_16718_),
    .B(_16719_),
    .Y(_04571_));
 sky130_fd_sc_hd__nor2_1 _38098_ (.A(\inst$top.soc.cpu.sink__payload$12[182] ),
    .B(net681),
    .Y(_16720_));
 sky130_fd_sc_hd__o21ai_1 _38099_ (.A1(_12298_),
    .A2(net637),
    .B1(net2067),
    .Y(_16721_));
 sky130_fd_sc_hd__nor2_4 _38100_ (.A(_16720_),
    .B(_16721_),
    .Y(_04572_));
 sky130_fd_sc_hd__nor2_1 _38101_ (.A(\inst$top.soc.cpu.sink__payload$12[183] ),
    .B(net678),
    .Y(_16722_));
 sky130_fd_sc_hd__nand2_1 _38102_ (.A(net678),
    .B(_12325_),
    .Y(_16723_));
 sky130_fd_sc_hd__nand2_1 _38103_ (.A(_16723_),
    .B(net2065),
    .Y(_16724_));
 sky130_fd_sc_hd__nor2_4 _38104_ (.A(_16722_),
    .B(_16724_),
    .Y(_04573_));
 sky130_fd_sc_hd__nor2_1 _38105_ (.A(\inst$top.soc.cpu.sink__payload$12[184] ),
    .B(net678),
    .Y(_16725_));
 sky130_fd_sc_hd__nand2_1 _38106_ (.A(net678),
    .B(_12349_),
    .Y(_16726_));
 sky130_fd_sc_hd__nand2_1 _38107_ (.A(_16726_),
    .B(net2065),
    .Y(_16727_));
 sky130_fd_sc_hd__nor2_4 _38108_ (.A(_16725_),
    .B(_16727_),
    .Y(_04574_));
 sky130_fd_sc_hd__nor2_1 _38109_ (.A(\inst$top.soc.cpu.sink__payload$12[185] ),
    .B(net666),
    .Y(_16728_));
 sky130_fd_sc_hd__nand2_1 _38110_ (.A(net666),
    .B(_12378_),
    .Y(_16729_));
 sky130_fd_sc_hd__nand2_1 _38111_ (.A(_16729_),
    .B(net2030),
    .Y(_16730_));
 sky130_fd_sc_hd__nor2_4 _38112_ (.A(_16728_),
    .B(_16730_),
    .Y(_04575_));
 sky130_fd_sc_hd__nor2_1 _38113_ (.A(\inst$top.soc.cpu.sink__payload$12[186] ),
    .B(net690),
    .Y(_16731_));
 sky130_fd_sc_hd__nand2_1 _38114_ (.A(net684),
    .B(_12414_),
    .Y(_16732_));
 sky130_fd_sc_hd__nand2_1 _38115_ (.A(_16732_),
    .B(net2066),
    .Y(_16733_));
 sky130_fd_sc_hd__nor2_4 _38116_ (.A(_16731_),
    .B(_16733_),
    .Y(_04576_));
 sky130_fd_sc_hd__nor2_1 _38117_ (.A(\inst$top.soc.cpu.sink__payload$12[187] ),
    .B(net682),
    .Y(_16734_));
 sky130_fd_sc_hd__nand2_1 _38118_ (.A(net682),
    .B(_12447_),
    .Y(_16735_));
 sky130_fd_sc_hd__nand2_1 _38119_ (.A(_16735_),
    .B(net2073),
    .Y(_16736_));
 sky130_fd_sc_hd__nor2_4 _38120_ (.A(_16734_),
    .B(_16736_),
    .Y(_04577_));
 sky130_fd_sc_hd__nor2_1 _38121_ (.A(\inst$top.soc.cpu.sink__payload$12[188] ),
    .B(net684),
    .Y(_16737_));
 sky130_fd_sc_hd__nand2_1 _38122_ (.A(net684),
    .B(_12475_),
    .Y(_16738_));
 sky130_fd_sc_hd__nand2_1 _38123_ (.A(_16738_),
    .B(net2065),
    .Y(_16739_));
 sky130_fd_sc_hd__nor2_4 _38124_ (.A(_16737_),
    .B(_16739_),
    .Y(_04578_));
 sky130_fd_sc_hd__nor2_1 _38125_ (.A(\inst$top.soc.cpu.sink__payload$12[189] ),
    .B(net684),
    .Y(_16740_));
 sky130_fd_sc_hd__nand2_1 _38126_ (.A(net677),
    .B(_12501_),
    .Y(_16741_));
 sky130_fd_sc_hd__nand2_1 _38127_ (.A(_16741_),
    .B(net2065),
    .Y(_16742_));
 sky130_fd_sc_hd__nor2_4 _38128_ (.A(_16740_),
    .B(_16742_),
    .Y(_04579_));
 sky130_fd_sc_hd__nor2_1 _38129_ (.A(\inst$top.soc.cpu.sink__payload$12[18] ),
    .B(net669),
    .Y(_16743_));
 sky130_fd_sc_hd__o21ai_1 _38130_ (.A1(\inst$top.soc.cpu.sink__payload$6[18] ),
    .A2(net625),
    .B1(net2037),
    .Y(_16744_));
 sky130_fd_sc_hd__nor2_4 _38131_ (.A(_16743_),
    .B(_16744_),
    .Y(_04580_));
 sky130_fd_sc_hd__nor2_1 _38133_ (.A(\inst$top.soc.cpu.sink__payload$12[190] ),
    .B(net684),
    .Y(_16746_));
 sky130_fd_sc_hd__nand2_1 _38134_ (.A(net684),
    .B(_12526_),
    .Y(_16747_));
 sky130_fd_sc_hd__nand2_1 _38135_ (.A(_16747_),
    .B(net2065),
    .Y(_16748_));
 sky130_fd_sc_hd__nor2_4 _38136_ (.A(_16746_),
    .B(_16748_),
    .Y(_04581_));
 sky130_fd_sc_hd__nor2_1 _38137_ (.A(\inst$top.soc.cpu.sink__payload$12[191] ),
    .B(net666),
    .Y(_16749_));
 sky130_fd_sc_hd__o21ai_1 _38138_ (.A1(_12551_),
    .A2(net623),
    .B1(net2029),
    .Y(_16750_));
 sky130_fd_sc_hd__nor2_4 _38139_ (.A(_16749_),
    .B(_16750_),
    .Y(_04582_));
 sky130_fd_sc_hd__nor2_1 _38140_ (.A(\inst$top.soc.cpu.d.sink__payload.branch_predict_taken ),
    .B(net673),
    .Y(_16751_));
 sky130_fd_sc_hd__o21ai_1 _38141_ (.A1(net831),
    .A2(net633),
    .B1(net2033),
    .Y(_16752_));
 sky130_fd_sc_hd__nor2_4 _38142_ (.A(_16751_),
    .B(_16752_),
    .Y(_04583_));
 sky130_fd_sc_hd__nor4_1 _38143_ (.A(net2821),
    .B(net2820),
    .C(_16052_),
    .D(_20299_),
    .Y(_16753_));
 sky130_fd_sc_hd__nand2_1 _38145_ (.A(net637),
    .B(_20361_),
    .Y(_16755_));
 sky130_fd_sc_hd__o21ai_1 _38146_ (.A1(_16753_),
    .A2(net637),
    .B1(_16755_),
    .Y(_16756_));
 sky130_fd_sc_hd__nor2_4 _38147_ (.A(net2955),
    .B(_16756_),
    .Y(_04584_));
 sky130_fd_sc_hd__nand2_1 _38148_ (.A(net653),
    .B(net2850),
    .Y(_16757_));
 sky130_fd_sc_hd__nand3_1 _38149_ (.A(net665),
    .B(_20354_),
    .C(net755),
    .Y(_16758_));
 sky130_fd_sc_hd__a21oi_4 _38151_ (.A1(_16757_),
    .A2(_16758_),
    .B1(net2993),
    .Y(_04585_));
 sky130_fd_sc_hd__nand2_1 _38152_ (.A(net641),
    .B(\inst$top.soc.cpu.d.sink__payload.csr_we ),
    .Y(_16760_));
 sky130_fd_sc_hd__a21oi_1 _38153_ (.A1(\inst$top.soc.cpu.sink__payload$6[45] ),
    .A2(_20347_),
    .B1(_16580_),
    .Y(_16761_));
 sky130_fd_sc_hd__nand3_1 _38154_ (.A(net665),
    .B(net755),
    .C(_16761_),
    .Y(_16762_));
 sky130_fd_sc_hd__a21oi_4 _38155_ (.A1(_16760_),
    .A2(_16762_),
    .B1(net2955),
    .Y(_04586_));
 sky130_fd_sc_hd__nor2_1 _38156_ (.A(net2842),
    .B(net686),
    .Y(_16763_));
 sky130_fd_sc_hd__o21ai_1 _38157_ (.A1(net2820),
    .A2(net639),
    .B1(net2076),
    .Y(_16764_));
 sky130_fd_sc_hd__nor2_4 _38158_ (.A(_16763_),
    .B(_16764_),
    .Y(_04587_));
 sky130_fd_sc_hd__nand2_1 _38159_ (.A(net653),
    .B(\inst$top.soc.cpu.d.sink__payload.csr_set ),
    .Y(_16765_));
 sky130_fd_sc_hd__nor2_1 _38160_ (.A(\inst$top.soc.cpu.sink__payload$6[44] ),
    .B(_16476_),
    .Y(_16766_));
 sky130_fd_sc_hd__nand3_1 _38161_ (.A(net665),
    .B(_16766_),
    .C(net755),
    .Y(_16767_));
 sky130_fd_sc_hd__a21oi_4 _38162_ (.A1(_16765_),
    .A2(_16767_),
    .B1(net2993),
    .Y(_04588_));
 sky130_fd_sc_hd__nor2_1 _38163_ (.A(\inst$top.soc.cpu.d.sink__payload.csr_clear ),
    .B(net692),
    .Y(_16768_));
 sky130_fd_sc_hd__o21ai_1 _38164_ (.A1(_16046_),
    .A2(net653),
    .B1(net2080),
    .Y(_16769_));
 sky130_fd_sc_hd__nor2_4 _38165_ (.A(_16768_),
    .B(_16769_),
    .Y(_04589_));
 sky130_fd_sc_hd__nor2_1 _38166_ (.A(\inst$top.soc.cpu.d.sink__payload.ecall ),
    .B(net692),
    .Y(_16770_));
 sky130_fd_sc_hd__nor2_1 _38167_ (.A(\inst$top.soc.cpu.sink__payload$6[57] ),
    .B(_16591_),
    .Y(_16771_));
 sky130_fd_sc_hd__nand3_1 _38168_ (.A(_16771_),
    .B(net2450),
    .C(net2496),
    .Y(_16772_));
 sky130_fd_sc_hd__nor2_1 _38169_ (.A(_16041_),
    .B(_20295_),
    .Y(_16773_));
 sky130_fd_sc_hd__inv_1 _38170_ (.A(_16773_),
    .Y(_16774_));
 sky130_fd_sc_hd__nor4_1 _38171_ (.A(_20236_),
    .B(_16772_),
    .C(_16593_),
    .D(_16774_),
    .Y(_16775_));
 sky130_fd_sc_hd__o21ai_1 _38173_ (.A1(_16775_),
    .A2(net644),
    .B1(net2080),
    .Y(_16777_));
 sky130_fd_sc_hd__nor2_4 _38174_ (.A(_16770_),
    .B(_16777_),
    .Y(_04590_));
 sky130_fd_sc_hd__nor2_1 _38175_ (.A(\inst$top.soc.cpu.sink__payload$12[19] ),
    .B(net683),
    .Y(_16778_));
 sky130_fd_sc_hd__o21ai_1 _38176_ (.A1(\inst$top.soc.cpu.sink__payload$6[19] ),
    .A2(net642),
    .B1(net2073),
    .Y(_16779_));
 sky130_fd_sc_hd__nor2_4 _38177_ (.A(_16778_),
    .B(_16779_),
    .Y(_04591_));
 sky130_fd_sc_hd__nor2_1 _38178_ (.A(\inst$top.soc.cpu.d.sink__payload.ebreak ),
    .B(net690),
    .Y(_16780_));
 sky130_fd_sc_hd__inv_1 _38179_ (.A(net1947),
    .Y(_16781_));
 sky130_fd_sc_hd__nor4_1 _38180_ (.A(_16781_),
    .B(_16772_),
    .C(_16593_),
    .D(_16774_),
    .Y(_16782_));
 sky130_fd_sc_hd__o21ai_1 _38181_ (.A1(_16782_),
    .A2(net644),
    .B1(net2078),
    .Y(_16783_));
 sky130_fd_sc_hd__nor2_4 _38182_ (.A(_16780_),
    .B(_16783_),
    .Y(_04592_));
 sky130_fd_sc_hd__nor2_1 _38183_ (.A(\inst$top.soc.cpu.d.sink__payload.mret ),
    .B(net690),
    .Y(_16784_));
 sky130_fd_sc_hd__nor2_1 _38184_ (.A(\inst$top.soc.cpu.sink__payload$6[63] ),
    .B(\inst$top.soc.cpu.sink__payload$6[62] ),
    .Y(_16785_));
 sky130_fd_sc_hd__nand4_1 _38185_ (.A(_16785_),
    .B(net2620),
    .C(net2465),
    .D(\inst$top.soc.cpu.sink__payload$6[61] ),
    .Y(_16786_));
 sky130_fd_sc_hd__nand2_1 _38186_ (.A(_16773_),
    .B(\inst$top.soc.cpu.sink__payload$6[60] ),
    .Y(_16787_));
 sky130_fd_sc_hd__or3_1 _38187_ (.A(_16772_),
    .B(_16786_),
    .C(_16787_),
    .X(_16788_));
 sky130_fd_sc_hd__nand2_1 _38188_ (.A(net690),
    .B(_16788_),
    .Y(_16789_));
 sky130_fd_sc_hd__nand2_1 _38189_ (.A(_16789_),
    .B(net2078),
    .Y(_16790_));
 sky130_fd_sc_hd__nor2_4 _38190_ (.A(_16784_),
    .B(_16790_),
    .Y(_04593_));
 sky130_fd_sc_hd__nor2_1 _38191_ (.A(\inst$top.soc.cpu.sink__payload$12[20] ),
    .B(net667),
    .Y(_16791_));
 sky130_fd_sc_hd__o21ai_1 _38192_ (.A1(\inst$top.soc.cpu.sink__payload$6[20] ),
    .A2(net623),
    .B1(net2030),
    .Y(_16792_));
 sky130_fd_sc_hd__nor2_4 _38193_ (.A(_16791_),
    .B(_16792_),
    .Y(_04594_));
 sky130_fd_sc_hd__nor2_1 _38195_ (.A(\inst$top.soc.cpu.sink__payload$12[21] ),
    .B(net669),
    .Y(_16794_));
 sky130_fd_sc_hd__o21ai_1 _38196_ (.A1(\inst$top.soc.cpu.sink__payload$6[21] ),
    .A2(net629),
    .B1(net2037),
    .Y(_16795_));
 sky130_fd_sc_hd__nor2_4 _38197_ (.A(_16794_),
    .B(_16795_),
    .Y(_04595_));
 sky130_fd_sc_hd__nor2_1 _38198_ (.A(\inst$top.soc.cpu.sink__payload$12[22] ),
    .B(net686),
    .Y(_16796_));
 sky130_fd_sc_hd__o21ai_1 _38199_ (.A1(\inst$top.soc.cpu.sink__payload$6[22] ),
    .A2(net639),
    .B1(net2073),
    .Y(_16797_));
 sky130_fd_sc_hd__nor2_4 _38200_ (.A(_16796_),
    .B(_16797_),
    .Y(_04596_));
 sky130_fd_sc_hd__nor2_1 _38201_ (.A(\inst$top.soc.cpu.sink__payload$12[23] ),
    .B(net683),
    .Y(_16798_));
 sky130_fd_sc_hd__o21ai_1 _38202_ (.A1(\inst$top.soc.cpu.sink__payload$6[23] ),
    .A2(net637),
    .B1(net2065),
    .Y(_16799_));
 sky130_fd_sc_hd__nor2_4 _38203_ (.A(_16798_),
    .B(_16799_),
    .Y(_04597_));
 sky130_fd_sc_hd__nor2_1 _38204_ (.A(\inst$top.soc.cpu.sink__payload$12[24] ),
    .B(net683),
    .Y(_16800_));
 sky130_fd_sc_hd__o21ai_1 _38206_ (.A1(\inst$top.soc.cpu.sink__payload$6[24] ),
    .A2(net637),
    .B1(net2066),
    .Y(_16802_));
 sky130_fd_sc_hd__nor2_4 _38207_ (.A(_16800_),
    .B(_16802_),
    .Y(_04598_));
 sky130_fd_sc_hd__nor2_1 _38208_ (.A(\inst$top.soc.cpu.sink__payload$12[25] ),
    .B(net683),
    .Y(_16803_));
 sky130_fd_sc_hd__o21ai_1 _38209_ (.A1(\inst$top.soc.cpu.sink__payload$6[25] ),
    .A2(net642),
    .B1(net2073),
    .Y(_16804_));
 sky130_fd_sc_hd__nor2_4 _38210_ (.A(_16803_),
    .B(_16804_),
    .Y(_04599_));
 sky130_fd_sc_hd__nor2_1 _38211_ (.A(\inst$top.soc.cpu.sink__payload$12[26] ),
    .B(net687),
    .Y(_16805_));
 sky130_fd_sc_hd__o21ai_1 _38212_ (.A1(\inst$top.soc.cpu.sink__payload$6[26] ),
    .A2(net642),
    .B1(net2073),
    .Y(_16806_));
 sky130_fd_sc_hd__nor2_4 _38213_ (.A(_16805_),
    .B(_16806_),
    .Y(_04600_));
 sky130_fd_sc_hd__nor2_1 _38214_ (.A(\inst$top.soc.cpu.sink__payload$12[27] ),
    .B(net683),
    .Y(_16807_));
 sky130_fd_sc_hd__o21ai_1 _38216_ (.A1(\inst$top.soc.cpu.sink__payload$6[27] ),
    .A2(net642),
    .B1(net2075),
    .Y(_16809_));
 sky130_fd_sc_hd__nor2_4 _38217_ (.A(_16807_),
    .B(_16809_),
    .Y(_04601_));
 sky130_fd_sc_hd__nor2_1 _38218_ (.A(\inst$top.soc.cpu.sink__payload$12[28] ),
    .B(net683),
    .Y(_16810_));
 sky130_fd_sc_hd__o21ai_1 _38219_ (.A1(\inst$top.soc.cpu.sink__payload$6[28] ),
    .A2(net642),
    .B1(net2075),
    .Y(_16811_));
 sky130_fd_sc_hd__nor2_4 _38220_ (.A(_16810_),
    .B(_16811_),
    .Y(_04602_));
 sky130_fd_sc_hd__nor2_1 _38221_ (.A(\inst$top.soc.cpu.sink__payload$12[29] ),
    .B(net683),
    .Y(_16812_));
 sky130_fd_sc_hd__o21ai_1 _38222_ (.A1(\inst$top.soc.cpu.sink__payload$6[29] ),
    .A2(net642),
    .B1(net2073),
    .Y(_16813_));
 sky130_fd_sc_hd__nor2_4 _38223_ (.A(_16812_),
    .B(_16813_),
    .Y(_04603_));
 sky130_fd_sc_hd__nor2_1 _38224_ (.A(\inst$top.soc.cpu.sink__payload$12[2] ),
    .B(net672),
    .Y(_16814_));
 sky130_fd_sc_hd__o21ai_1 _38225_ (.A1(\inst$top.soc.cpu.sink__payload$6[2] ),
    .A2(net624),
    .B1(net2029),
    .Y(_16815_));
 sky130_fd_sc_hd__nor2_4 _38226_ (.A(_16814_),
    .B(_16815_),
    .Y(_04604_));
 sky130_fd_sc_hd__nor2_1 _38228_ (.A(\inst$top.soc.cpu.sink__payload$12[30] ),
    .B(net684),
    .Y(_16817_));
 sky130_fd_sc_hd__o21ai_1 _38229_ (.A1(\inst$top.soc.cpu.sink__payload$6[30] ),
    .A2(net642),
    .B1(net2074),
    .Y(_16818_));
 sky130_fd_sc_hd__nor2_4 _38230_ (.A(_16817_),
    .B(_16818_),
    .Y(_04605_));
 sky130_fd_sc_hd__nor2_1 _38231_ (.A(\inst$top.soc.cpu.sink__payload$12[31] ),
    .B(net685),
    .Y(_16819_));
 sky130_fd_sc_hd__o21ai_1 _38232_ (.A1(\inst$top.soc.cpu.sink__payload$6[31] ),
    .A2(net641),
    .B1(net2074),
    .Y(_16820_));
 sky130_fd_sc_hd__nor2_4 _38233_ (.A(_16819_),
    .B(_16820_),
    .Y(_04606_));
 sky130_fd_sc_hd__nor2_1 _38234_ (.A(\inst$top.soc.cpu.sink__payload$12[32] ),
    .B(net690),
    .Y(_16821_));
 sky130_fd_sc_hd__o21ai_1 _38235_ (.A1(\inst$top.soc.cpu.sink__payload$6[32] ),
    .A2(net644),
    .B1(net2078),
    .Y(_16822_));
 sky130_fd_sc_hd__nor2_4 _38236_ (.A(_16821_),
    .B(_16822_),
    .Y(_04607_));
 sky130_fd_sc_hd__nor2_1 _38237_ (.A(\inst$top.soc.cpu.sink__payload$12[33] ),
    .B(net679),
    .Y(_16823_));
 sky130_fd_sc_hd__o21ai_1 _38239_ (.A1(\inst$top.soc.cpu.sink__payload$6[33] ),
    .A2(net634),
    .B1(net2044),
    .Y(_16825_));
 sky130_fd_sc_hd__nor2_4 _38240_ (.A(_16823_),
    .B(_16825_),
    .Y(_04608_));
 sky130_fd_sc_hd__nor2_1 _38241_ (.A(\inst$top.soc.cpu.sink__payload$12[34] ),
    .B(net668),
    .Y(_16826_));
 sky130_fd_sc_hd__o21ai_2 _38242_ (.A1(\inst$top.soc.cpu.sink__payload$6[34] ),
    .A2(net641),
    .B1(net2074),
    .Y(_16827_));
 sky130_fd_sc_hd__nor2_4 _38243_ (.A(_16826_),
    .B(_16827_),
    .Y(_04609_));
 sky130_fd_sc_hd__nor2_1 _38244_ (.A(\inst$top.soc.cpu.sink__payload$12[35] ),
    .B(net668),
    .Y(_16828_));
 sky130_fd_sc_hd__o21ai_4 _38245_ (.A1(\inst$top.soc.cpu.sink__payload$6[35] ),
    .A2(net646),
    .B1(net2077),
    .Y(_16829_));
 sky130_fd_sc_hd__nor2_4 _38246_ (.A(_16828_),
    .B(_16829_),
    .Y(_04610_));
 sky130_fd_sc_hd__nor2_1 _38247_ (.A(\inst$top.soc.cpu.sink__payload$12[36] ),
    .B(net680),
    .Y(_16830_));
 sky130_fd_sc_hd__o21ai_1 _38250_ (.A1(\inst$top.soc.cpu.sink__payload$6[36] ),
    .A2(net641),
    .B1(net2074),
    .Y(_16833_));
 sky130_fd_sc_hd__nor2_4 _38251_ (.A(_16830_),
    .B(_16833_),
    .Y(_04611_));
 sky130_fd_sc_hd__nor2_1 _38252_ (.A(\inst$top.soc.cpu.sink__payload$12[37] ),
    .B(net673),
    .Y(_16834_));
 sky130_fd_sc_hd__o21ai_2 _38253_ (.A1(\inst$top.soc.cpu.sink__payload$6[37] ),
    .A2(net641),
    .B1(net2074),
    .Y(_16835_));
 sky130_fd_sc_hd__nor2_4 _38254_ (.A(_16834_),
    .B(_16835_),
    .Y(_04612_));
 sky130_fd_sc_hd__nor2_1 _38255_ (.A(\inst$top.soc.cpu.sink__payload$12[38] ),
    .B(net673),
    .Y(_16836_));
 sky130_fd_sc_hd__o21ai_2 _38256_ (.A1(net2821),
    .A2(net643),
    .B1(net2077),
    .Y(_16837_));
 sky130_fd_sc_hd__nor2_4 _38257_ (.A(_16836_),
    .B(_16837_),
    .Y(_04613_));
 sky130_fd_sc_hd__nor2_1 _38258_ (.A(\inst$top.soc.cpu.sink__payload$12[3] ),
    .B(net667),
    .Y(_16838_));
 sky130_fd_sc_hd__o21ai_1 _38259_ (.A1(\inst$top.soc.cpu.sink__payload$6[3] ),
    .A2(net624),
    .B1(net2029),
    .Y(_16839_));
 sky130_fd_sc_hd__nor2_4 _38260_ (.A(_16838_),
    .B(_16839_),
    .Y(_04614_));
 sky130_fd_sc_hd__nor2_1 _38262_ (.A(\inst$top.soc.cpu.sink__payload$12[4] ),
    .B(net671),
    .Y(_16841_));
 sky130_fd_sc_hd__o21ai_1 _38263_ (.A1(\inst$top.soc.cpu.sink__payload$6[4] ),
    .A2(net624),
    .B1(net2029),
    .Y(_16842_));
 sky130_fd_sc_hd__nor2_4 _38264_ (.A(_16841_),
    .B(_16842_),
    .Y(_04615_));
 sky130_fd_sc_hd__nor2_1 _38265_ (.A(\inst$top.soc.cpu.sink__payload$12[52] ),
    .B(net673),
    .Y(_16843_));
 sky130_fd_sc_hd__o21ai_1 _38266_ (.A1(net2687),
    .A2(net634),
    .B1(net2097),
    .Y(_16844_));
 sky130_fd_sc_hd__nor2_4 _38267_ (.A(_16843_),
    .B(_16844_),
    .Y(_04616_));
 sky130_fd_sc_hd__nor2_1 _38268_ (.A(\inst$top.soc.cpu.sink__payload$12[53] ),
    .B(net692),
    .Y(_16845_));
 sky130_fd_sc_hd__o21ai_1 _38269_ (.A1(net2620),
    .A2(net645),
    .B1(net2080),
    .Y(_16846_));
 sky130_fd_sc_hd__nor2_4 _38270_ (.A(_16845_),
    .B(_16846_),
    .Y(_04617_));
 sky130_fd_sc_hd__nor2_1 _38271_ (.A(\inst$top.soc.cpu.sink__payload$12[54] ),
    .B(net702),
    .Y(_16847_));
 sky130_fd_sc_hd__o21ai_1 _38273_ (.A1(net2608),
    .A2(net655),
    .B1(net2178),
    .Y(_16849_));
 sky130_fd_sc_hd__nor2_4 _38274_ (.A(_16847_),
    .B(_16849_),
    .Y(_04618_));
 sky130_fd_sc_hd__nor2_1 _38275_ (.A(\inst$top.soc.cpu.sink__payload$12[55] ),
    .B(net691),
    .Y(_16850_));
 sky130_fd_sc_hd__o21ai_1 _38276_ (.A1(net2597),
    .A2(net645),
    .B1(net2107),
    .Y(_16851_));
 sky130_fd_sc_hd__nor2_4 _38277_ (.A(_16850_),
    .B(_16851_),
    .Y(_04619_));
 sky130_fd_sc_hd__nor2_1 _38278_ (.A(\inst$top.soc.cpu.sink__payload$12[56] ),
    .B(net691),
    .Y(_16852_));
 sky130_fd_sc_hd__o21ai_1 _38279_ (.A1(net2590),
    .A2(net645),
    .B1(net2111),
    .Y(_16853_));
 sky130_fd_sc_hd__nor2_4 _38280_ (.A(_16852_),
    .B(_16853_),
    .Y(_04620_));
 sky130_fd_sc_hd__nor2_1 _38281_ (.A(\inst$top.soc.cpu.sink__payload$12[57] ),
    .B(net671),
    .Y(_16854_));
 sky130_fd_sc_hd__o21ai_4 _38283_ (.A1(\inst$top.soc.cpu.sink__payload$6[57] ),
    .A2(net645),
    .B1(net2075),
    .Y(_16856_));
 sky130_fd_sc_hd__nor2_4 _38284_ (.A(_16854_),
    .B(_16856_),
    .Y(_04621_));
 sky130_fd_sc_hd__nor2_1 _38285_ (.A(\inst$top.soc.cpu.sink__payload$12[58] ),
    .B(net691),
    .Y(_16857_));
 sky130_fd_sc_hd__o21ai_1 _38286_ (.A1(\inst$top.soc.cpu.sink__payload$6[58] ),
    .A2(net642),
    .B1(net2075),
    .Y(_16858_));
 sky130_fd_sc_hd__nor2_4 _38287_ (.A(_16857_),
    .B(_16858_),
    .Y(_04622_));
 sky130_fd_sc_hd__nor2_1 _38288_ (.A(\inst$top.soc.cpu.sink__payload$12[59] ),
    .B(net690),
    .Y(_16859_));
 sky130_fd_sc_hd__o21ai_1 _38289_ (.A1(\inst$top.soc.cpu.sink__payload$6[59] ),
    .A2(net641),
    .B1(net2075),
    .Y(_16860_));
 sky130_fd_sc_hd__nor2_4 _38290_ (.A(_16859_),
    .B(_16860_),
    .Y(_04623_));
 sky130_fd_sc_hd__nor2_1 _38291_ (.A(\inst$top.soc.cpu.sink__payload$12[5] ),
    .B(net679),
    .Y(_16861_));
 sky130_fd_sc_hd__o21ai_1 _38292_ (.A1(\inst$top.soc.cpu.sink__payload$6[5] ),
    .A2(net630),
    .B1(net2040),
    .Y(_16862_));
 sky130_fd_sc_hd__nor2_4 _38293_ (.A(_16861_),
    .B(_16862_),
    .Y(_04624_));
 sky130_fd_sc_hd__nand2_1 _38294_ (.A(net690),
    .B(\inst$top.soc.cpu.sink__payload$6[60] ),
    .Y(_16863_));
 sky130_fd_sc_hd__nand2_1 _38295_ (.A(net644),
    .B(\inst$top.soc.cpu.sink__payload$12[60] ),
    .Y(_16864_));
 sky130_fd_sc_hd__a21oi_4 _38296_ (.A1(_16863_),
    .A2(_16864_),
    .B1(net2955),
    .Y(_04625_));
 sky130_fd_sc_hd__nor2_1 _38298_ (.A(\inst$top.soc.cpu.sink__payload$12[61] ),
    .B(net690),
    .Y(_16866_));
 sky130_fd_sc_hd__o21ai_1 _38299_ (.A1(\inst$top.soc.cpu.sink__payload$6[61] ),
    .A2(net644),
    .B1(net2078),
    .Y(_16867_));
 sky130_fd_sc_hd__nor2_4 _38300_ (.A(_16866_),
    .B(_16867_),
    .Y(_04626_));
 sky130_fd_sc_hd__nand2_1 _38301_ (.A(net690),
    .B(\inst$top.soc.cpu.sink__payload$6[62] ),
    .Y(_16868_));
 sky130_fd_sc_hd__nand2_1 _38302_ (.A(net644),
    .B(\inst$top.soc.cpu.sink__payload$12[62] ),
    .Y(_16869_));
 sky130_fd_sc_hd__a21oi_4 _38303_ (.A1(_16868_),
    .A2(_16869_),
    .B1(net2955),
    .Y(_04627_));
 sky130_fd_sc_hd__nor2_1 _38304_ (.A(\inst$top.soc.cpu.sink__payload$12[63] ),
    .B(net671),
    .Y(_16870_));
 sky130_fd_sc_hd__o21ai_1 _38305_ (.A1(\inst$top.soc.cpu.sink__payload$6[63] ),
    .A2(net644),
    .B1(net2078),
    .Y(_16871_));
 sky130_fd_sc_hd__nor2_4 _38306_ (.A(_16870_),
    .B(_16871_),
    .Y(_04628_));
 sky130_fd_sc_hd__nor2_1 _38307_ (.A(\inst$top.soc.cpu.sink__payload$12[6] ),
    .B(net679),
    .Y(_16872_));
 sky130_fd_sc_hd__o21ai_1 _38308_ (.A1(\inst$top.soc.cpu.sink__payload$6[6] ),
    .A2(net629),
    .B1(net2040),
    .Y(_16873_));
 sky130_fd_sc_hd__nor2_4 _38309_ (.A(_16872_),
    .B(_16873_),
    .Y(_04629_));
 sky130_fd_sc_hd__nor2_1 _38310_ (.A(\inst$top.soc.cpu.sink__payload$12[7] ),
    .B(net681),
    .Y(_16874_));
 sky130_fd_sc_hd__o21ai_1 _38312_ (.A1(\inst$top.soc.cpu.sink__payload$6[7] ),
    .A2(net637),
    .B1(net2065),
    .Y(_16876_));
 sky130_fd_sc_hd__nor2_4 _38313_ (.A(_16874_),
    .B(_16876_),
    .Y(_04630_));
 sky130_fd_sc_hd__nor2_1 _38314_ (.A(\inst$top.soc.cpu.sink__payload$12[8] ),
    .B(net680),
    .Y(_16877_));
 sky130_fd_sc_hd__o21ai_1 _38315_ (.A1(\inst$top.soc.cpu.sink__payload$6[8] ),
    .A2(net630),
    .B1(net2041),
    .Y(_16878_));
 sky130_fd_sc_hd__nor2_4 _38316_ (.A(_16877_),
    .B(_16878_),
    .Y(_04631_));
 sky130_fd_sc_hd__nor2_1 _38317_ (.A(\inst$top.soc.cpu.d.sink__payload.illegal ),
    .B(net691),
    .Y(_16879_));
 sky130_fd_sc_hd__nor4_1 _38318_ (.A(_16781_),
    .B(_16772_),
    .C(_16593_),
    .D(_16774_),
    .Y(_16880_));
 sky130_fd_sc_hd__nor3_1 _38319_ (.A(\inst$top.soc.cpu.sink__payload$6[61] ),
    .B(net2590),
    .C(_16781_),
    .Y(_16881_));
 sky130_fd_sc_hd__nand4_1 _38320_ (.A(_16881_),
    .B(net1942),
    .C(_16771_),
    .D(_16785_),
    .Y(_16882_));
 sky130_fd_sc_hd__o21ai_0 _38321_ (.A1(_16787_),
    .A2(_16882_),
    .B1(_16788_),
    .Y(_16883_));
 sky130_fd_sc_hd__nand2_1 _38322_ (.A(_16589_),
    .B(_16596_),
    .Y(_16884_));
 sky130_fd_sc_hd__nor4_1 _38323_ (.A(_16775_),
    .B(_16880_),
    .C(_16883_),
    .D(_16884_),
    .Y(_16885_));
 sky130_fd_sc_hd__nor3_1 _38324_ (.A(_16647_),
    .B(_16631_),
    .C(_16638_),
    .Y(_16886_));
 sky130_fd_sc_hd__inv_1 _38325_ (.A(_16614_),
    .Y(_16887_));
 sky130_fd_sc_hd__nand4_1 _38326_ (.A(_16887_),
    .B(_11910_),
    .C(_16477_),
    .D(_16610_),
    .Y(_16888_));
 sky130_fd_sc_hd__nand2_1 _38327_ (.A(_16579_),
    .B(_16582_),
    .Y(_16889_));
 sky130_fd_sc_hd__nor2_1 _38328_ (.A(_16888_),
    .B(_16889_),
    .Y(_16890_));
 sky130_fd_sc_hd__nand2_1 _38329_ (.A(\inst$top.soc.cpu.sink__payload$6[32] ),
    .B(\inst$top.soc.cpu.sink__payload$6[33] ),
    .Y(_16891_));
 sky130_fd_sc_hd__a41o_1 _38330_ (.A1(_16576_),
    .A2(_16885_),
    .A3(_16886_),
    .A4(_16890_),
    .B1(_16891_),
    .X(_16892_));
 sky130_fd_sc_hd__o21ai_1 _38331_ (.A1(_16892_),
    .A2(net644),
    .B1(net2078),
    .Y(_16893_));
 sky130_fd_sc_hd__nor2_4 _38332_ (.A(_16879_),
    .B(_16893_),
    .Y(_04632_));
 sky130_fd_sc_hd__nor2_1 _38333_ (.A(\inst$top.soc.cpu.sink__payload$12[39] ),
    .B(net697),
    .Y(_16894_));
 sky130_fd_sc_hd__o21ai_1 _38335_ (.A1(\inst$top.soc.cpu.sink__payload$6[39] ),
    .A2(net651),
    .B1(net2143),
    .Y(_16896_));
 sky130_fd_sc_hd__nor2_4 _38336_ (.A(_16894_),
    .B(_16896_),
    .Y(_04633_));
 sky130_fd_sc_hd__nor2_1 _38337_ (.A(\inst$top.soc.cpu.sink__payload$12[40] ),
    .B(net696),
    .Y(_16897_));
 sky130_fd_sc_hd__o21ai_1 _38338_ (.A1(\inst$top.soc.cpu.sink__payload$6[40] ),
    .A2(net650),
    .B1(net2143),
    .Y(_16898_));
 sky130_fd_sc_hd__nor2_4 _38339_ (.A(_16897_),
    .B(_16898_),
    .Y(_04634_));
 sky130_fd_sc_hd__nor2_1 _38340_ (.A(\inst$top.soc.cpu.sink__payload$12[41] ),
    .B(net696),
    .Y(_16899_));
 sky130_fd_sc_hd__o21ai_1 _38341_ (.A1(\inst$top.soc.cpu.sink__payload$6[41] ),
    .A2(net650),
    .B1(net2143),
    .Y(_16900_));
 sky130_fd_sc_hd__nor2_4 _38342_ (.A(_16899_),
    .B(_16900_),
    .Y(_04635_));
 sky130_fd_sc_hd__nor2_1 _38343_ (.A(\inst$top.soc.cpu.sink__payload$12[42] ),
    .B(net693),
    .Y(_16901_));
 sky130_fd_sc_hd__o21ai_1 _38344_ (.A1(\inst$top.soc.cpu.sink__payload$6[42] ),
    .A2(net649),
    .B1(net2143),
    .Y(_16902_));
 sky130_fd_sc_hd__nor2_4 _38345_ (.A(_16901_),
    .B(_16902_),
    .Y(_04636_));
 sky130_fd_sc_hd__nor2_1 _38347_ (.A(\inst$top.soc.cpu.sink__payload$12[9] ),
    .B(net681),
    .Y(_16904_));
 sky130_fd_sc_hd__o21ai_1 _38348_ (.A1(\inst$top.soc.cpu.sink__payload$6[9] ),
    .A2(net630),
    .B1(net2067),
    .Y(_16905_));
 sky130_fd_sc_hd__nor2_4 _38349_ (.A(_16904_),
    .B(_16905_),
    .Y(_04637_));
 sky130_fd_sc_hd__o21ai_0 _38350_ (.A1(\inst$top.soc.cpu.sink__payload$12[40] ),
    .A2(net1914),
    .B1(net2143),
    .Y(_16906_));
 sky130_fd_sc_hd__a21oi_1 _38351_ (.A1(_11885_),
    .A2(net1914),
    .B1(_16906_),
    .Y(_04638_));
 sky130_fd_sc_hd__o21ai_0 _38353_ (.A1(\inst$top.soc.cpu.sink__payload$18[101] ),
    .A2(net2275),
    .B1(net2150),
    .Y(_16908_));
 sky130_fd_sc_hd__a21oi_1 _38354_ (.A1(_20317_),
    .A2(net2275),
    .B1(_16908_),
    .Y(_04639_));
 sky130_fd_sc_hd__o21ai_0 _38355_ (.A1(\inst$top.soc.cpu.sink__payload$12[42] ),
    .A2(net1914),
    .B1(net2150),
    .Y(_16909_));
 sky130_fd_sc_hd__a21oi_1 _38356_ (.A1(_11724_),
    .A2(net1914),
    .B1(_16909_),
    .Y(_04640_));
 sky130_fd_sc_hd__o21ai_0 _38357_ (.A1(\inst$top.soc.cpu.sink__payload$12[100] ),
    .A2(net1914),
    .B1(net2150),
    .Y(_16910_));
 sky130_fd_sc_hd__a21oi_1 _38358_ (.A1(_20271_),
    .A2(net1914),
    .B1(_16910_),
    .Y(_04641_));
 sky130_fd_sc_hd__o21ai_0 _38359_ (.A1(\inst$top.soc.cpu.d.sink__payload$6.rd_we ),
    .A2(net2267),
    .B1(net2144),
    .Y(_16911_));
 sky130_fd_sc_hd__a21oi_1 _38360_ (.A1(_20138_),
    .A2(net2267),
    .B1(_16911_),
    .Y(_04642_));
 sky130_fd_sc_hd__nor3_1 _38362_ (.A(\inst$top.soc.cpu.d.sink__payload.bypass_x ),
    .B(\inst$top.soc.cpu.d.sink__payload.bypass_m ),
    .C(net1914),
    .Y(_16913_));
 sky130_fd_sc_hd__a211oi_1 _38363_ (.A1(_20278_),
    .A2(net1914),
    .B1(net2993),
    .C1(_16913_),
    .Y(_04643_));
 sky130_fd_sc_hd__inv_1 _38364_ (.A(\inst$top.soc.cpu.sink__payload$12[143] ),
    .Y(_16914_));
 sky130_fd_sc_hd__o21ai_0 _38365_ (.A1(\inst$top.soc.cpu.sink__payload$18[106] ),
    .A2(net2277),
    .B1(net2178),
    .Y(_16915_));
 sky130_fd_sc_hd__a21oi_1 _38366_ (.A1(_16914_),
    .A2(net2277),
    .B1(_16915_),
    .Y(_04644_));
 sky130_fd_sc_hd__o21ai_0 _38367_ (.A1(\inst$top.soc.cpu.sink__payload$18[107] ),
    .A2(net2276),
    .B1(net2146),
    .Y(_16916_));
 sky130_fd_sc_hd__a21oi_1 _38368_ (.A1(_09912_),
    .A2(net2276),
    .B1(_16916_),
    .Y(_04645_));
 sky130_fd_sc_hd__o21ai_0 _38369_ (.A1(net2842),
    .A2(net1913),
    .B1(net2141),
    .Y(_16917_));
 sky130_fd_sc_hd__a21oi_1 _38370_ (.A1(_11745_),
    .A2(net1913),
    .B1(_16917_),
    .Y(_04646_));
 sky130_fd_sc_hd__o21ai_0 _38372_ (.A1(\inst$top.soc.cpu.sink__payload$18[109] ),
    .A2(net2276),
    .B1(net2146),
    .Y(_16919_));
 sky130_fd_sc_hd__a21oi_1 _38373_ (.A1(_12982_),
    .A2(net2276),
    .B1(_16919_),
    .Y(_04647_));
 sky130_fd_sc_hd__o21ai_0 _38374_ (.A1(\inst$top.soc.cpu.sink__payload$18[10] ),
    .A2(net2240),
    .B1(net2070),
    .Y(_16920_));
 sky130_fd_sc_hd__a21oi_1 _38375_ (.A1(_20705_),
    .A2(net2240),
    .B1(_16920_),
    .Y(_04648_));
 sky130_fd_sc_hd__o21ai_0 _38376_ (.A1(\inst$top.soc.cpu.sink__payload$18[110] ),
    .A2(net2278),
    .B1(net2148),
    .Y(_16921_));
 sky130_fd_sc_hd__a21oi_1 _38377_ (.A1(_13686_),
    .A2(net2278),
    .B1(_16921_),
    .Y(_04649_));
 sky130_fd_sc_hd__o21ai_0 _38379_ (.A1(\inst$top.soc.cpu.sink__payload$18[111] ),
    .A2(net2276),
    .B1(net2149),
    .Y(_16923_));
 sky130_fd_sc_hd__a21oi_1 _38380_ (.A1(_14261_),
    .A2(net2276),
    .B1(_16923_),
    .Y(_04650_));
 sky130_fd_sc_hd__a21oi_1 _38382_ (.A1(net1916),
    .A2(_14377_),
    .B1(net2993),
    .Y(_16925_));
 sky130_fd_sc_hd__o21ai_0 _38383_ (.A1(net1916),
    .A2(_14376_),
    .B1(_16925_),
    .Y(_16926_));
 sky130_fd_sc_hd__inv_2 _38384_ (.A(_16926_),
    .Y(_04651_));
 sky130_fd_sc_hd__o21ai_0 _38386_ (.A1(\inst$top.soc.cpu.sink__payload$18[113] ),
    .A2(net2277),
    .B1(net2149),
    .Y(_16928_));
 sky130_fd_sc_hd__a21oi_1 _38387_ (.A1(_14413_),
    .A2(net2276),
    .B1(_16928_),
    .Y(_04652_));
 sky130_fd_sc_hd__o21ai_0 _38388_ (.A1(\inst$top.soc.cpu.sink__payload$18[114] ),
    .A2(net2279),
    .B1(net2155),
    .Y(_16929_));
 sky130_fd_sc_hd__a21oi_1 _38389_ (.A1(_14444_),
    .A2(net2279),
    .B1(_16929_),
    .Y(_04653_));
 sky130_fd_sc_hd__o21ai_0 _38390_ (.A1(\inst$top.soc.cpu.sink__payload$18[115] ),
    .A2(net2290),
    .B1(net2172),
    .Y(_16930_));
 sky130_fd_sc_hd__a21oi_1 _38391_ (.A1(_14471_),
    .A2(net2289),
    .B1(_16930_),
    .Y(_04654_));
 sky130_fd_sc_hd__a21oi_1 _38392_ (.A1(net1910),
    .A2(_14493_),
    .B1(net2993),
    .Y(_16931_));
 sky130_fd_sc_hd__o21ai_0 _38393_ (.A1(net1910),
    .A2(net620),
    .B1(_16931_),
    .Y(_16932_));
 sky130_fd_sc_hd__inv_2 _38394_ (.A(_16932_),
    .Y(_04655_));
 sky130_fd_sc_hd__o21ai_0 _38395_ (.A1(\inst$top.soc.cpu.sink__payload$18[117] ),
    .A2(net2289),
    .B1(net2172),
    .Y(_16933_));
 sky130_fd_sc_hd__a21oi_1 _38396_ (.A1(_14530_),
    .A2(net2289),
    .B1(_16933_),
    .Y(_04656_));
 sky130_fd_sc_hd__o21ai_0 _38397_ (.A1(\inst$top.soc.cpu.sink__payload$18[118] ),
    .A2(net2290),
    .B1(net2172),
    .Y(_16934_));
 sky130_fd_sc_hd__a21oi_1 _38398_ (.A1(_14561_),
    .A2(net2289),
    .B1(_16934_),
    .Y(_04657_));
 sky130_fd_sc_hd__o21ai_0 _38399_ (.A1(\inst$top.soc.cpu.sink__payload$18[119] ),
    .A2(net2280),
    .B1(net2155),
    .Y(_16935_));
 sky130_fd_sc_hd__a21oi_1 _38400_ (.A1(_13095_),
    .A2(net2280),
    .B1(_16935_),
    .Y(_04658_));
 sky130_fd_sc_hd__o21ai_0 _38402_ (.A1(\inst$top.soc.cpu.sink__payload$18[11] ),
    .A2(net2230),
    .B1(net2093),
    .Y(_16937_));
 sky130_fd_sc_hd__a21oi_1 _38403_ (.A1(_20726_),
    .A2(net2230),
    .B1(_16937_),
    .Y(_04659_));
 sky130_fd_sc_hd__a21oi_1 _38405_ (.A1(net1917),
    .A2(_13101_),
    .B1(net3006),
    .Y(_16939_));
 sky130_fd_sc_hd__o21ai_0 _38406_ (.A1(net1917),
    .A2(_13190_),
    .B1(_16939_),
    .Y(_16940_));
 sky130_fd_sc_hd__inv_2 _38407_ (.A(_16940_),
    .Y(_04660_));
 sky130_fd_sc_hd__nor2_1 _38409_ (.A(net1924),
    .B(_13228_),
    .Y(_16942_));
 sky130_fd_sc_hd__a211oi_2 _38410_ (.A1(_13229_),
    .A2(net1924),
    .B1(net3004),
    .C1(_16942_),
    .Y(_04661_));
 sky130_fd_sc_hd__nor2_1 _38411_ (.A(net1911),
    .B(net602),
    .Y(_16943_));
 sky130_fd_sc_hd__a211oi_1 _38412_ (.A1(_13246_),
    .A2(net1910),
    .B1(net3005),
    .C1(_16943_),
    .Y(_04662_));
 sky130_fd_sc_hd__o21ai_0 _38413_ (.A1(\inst$top.soc.cpu.sink__payload$18[123] ),
    .A2(net2289),
    .B1(net2172),
    .Y(_16944_));
 sky130_fd_sc_hd__a21oi_1 _38414_ (.A1(_14628_),
    .A2(net2289),
    .B1(_16944_),
    .Y(_04663_));
 sky130_fd_sc_hd__nor2_1 _38415_ (.A(net1915),
    .B(_13387_),
    .Y(_16945_));
 sky130_fd_sc_hd__a211oi_1 _38416_ (.A1(_13388_),
    .A2(net1915),
    .B1(net2994),
    .C1(_16945_),
    .Y(_04664_));
 sky130_fd_sc_hd__a21oi_1 _38417_ (.A1(net1916),
    .A2(_13402_),
    .B1(net3006),
    .Y(_16946_));
 sky130_fd_sc_hd__o21ai_0 _38418_ (.A1(net1916),
    .A2(_13462_),
    .B1(_16946_),
    .Y(_16947_));
 sky130_fd_sc_hd__inv_2 _38419_ (.A(_16947_),
    .Y(_04665_));
 sky130_fd_sc_hd__o21ai_0 _38420_ (.A1(\inst$top.soc.cpu.sink__payload$18[126] ),
    .A2(net2293),
    .B1(net2174),
    .Y(_16948_));
 sky130_fd_sc_hd__a21oi_1 _38421_ (.A1(_14660_),
    .A2(net2293),
    .B1(_16948_),
    .Y(_04666_));
 sky130_fd_sc_hd__o21ai_0 _38423_ (.A1(\inst$top.soc.cpu.sink__payload$18[127] ),
    .A2(net2277),
    .B1(net2178),
    .Y(_16950_));
 sky130_fd_sc_hd__a21oi_1 _38424_ (.A1(_13575_),
    .A2(net2277),
    .B1(_16950_),
    .Y(_04667_));
 sky130_fd_sc_hd__nor2_1 _38425_ (.A(net1910),
    .B(_13660_),
    .Y(_16951_));
 sky130_fd_sc_hd__a211oi_1 _38426_ (.A1(_13593_),
    .A2(net1910),
    .B1(net3005),
    .C1(_16951_),
    .Y(_04668_));
 sky130_fd_sc_hd__nor2_1 _38427_ (.A(net1918),
    .B(_13732_),
    .Y(_16952_));
 sky130_fd_sc_hd__a211oi_1 _38428_ (.A1(_13735_),
    .A2(net1917),
    .B1(net3006),
    .C1(_16952_),
    .Y(_04669_));
 sky130_fd_sc_hd__o21ai_0 _38430_ (.A1(\inst$top.soc.cpu.sink__payload$18[12] ),
    .A2(net2229),
    .B1(net2045),
    .Y(_16954_));
 sky130_fd_sc_hd__a21oi_1 _38431_ (.A1(_20751_),
    .A2(net2229),
    .B1(_16954_),
    .Y(_04670_));
 sky130_fd_sc_hd__nor2_1 _38432_ (.A(net1917),
    .B(_13793_),
    .Y(_16955_));
 sky130_fd_sc_hd__a211oi_1 _38433_ (.A1(_13748_),
    .A2(net1917),
    .B1(net3006),
    .C1(_16955_),
    .Y(_04671_));
 sky130_fd_sc_hd__nor2_1 _38435_ (.A(net1924),
    .B(net603),
    .Y(_16957_));
 sky130_fd_sc_hd__a211oi_2 _38436_ (.A1(_13802_),
    .A2(net1924),
    .B1(net3010),
    .C1(_16957_),
    .Y(_04672_));
 sky130_fd_sc_hd__nor2_1 _38437_ (.A(net1917),
    .B(_13898_),
    .Y(_16958_));
 sky130_fd_sc_hd__a211oi_1 _38438_ (.A1(_13901_),
    .A2(net1917),
    .B1(net3005),
    .C1(_16958_),
    .Y(_04673_));
 sky130_fd_sc_hd__nor2_1 _38439_ (.A(net1916),
    .B(_13947_),
    .Y(_16959_));
 sky130_fd_sc_hd__a211oi_2 _38440_ (.A1(_13950_),
    .A2(net1916),
    .B1(net3006),
    .C1(_16959_),
    .Y(_04674_));
 sky130_fd_sc_hd__nor2_1 _38441_ (.A(net1916),
    .B(_13997_),
    .Y(_16960_));
 sky130_fd_sc_hd__a211oi_2 _38442_ (.A1(_14000_),
    .A2(net1916),
    .B1(net3005),
    .C1(_16960_),
    .Y(_04675_));
 sky130_fd_sc_hd__nor2_1 _38443_ (.A(net1910),
    .B(_14058_),
    .Y(_16961_));
 sky130_fd_sc_hd__a211oi_2 _38444_ (.A1(_14012_),
    .A2(net1912),
    .B1(net3005),
    .C1(_16961_),
    .Y(_04676_));
 sky130_fd_sc_hd__nor2_1 _38445_ (.A(net1910),
    .B(_14118_),
    .Y(_16962_));
 sky130_fd_sc_hd__a211oi_1 _38446_ (.A1(_14066_),
    .A2(net1910),
    .B1(net3005),
    .C1(_16962_),
    .Y(_04677_));
 sky130_fd_sc_hd__nor2_1 _38447_ (.A(net1924),
    .B(_14161_),
    .Y(_16963_));
 sky130_fd_sc_hd__a211oi_2 _38448_ (.A1(_14164_),
    .A2(net1924),
    .B1(net3010),
    .C1(_16963_),
    .Y(_04678_));
 sky130_fd_sc_hd__nor2_1 _38449_ (.A(net1916),
    .B(_14225_),
    .Y(_16964_));
 sky130_fd_sc_hd__a211oi_2 _38450_ (.A1(_14228_),
    .A2(net1916),
    .B1(net3005),
    .C1(_16964_),
    .Y(_04679_));
 sky130_fd_sc_hd__o21ai_0 _38451_ (.A1(\inst$top.soc.cpu.sink__payload$18[139] ),
    .A2(net2284),
    .B1(net2149),
    .Y(_16965_));
 sky130_fd_sc_hd__a21oi_1 _38452_ (.A1(_14313_),
    .A2(net2277),
    .B1(_16965_),
    .Y(_04680_));
 sky130_fd_sc_hd__o21ai_0 _38453_ (.A1(\inst$top.soc.cpu.sink__payload$18[13] ),
    .A2(net2249),
    .B1(net2069),
    .Y(_16966_));
 sky130_fd_sc_hd__a21oi_1 _38454_ (.A1(_20771_),
    .A2(net2239),
    .B1(_16966_),
    .Y(_04681_));
 sky130_fd_sc_hd__o21ai_0 _38455_ (.A1(\inst$top.soc.cpu.sink__payload$18[140] ),
    .A2(net2277),
    .B1(net2146),
    .Y(_16967_));
 sky130_fd_sc_hd__a21oi_1 _38456_ (.A1(_14349_),
    .A2(net2277),
    .B1(_16967_),
    .Y(_04682_));
 sky130_fd_sc_hd__nor2_1 _38457_ (.A(\inst$top.soc.cpu.d.sink__payload.shift ),
    .B(net1913),
    .Y(_16968_));
 sky130_fd_sc_hd__o21ai_0 _38458_ (.A1(net2834),
    .A2(net2276),
    .B1(net2146),
    .Y(_16969_));
 sky130_fd_sc_hd__nor2_1 _38459_ (.A(_16968_),
    .B(_16969_),
    .Y(_04683_));
 sky130_fd_sc_hd__o21ai_0 _38460_ (.A1(\inst$top.soc.cpu.d.sink__payload.load ),
    .A2(net1903),
    .B1(net2075),
    .Y(_16970_));
 sky130_fd_sc_hd__a21oi_1 _38461_ (.A1(_20187_),
    .A2(net1903),
    .B1(_16970_),
    .Y(_04684_));
 sky130_fd_sc_hd__nand2_1 _38462_ (.A(net1903),
    .B(\inst$top.soc.cpu.d.sink__payload$6.store ),
    .Y(_16971_));
 sky130_fd_sc_hd__nand2_1 _38463_ (.A(net2238),
    .B(\inst$top.soc.cpu.d.sink__payload.store ),
    .Y(_16972_));
 sky130_fd_sc_hd__a21oi_1 _38464_ (.A1(_16971_),
    .A2(_16972_),
    .B1(net2955),
    .Y(_04685_));
 sky130_fd_sc_hd__o21ai_0 _38465_ (.A1(\inst$top.soc.cpu.sink__payload$18[14] ),
    .A2(net2239),
    .B1(net2068),
    .Y(_16973_));
 sky130_fd_sc_hd__a21oi_1 _38466_ (.A1(_20789_),
    .A2(net2239),
    .B1(_16973_),
    .Y(_04686_));
 sky130_fd_sc_hd__o21ai_0 _38467_ (.A1(\inst$top.soc.cpu.sink__payload$18[15] ),
    .A2(net2241),
    .B1(net2071),
    .Y(_16974_));
 sky130_fd_sc_hd__a21oi_1 _38468_ (.A1(_20807_),
    .A2(net2241),
    .B1(_16974_),
    .Y(_04687_));
 sky130_fd_sc_hd__o21ai_0 _38470_ (.A1(\inst$top.soc.cpu.sink__payload$18[16] ),
    .A2(net2232),
    .B1(net2097),
    .Y(_16976_));
 sky130_fd_sc_hd__a21oi_1 _38471_ (.A1(_05598_),
    .A2(net2232),
    .B1(_16976_),
    .Y(_04688_));
 sky130_fd_sc_hd__inv_1 _38472_ (.A(\inst$top.soc.cpu.d.sink__payload.compare ),
    .Y(_16977_));
 sky130_fd_sc_hd__o21ai_0 _38473_ (.A1(net2829),
    .A2(net2277),
    .B1(net2178),
    .Y(_16978_));
 sky130_fd_sc_hd__a21oi_1 _38474_ (.A1(_16977_),
    .A2(net2284),
    .B1(_16978_),
    .Y(_04689_));
 sky130_fd_sc_hd__nor2_1 _38475_ (.A(\inst$top.soc.cpu.d.sink__payload.multiply ),
    .B(net1915),
    .Y(_16979_));
 sky130_fd_sc_hd__o21ai_0 _38476_ (.A1(\inst$top.soc.cpu.d.sink__payload$6.multiply ),
    .A2(net2279),
    .B1(net2147),
    .Y(_16980_));
 sky130_fd_sc_hd__nor2_1 _38477_ (.A(_16979_),
    .B(_16980_),
    .Y(_04690_));
 sky130_fd_sc_hd__o21ai_0 _38479_ (.A1(\inst$top.soc.cpu.d.sink__payload.divide ),
    .A2(net1913),
    .B1(net2149),
    .Y(_16982_));
 sky130_fd_sc_hd__a21oi_1 _38480_ (.A1(net2012),
    .A2(net1912),
    .B1(_16982_),
    .Y(_04691_));
 sky130_fd_sc_hd__o21ai_0 _38481_ (.A1(\inst$top.soc.cpu.d.sink__payload$6.condition_met ),
    .A2(net2276),
    .B1(net2146),
    .Y(_16983_));
 sky130_fd_sc_hd__nand2_1 _38482_ (.A(_14331_),
    .B(net1739),
    .Y(_16984_));
 sky130_fd_sc_hd__nand3_1 _38483_ (.A(_14328_),
    .B(net1480),
    .C(_14330_),
    .Y(_16985_));
 sky130_fd_sc_hd__nand4_1 _38484_ (.A(_16984_),
    .B(_16985_),
    .C(_09916_),
    .D(net2866),
    .Y(_16986_));
 sky130_fd_sc_hd__nand3_1 _38485_ (.A(_14340_),
    .B(net2005),
    .C(_02925_),
    .Y(_16987_));
 sky130_fd_sc_hd__nand3_1 _38486_ (.A(_14342_),
    .B(_16986_),
    .C(_16987_),
    .Y(_16988_));
 sky130_fd_sc_hd__inv_1 _38487_ (.A(_16986_),
    .Y(_16989_));
 sky130_fd_sc_hd__nand2_1 _38488_ (.A(_14857_),
    .B(_16989_),
    .Y(_16990_));
 sky130_fd_sc_hd__nand2_1 _38489_ (.A(_16988_),
    .B(_16990_),
    .Y(_16991_));
 sky130_fd_sc_hd__nor2_1 _38490_ (.A(\inst$top.soc.cpu.d.sink__payload.compare ),
    .B(_09447_),
    .Y(_16992_));
 sky130_fd_sc_hd__inv_1 _38491_ (.A(_16992_),
    .Y(_16993_));
 sky130_fd_sc_hd__o21ai_0 _38492_ (.A1(_09912_),
    .A2(_16977_),
    .B1(_16993_),
    .Y(_16994_));
 sky130_fd_sc_hd__nand2_1 _38493_ (.A(_16991_),
    .B(_16994_),
    .Y(_16995_));
 sky130_fd_sc_hd__nor3_1 _38494_ (.A(_09916_),
    .B(_02928_),
    .C(_14293_),
    .Y(_16996_));
 sky130_fd_sc_hd__nand2_1 _38495_ (.A(_16996_),
    .B(_14140_),
    .Y(_16997_));
 sky130_fd_sc_hd__nor4_1 _38496_ (.A(_13539_),
    .B(_13435_),
    .C(_13918_),
    .D(_16997_),
    .Y(_16998_));
 sky130_fd_sc_hd__nor3_1 _38497_ (.A(_03083_),
    .B(_13063_),
    .C(_13042_),
    .Y(_16999_));
 sky130_fd_sc_hd__nor4_1 _38498_ (.A(_13054_),
    .B(_13174_),
    .C(_13160_),
    .D(_13205_),
    .Y(_17000_));
 sky130_fd_sc_hd__nand3_1 _38499_ (.A(_16998_),
    .B(_16999_),
    .C(_17000_),
    .Y(_17001_));
 sky130_fd_sc_hd__o2111ai_1 _38500_ (.A1(\inst$top.soc.cpu.d.sink__payload.csr_fmt_i ),
    .A2(_17001_),
    .B1(_09912_),
    .C1(\inst$top.soc.cpu.sink__payload$12[143] ),
    .D1(_16977_),
    .Y(_17002_));
 sky130_fd_sc_hd__inv_1 _38501_ (.A(_17002_),
    .Y(_17003_));
 sky130_fd_sc_hd__nand2_1 _38502_ (.A(_16995_),
    .B(_17003_),
    .Y(_17004_));
 sky130_fd_sc_hd__nand3_1 _38503_ (.A(_13922_),
    .B(_14140_),
    .C(_16996_),
    .Y(_17005_));
 sky130_fd_sc_hd__nand2_1 _38504_ (.A(_14142_),
    .B(_16996_),
    .Y(_17006_));
 sky130_fd_sc_hd__nor3_1 _38505_ (.A(_09916_),
    .B(_02928_),
    .C(_14295_),
    .Y(_17007_));
 sky130_fd_sc_hd__a211oi_1 _38506_ (.A1(_02922_),
    .A2(_02930_),
    .B1(_02921_),
    .C1(_17007_),
    .Y(_17008_));
 sky130_fd_sc_hd__nand3_1 _38507_ (.A(_17005_),
    .B(_17006_),
    .C(_17008_),
    .Y(_17009_));
 sky130_fd_sc_hd__nand2_1 _38508_ (.A(_17009_),
    .B(net2867),
    .Y(_17010_));
 sky130_fd_sc_hd__a211oi_1 _38509_ (.A1(_09916_),
    .A2(_02678_),
    .B1(net2867),
    .C1(_02691_),
    .Y(_17011_));
 sky130_fd_sc_hd__nor3_1 _38510_ (.A(_02922_),
    .B(_14326_),
    .C(_14281_),
    .Y(_17012_));
 sky130_fd_sc_hd__nand2_1 _38511_ (.A(_14133_),
    .B(_17012_),
    .Y(_17013_));
 sky130_fd_sc_hd__o311ai_0 _38512_ (.A1(_02922_),
    .A2(_14326_),
    .A3(_14285_),
    .B1(_17011_),
    .C1(_17013_),
    .Y(_17014_));
 sky130_fd_sc_hd__nand2_1 _38513_ (.A(_17010_),
    .B(_17014_),
    .Y(_17015_));
 sky130_fd_sc_hd__nand2_1 _38514_ (.A(_16993_),
    .B(_16914_),
    .Y(_17016_));
 sky130_fd_sc_hd__nand2_1 _38515_ (.A(_16977_),
    .B(\inst$top.soc.cpu.sink__payload$12[143] ),
    .Y(_17017_));
 sky130_fd_sc_hd__nand3_1 _38516_ (.A(_17001_),
    .B(_16994_),
    .C(_17017_),
    .Y(_17018_));
 sky130_fd_sc_hd__a31oi_1 _38517_ (.A1(_17015_),
    .A2(\inst$top.soc.cpu.sink__payload$12[144] ),
    .A3(_17016_),
    .B1(_17018_),
    .Y(_17019_));
 sky130_fd_sc_hd__nand3_1 _38518_ (.A(_17016_),
    .B(\inst$top.soc.cpu.sink__payload$12[144] ),
    .C(_17017_),
    .Y(_17020_));
 sky130_fd_sc_hd__nand3_1 _38519_ (.A(_16988_),
    .B(_16990_),
    .C(_17020_),
    .Y(_17021_));
 sky130_fd_sc_hd__nand2_1 _38520_ (.A(_17019_),
    .B(_17021_),
    .Y(_17022_));
 sky130_fd_sc_hd__nor2_1 _38521_ (.A(_12969_),
    .B(_16993_),
    .Y(_17023_));
 sky130_fd_sc_hd__nor4_1 _38522_ (.A(\inst$top.soc.cpu.sink__payload$12[144] ),
    .B(\inst$top.soc.cpu.sink__payload$12[143] ),
    .C(_16992_),
    .D(_17001_),
    .Y(_17024_));
 sky130_fd_sc_hd__a21oi_1 _38523_ (.A1(_17015_),
    .A2(_17023_),
    .B1(_17024_),
    .Y(_17025_));
 sky130_fd_sc_hd__nand3_1 _38524_ (.A(_17004_),
    .B(_17022_),
    .C(_17025_),
    .Y(_17026_));
 sky130_fd_sc_hd__nor2_1 _38525_ (.A(net1912),
    .B(_17026_),
    .Y(_17027_));
 sky130_fd_sc_hd__nor2_1 _38526_ (.A(_16983_),
    .B(_17027_),
    .Y(_04692_));
 sky130_fd_sc_hd__o21ai_0 _38527_ (.A1(\inst$top.soc.cpu.sink__payload$18[17] ),
    .A2(net2232),
    .B1(net2097),
    .Y(_17028_));
 sky130_fd_sc_hd__a21oi_1 _38528_ (.A1(_05622_),
    .A2(net2234),
    .B1(_17028_),
    .Y(_04693_));
 sky130_fd_sc_hd__nand2_1 _38529_ (.A(net2851),
    .B(\inst$top.soc.cpu.d.sink__payload.rs1_re ),
    .Y(_17029_));
 sky130_fd_sc_hd__nand3_1 _38530_ (.A(net2226),
    .B(\inst$top.soc.cpu.sink__payload$12[109] ),
    .C(_17029_),
    .Y(_17030_));
 sky130_fd_sc_hd__nand2_1 _38531_ (.A(net1888),
    .B(\inst$top.soc.cpu.sink__payload$18[180] ),
    .Y(_17031_));
 sky130_fd_sc_hd__a21oi_1 _38532_ (.A1(_17030_),
    .A2(_17031_),
    .B1(net2939),
    .Y(_04694_));
 sky130_fd_sc_hd__a21oi_1 _38534_ (.A1(\inst$top.soc.cpu.sink__payload$12[110] ),
    .A2(_17029_),
    .B1(net1902),
    .Y(_17033_));
 sky130_fd_sc_hd__inv_1 _38535_ (.A(_17029_),
    .Y(_17034_));
 sky130_fd_sc_hd__nand2_1 _38537_ (.A(_13681_),
    .B(net1865),
    .Y(_17036_));
 sky130_fd_sc_hd__o21ai_0 _38538_ (.A1(\inst$top.soc.cpu.sink__payload$18[181] ),
    .A2(net2247),
    .B1(net2078),
    .Y(_17037_));
 sky130_fd_sc_hd__a21oi_1 _38539_ (.A1(_17033_),
    .A2(_17036_),
    .B1(_17037_),
    .Y(_04695_));
 sky130_fd_sc_hd__nand2_1 _38541_ (.A(net869),
    .B(net1863),
    .Y(_17039_));
 sky130_fd_sc_hd__a21oi_1 _38542_ (.A1(\inst$top.soc.cpu.sink__payload$12[162] ),
    .A2(_17029_),
    .B1(net1881),
    .Y(_17040_));
 sky130_fd_sc_hd__a221oi_1 _38543_ (.A1(_11843_),
    .A2(net1881),
    .B1(_17039_),
    .B2(_17040_),
    .C1(net2936),
    .Y(_04696_));
 sky130_fd_sc_hd__nand2_1 _38544_ (.A(net830),
    .B(net1863),
    .Y(_17041_));
 sky130_fd_sc_hd__a21oi_1 _38545_ (.A1(\inst$top.soc.cpu.sink__payload$12[163] ),
    .A2(_17029_),
    .B1(net1881),
    .Y(_17042_));
 sky130_fd_sc_hd__a221oi_1 _38546_ (.A1(_11858_),
    .A2(net1887),
    .B1(_17041_),
    .B2(_17042_),
    .C1(net2939),
    .Y(_04697_));
 sky130_fd_sc_hd__nand2_1 _38547_ (.A(net812),
    .B(net1863),
    .Y(_17043_));
 sky130_fd_sc_hd__a21oi_1 _38548_ (.A1(\inst$top.soc.cpu.sink__payload$12[164] ),
    .A2(_17029_),
    .B1(net1881),
    .Y(_17044_));
 sky130_fd_sc_hd__a221oi_1 _38549_ (.A1(_11865_),
    .A2(net1881),
    .B1(_17043_),
    .B2(_17044_),
    .C1(net2936),
    .Y(_04698_));
 sky130_fd_sc_hd__a21oi_1 _38550_ (.A1(_14434_),
    .A2(net1861),
    .B1(net1888),
    .Y(_17045_));
 sky130_fd_sc_hd__o21ai_0 _38551_ (.A1(\inst$top.soc.cpu.sink__payload$12[165] ),
    .A2(net1861),
    .B1(_17045_),
    .Y(_17046_));
 sky130_fd_sc_hd__nand2_1 _38552_ (.A(net1888),
    .B(\inst$top.soc.cpu.sink__payload$18[185] ),
    .Y(_17047_));
 sky130_fd_sc_hd__a21oi_1 _38553_ (.A1(_17046_),
    .A2(_17047_),
    .B1(net2939),
    .Y(_04699_));
 sky130_fd_sc_hd__a21oi_1 _38554_ (.A1(_14863_),
    .A2(net1861),
    .B1(net1888),
    .Y(_17048_));
 sky130_fd_sc_hd__o21ai_0 _38555_ (.A1(\inst$top.soc.cpu.sink__payload$12[166] ),
    .A2(net1861),
    .B1(_17048_),
    .Y(_17049_));
 sky130_fd_sc_hd__nand2_1 _38556_ (.A(net1887),
    .B(\inst$top.soc.cpu.sink__payload$18[186] ),
    .Y(_17050_));
 sky130_fd_sc_hd__a21oi_1 _38557_ (.A1(_17049_),
    .A2(_17050_),
    .B1(net2939),
    .Y(_04700_));
 sky130_fd_sc_hd__a21oi_1 _38558_ (.A1(_14866_),
    .A2(net1863),
    .B1(net1881),
    .Y(_17051_));
 sky130_fd_sc_hd__o21ai_0 _38559_ (.A1(\inst$top.soc.cpu.sink__payload$12[167] ),
    .A2(net1863),
    .B1(_17051_),
    .Y(_17052_));
 sky130_fd_sc_hd__nand2_1 _38560_ (.A(net1882),
    .B(\inst$top.soc.cpu.sink__payload$18[187] ),
    .Y(_17053_));
 sky130_fd_sc_hd__a21oi_1 _38561_ (.A1(_17052_),
    .A2(_17053_),
    .B1(net2938),
    .Y(_04701_));
 sky130_fd_sc_hd__a21oi_1 _38562_ (.A1(net734),
    .A2(net1864),
    .B1(net1896),
    .Y(_17054_));
 sky130_fd_sc_hd__o21ai_0 _38563_ (.A1(\inst$top.soc.cpu.sink__payload$12[168] ),
    .A2(net1864),
    .B1(_17054_),
    .Y(_17055_));
 sky130_fd_sc_hd__nand2_1 _38564_ (.A(net1896),
    .B(\inst$top.soc.cpu.sink__payload$18[188] ),
    .Y(_17056_));
 sky130_fd_sc_hd__a21oi_1 _38566_ (.A1(_17055_),
    .A2(_17056_),
    .B1(net2952),
    .Y(_04702_));
 sky130_fd_sc_hd__a21oi_1 _38567_ (.A1(net662),
    .A2(net1862),
    .B1(net1889),
    .Y(_17058_));
 sky130_fd_sc_hd__o21ai_0 _38568_ (.A1(\inst$top.soc.cpu.sink__payload$12[169] ),
    .A2(net1862),
    .B1(_17058_),
    .Y(_17059_));
 sky130_fd_sc_hd__nand2_1 _38569_ (.A(net1889),
    .B(\inst$top.soc.cpu.sink__payload$18[189] ),
    .Y(_17060_));
 sky130_fd_sc_hd__a21oi_1 _38570_ (.A1(_17059_),
    .A2(_17060_),
    .B1(net2941),
    .Y(_04703_));
 sky130_fd_sc_hd__o21ai_0 _38572_ (.A1(\inst$top.soc.cpu.sink__payload$18[18] ),
    .A2(net2233),
    .B1(net2093),
    .Y(_17062_));
 sky130_fd_sc_hd__a21oi_1 _38573_ (.A1(_05644_),
    .A2(net2233),
    .B1(_17062_),
    .Y(_04704_));
 sky130_fd_sc_hd__a21oi_1 _38575_ (.A1(_14870_),
    .A2(net1864),
    .B1(net1896),
    .Y(_17064_));
 sky130_fd_sc_hd__o21ai_0 _38576_ (.A1(\inst$top.soc.cpu.sink__payload$12[170] ),
    .A2(net1864),
    .B1(_17064_),
    .Y(_17065_));
 sky130_fd_sc_hd__nand2_1 _38577_ (.A(net1894),
    .B(\inst$top.soc.cpu.sink__payload$18[190] ),
    .Y(_17066_));
 sky130_fd_sc_hd__a21oi_1 _38578_ (.A1(_17065_),
    .A2(_17066_),
    .B1(net2953),
    .Y(_04705_));
 sky130_fd_sc_hd__nand2_1 _38581_ (.A(_14872_),
    .B(net1861),
    .Y(_17069_));
 sky130_fd_sc_hd__o211ai_1 _38582_ (.A1(\inst$top.soc.cpu.sink__payload$12[171] ),
    .A2(net1861),
    .B1(net2237),
    .C1(_17069_),
    .Y(_17070_));
 sky130_fd_sc_hd__nand2_1 _38584_ (.A(net1887),
    .B(\inst$top.soc.cpu.sink__payload$18[191] ),
    .Y(_17072_));
 sky130_fd_sc_hd__a21oi_1 _38585_ (.A1(_17070_),
    .A2(_17072_),
    .B1(net2939),
    .Y(_04706_));
 sky130_fd_sc_hd__nand2_1 _38586_ (.A(_13217_),
    .B(net1862),
    .Y(_17073_));
 sky130_fd_sc_hd__o211ai_1 _38587_ (.A1(\inst$top.soc.cpu.sink__payload$12[172] ),
    .A2(net1862),
    .B1(net2237),
    .C1(_17073_),
    .Y(_17074_));
 sky130_fd_sc_hd__nand2_1 _38588_ (.A(net1889),
    .B(\inst$top.soc.cpu.sink__payload$18[192] ),
    .Y(_17075_));
 sky130_fd_sc_hd__a21oi_1 _38589_ (.A1(_17074_),
    .A2(_17075_),
    .B1(net2941),
    .Y(_04707_));
 sky130_fd_sc_hd__a21oi_1 _38590_ (.A1(_14823_),
    .A2(net1864),
    .B1(net1896),
    .Y(_17076_));
 sky130_fd_sc_hd__o21ai_0 _38591_ (.A1(\inst$top.soc.cpu.sink__payload$12[173] ),
    .A2(net1864),
    .B1(_17076_),
    .Y(_17077_));
 sky130_fd_sc_hd__nand2_1 _38592_ (.A(net1896),
    .B(\inst$top.soc.cpu.sink__payload$18[193] ),
    .Y(_17078_));
 sky130_fd_sc_hd__a21oi_1 _38593_ (.A1(_17077_),
    .A2(_17078_),
    .B1(net2952),
    .Y(_04708_));
 sky130_fd_sc_hd__a21oi_1 _38594_ (.A1(_13327_),
    .A2(net1864),
    .B1(net1896),
    .Y(_17079_));
 sky130_fd_sc_hd__o21ai_0 _38595_ (.A1(\inst$top.soc.cpu.sink__payload$12[174] ),
    .A2(net1864),
    .B1(_17079_),
    .Y(_17080_));
 sky130_fd_sc_hd__nand2_1 _38596_ (.A(net1896),
    .B(\inst$top.soc.cpu.sink__payload$18[194] ),
    .Y(_17081_));
 sky130_fd_sc_hd__a21oi_1 _38597_ (.A1(_17080_),
    .A2(_17081_),
    .B1(net2952),
    .Y(_04709_));
 sky130_fd_sc_hd__nand2_1 _38598_ (.A(_14826_),
    .B(net1865),
    .Y(_17082_));
 sky130_fd_sc_hd__o211ai_1 _38599_ (.A1(\inst$top.soc.cpu.sink__payload$12[175] ),
    .A2(net1865),
    .B1(net2241),
    .C1(_17082_),
    .Y(_17083_));
 sky130_fd_sc_hd__nand2_1 _38600_ (.A(net1894),
    .B(\inst$top.soc.cpu.sink__payload$18[195] ),
    .Y(_17084_));
 sky130_fd_sc_hd__a21oi_1 _38601_ (.A1(_17083_),
    .A2(_17084_),
    .B1(net2953),
    .Y(_04710_));
 sky130_fd_sc_hd__a21oi_1 _38602_ (.A1(_13448_),
    .A2(net1862),
    .B1(net1889),
    .Y(_17085_));
 sky130_fd_sc_hd__o21ai_0 _38603_ (.A1(\inst$top.soc.cpu.sink__payload$12[176] ),
    .A2(net1862),
    .B1(_17085_),
    .Y(_17086_));
 sky130_fd_sc_hd__nand2_1 _38604_ (.A(net1890),
    .B(\inst$top.soc.cpu.sink__payload$18[196] ),
    .Y(_17087_));
 sky130_fd_sc_hd__a21oi_1 _38605_ (.A1(_17086_),
    .A2(_17087_),
    .B1(net2941),
    .Y(_04711_));
 sky130_fd_sc_hd__a21oi_1 _38606_ (.A1(_13515_),
    .A2(net1864),
    .B1(net1889),
    .Y(_17088_));
 sky130_fd_sc_hd__o21ai_0 _38607_ (.A1(\inst$top.soc.cpu.sink__payload$12[177] ),
    .A2(net1864),
    .B1(_17088_),
    .Y(_17089_));
 sky130_fd_sc_hd__nand2_1 _38608_ (.A(net1890),
    .B(\inst$top.soc.cpu.sink__payload$18[197] ),
    .Y(_17090_));
 sky130_fd_sc_hd__a21oi_1 _38609_ (.A1(_17089_),
    .A2(_17090_),
    .B1(net2941),
    .Y(_04712_));
 sky130_fd_sc_hd__nand2_1 _38611_ (.A(_13564_),
    .B(net1861),
    .Y(_17092_));
 sky130_fd_sc_hd__o211ai_1 _38612_ (.A1(\inst$top.soc.cpu.sink__payload$12[178] ),
    .A2(net1861),
    .B1(net2237),
    .C1(_17092_),
    .Y(_17093_));
 sky130_fd_sc_hd__nand2_1 _38613_ (.A(net1888),
    .B(\inst$top.soc.cpu.sink__payload$18[198] ),
    .Y(_17094_));
 sky130_fd_sc_hd__a21oi_1 _38615_ (.A1(_17093_),
    .A2(_17094_),
    .B1(net2941),
    .Y(_04713_));
 sky130_fd_sc_hd__nand2_1 _38617_ (.A(_13653_),
    .B(net1862),
    .Y(_17097_));
 sky130_fd_sc_hd__o211ai_1 _38618_ (.A1(\inst$top.soc.cpu.sink__payload$12[179] ),
    .A2(net1862),
    .B1(net2237),
    .C1(_17097_),
    .Y(_17098_));
 sky130_fd_sc_hd__nand2_1 _38619_ (.A(net1889),
    .B(\inst$top.soc.cpu.sink__payload$18[199] ),
    .Y(_17099_));
 sky130_fd_sc_hd__a21oi_1 _38620_ (.A1(_17098_),
    .A2(_17099_),
    .B1(net2943),
    .Y(_04714_));
 sky130_fd_sc_hd__o21ai_0 _38621_ (.A1(\inst$top.soc.cpu.sink__payload$18[19] ),
    .A2(net2232),
    .B1(net2097),
    .Y(_17100_));
 sky130_fd_sc_hd__a21oi_1 _38622_ (.A1(_05666_),
    .A2(net2232),
    .B1(_17100_),
    .Y(_04715_));
 sky130_fd_sc_hd__nand2_1 _38623_ (.A(_13729_),
    .B(net1861),
    .Y(_17101_));
 sky130_fd_sc_hd__o211ai_1 _38624_ (.A1(\inst$top.soc.cpu.sink__payload$12[180] ),
    .A2(net1861),
    .B1(net2237),
    .C1(_17101_),
    .Y(_17102_));
 sky130_fd_sc_hd__nand2_1 _38625_ (.A(net1888),
    .B(\inst$top.soc.cpu.sink__payload$18[200] ),
    .Y(_17103_));
 sky130_fd_sc_hd__a21oi_1 _38626_ (.A1(_17102_),
    .A2(_17103_),
    .B1(net2939),
    .Y(_04716_));
 sky130_fd_sc_hd__nand2_1 _38627_ (.A(_13780_),
    .B(net1862),
    .Y(_17104_));
 sky130_fd_sc_hd__o211ai_1 _38628_ (.A1(\inst$top.soc.cpu.sink__payload$12[181] ),
    .A2(net1862),
    .B1(net2237),
    .C1(_17104_),
    .Y(_17105_));
 sky130_fd_sc_hd__nand2_1 _38630_ (.A(net1889),
    .B(\inst$top.soc.cpu.sink__payload$18[201] ),
    .Y(_17107_));
 sky130_fd_sc_hd__a21oi_1 _38631_ (.A1(_17105_),
    .A2(_17107_),
    .B1(net2941),
    .Y(_04717_));
 sky130_fd_sc_hd__nand2_1 _38632_ (.A(_14838_),
    .B(net1867),
    .Y(_17108_));
 sky130_fd_sc_hd__o211ai_1 _38633_ (.A1(\inst$top.soc.cpu.sink__payload$12[182] ),
    .A2(net1867),
    .B1(net2238),
    .C1(_17108_),
    .Y(_17109_));
 sky130_fd_sc_hd__nand2_1 _38634_ (.A(net1896),
    .B(\inst$top.soc.cpu.sink__payload$18[202] ),
    .Y(_17110_));
 sky130_fd_sc_hd__a21oi_1 _38635_ (.A1(_17109_),
    .A2(_17110_),
    .B1(net2952),
    .Y(_04718_));
 sky130_fd_sc_hd__nand2_1 _38636_ (.A(_14841_),
    .B(net1865),
    .Y(_17111_));
 sky130_fd_sc_hd__o211ai_1 _38637_ (.A1(\inst$top.soc.cpu.sink__payload$12[183] ),
    .A2(net1865),
    .B1(net2238),
    .C1(_17111_),
    .Y(_17112_));
 sky130_fd_sc_hd__nand2_1 _38638_ (.A(net1894),
    .B(\inst$top.soc.cpu.sink__payload$18[203] ),
    .Y(_17113_));
 sky130_fd_sc_hd__a21oi_1 _38639_ (.A1(_17112_),
    .A2(_17113_),
    .B1(net2954),
    .Y(_04719_));
 sky130_fd_sc_hd__nand2_1 _38640_ (.A(_14843_),
    .B(net1865),
    .Y(_17114_));
 sky130_fd_sc_hd__o211ai_1 _38641_ (.A1(\inst$top.soc.cpu.sink__payload$12[184] ),
    .A2(net1865),
    .B1(net2238),
    .C1(_17114_),
    .Y(_17115_));
 sky130_fd_sc_hd__nand2_1 _38642_ (.A(net1894),
    .B(\inst$top.soc.cpu.sink__payload$18[204] ),
    .Y(_17116_));
 sky130_fd_sc_hd__a21oi_1 _38643_ (.A1(_17115_),
    .A2(_17116_),
    .B1(net2954),
    .Y(_04720_));
 sky130_fd_sc_hd__a21oi_1 _38644_ (.A1(_13990_),
    .A2(net1863),
    .B1(net1881),
    .Y(_17117_));
 sky130_fd_sc_hd__o21ai_0 _38645_ (.A1(\inst$top.soc.cpu.sink__payload$12[185] ),
    .A2(net1863),
    .B1(_17117_),
    .Y(_17118_));
 sky130_fd_sc_hd__nand2_1 _38646_ (.A(net1882),
    .B(\inst$top.soc.cpu.sink__payload$18[205] ),
    .Y(_17119_));
 sky130_fd_sc_hd__a21oi_1 _38647_ (.A1(_17118_),
    .A2(_17119_),
    .B1(net2938),
    .Y(_04721_));
 sky130_fd_sc_hd__nand2_1 _38648_ (.A(_14046_),
    .B(net1866),
    .Y(_17120_));
 sky130_fd_sc_hd__o211ai_1 _38649_ (.A1(\inst$top.soc.cpu.sink__payload$12[186] ),
    .A2(net1866),
    .B1(net2250),
    .C1(_17120_),
    .Y(_17121_));
 sky130_fd_sc_hd__nand2_1 _38650_ (.A(net1894),
    .B(\inst$top.soc.cpu.sink__payload$18[206] ),
    .Y(_17122_));
 sky130_fd_sc_hd__a21oi_1 _38651_ (.A1(_17121_),
    .A2(_17122_),
    .B1(net2954),
    .Y(_04722_));
 sky130_fd_sc_hd__nor2_1 _38652_ (.A(\inst$top.soc.cpu.sink__payload$12[187] ),
    .B(net1865),
    .Y(_17123_));
 sky130_fd_sc_hd__nor2_1 _38653_ (.A(_17123_),
    .B(net1904),
    .Y(_17124_));
 sky130_fd_sc_hd__o21ai_0 _38654_ (.A1(_17029_),
    .A2(_14848_),
    .B1(_17124_),
    .Y(_17125_));
 sky130_fd_sc_hd__nand2_1 _38655_ (.A(net1901),
    .B(\inst$top.soc.cpu.sink__payload$18[207] ),
    .Y(_17126_));
 sky130_fd_sc_hd__a21oi_1 _38656_ (.A1(_17125_),
    .A2(_17126_),
    .B1(net2955),
    .Y(_04723_));
 sky130_fd_sc_hd__nand2_1 _38657_ (.A(_14850_),
    .B(net1866),
    .Y(_17127_));
 sky130_fd_sc_hd__o211ai_1 _38658_ (.A1(\inst$top.soc.cpu.sink__payload$12[188] ),
    .A2(net1866),
    .B1(net2250),
    .C1(_17127_),
    .Y(_17128_));
 sky130_fd_sc_hd__nand2_1 _38659_ (.A(net1901),
    .B(\inst$top.soc.cpu.sink__payload$18[208] ),
    .Y(_17129_));
 sky130_fd_sc_hd__a21oi_1 _38661_ (.A1(_17128_),
    .A2(_17129_),
    .B1(net2954),
    .Y(_04724_));
 sky130_fd_sc_hd__nand2_1 _38662_ (.A(_14853_),
    .B(net1866),
    .Y(_17131_));
 sky130_fd_sc_hd__o211ai_1 _38663_ (.A1(\inst$top.soc.cpu.sink__payload$12[189] ),
    .A2(net1865),
    .B1(net2238),
    .C1(_17131_),
    .Y(_17132_));
 sky130_fd_sc_hd__nand2_1 _38664_ (.A(net1894),
    .B(\inst$top.soc.cpu.sink__payload$18[209] ),
    .Y(_17133_));
 sky130_fd_sc_hd__a21oi_1 _38665_ (.A1(_17132_),
    .A2(_17133_),
    .B1(net2954),
    .Y(_04725_));
 sky130_fd_sc_hd__o21ai_0 _38666_ (.A1(\inst$top.soc.cpu.sink__payload$18[20] ),
    .A2(net2231),
    .B1(net2094),
    .Y(_17134_));
 sky130_fd_sc_hd__a21oi_1 _38667_ (.A1(_12244_),
    .A2(net2231),
    .B1(_17134_),
    .Y(_04726_));
 sky130_fd_sc_hd__nand2_1 _38668_ (.A(_14855_),
    .B(net1865),
    .Y(_17135_));
 sky130_fd_sc_hd__o211ai_1 _38669_ (.A1(\inst$top.soc.cpu.sink__payload$12[190] ),
    .A2(net1866),
    .B1(net2238),
    .C1(_17135_),
    .Y(_17136_));
 sky130_fd_sc_hd__nand2_1 _38670_ (.A(net1894),
    .B(\inst$top.soc.cpu.sink__payload$18[210] ),
    .Y(_17137_));
 sky130_fd_sc_hd__a21oi_1 _38671_ (.A1(_17136_),
    .A2(_17137_),
    .B1(net2954),
    .Y(_04727_));
 sky130_fd_sc_hd__nand2_1 _38672_ (.A(_14857_),
    .B(net1863),
    .Y(_17138_));
 sky130_fd_sc_hd__o211ai_1 _38673_ (.A1(\inst$top.soc.cpu.sink__payload$12[191] ),
    .A2(net1863),
    .B1(net2237),
    .C1(_17138_),
    .Y(_17139_));
 sky130_fd_sc_hd__nand2_1 _38674_ (.A(net1882),
    .B(\inst$top.soc.cpu.sink__payload$18[211] ),
    .Y(_17140_));
 sky130_fd_sc_hd__a21oi_1 _38675_ (.A1(_17139_),
    .A2(_17140_),
    .B1(net2938),
    .Y(_04728_));
 sky130_fd_sc_hd__nand2_1 _38676_ (.A(_17026_),
    .B(\inst$top.soc.cpu.d.sink__payload.branch ),
    .Y(_17141_));
 sky130_fd_sc_hd__nor2_1 _38677_ (.A(net2852),
    .B(net1903),
    .Y(_17142_));
 sky130_fd_sc_hd__o21ai_0 _38678_ (.A1(\inst$top.soc.cpu.d.sink__payload$6.branch_taken ),
    .A2(net2247),
    .B1(net2080),
    .Y(_17143_));
 sky130_fd_sc_hd__a21oi_1 _38679_ (.A1(_17141_),
    .A2(_17142_),
    .B1(_17143_),
    .Y(_04729_));
 sky130_fd_sc_hd__o21ai_0 _38680_ (.A1(\inst$top.soc.cpu.d.sink__payload.branch_predict_taken ),
    .A2(net1887),
    .B1(net2042),
    .Y(_17144_));
 sky130_fd_sc_hd__a21oi_1 _38681_ (.A1(_02864_),
    .A2(net1887),
    .B1(_17144_),
    .Y(_04730_));
 sky130_fd_sc_hd__nor2_1 _38682_ (.A(\inst$top.soc.cpu.d.sink__payload.csr_we ),
    .B(net1895),
    .Y(_17145_));
 sky130_fd_sc_hd__o21ai_0 _38683_ (.A1(\inst$top.soc.cpu.d.sink__payload$6.csr_we ),
    .A2(net2238),
    .B1(net2066),
    .Y(_17146_));
 sky130_fd_sc_hd__nor2_1 _38684_ (.A(_17145_),
    .B(_17146_),
    .Y(_04731_));
 sky130_fd_sc_hd__nor2_1 _38685_ (.A(\inst$top.soc.cpu.d.sink__payload.csr_clear ),
    .B(\inst$top.soc.cpu.d.sink__payload.csr_set ),
    .Y(_17147_));
 sky130_fd_sc_hd__inv_1 _38686_ (.A(net1994),
    .Y(_17148_));
 sky130_fd_sc_hd__nand2_1 _38687_ (.A(_12979_),
    .B(net1859),
    .Y(_17149_));
 sky130_fd_sc_hd__nand2_1 _38689_ (.A(_03082_),
    .B(net1995),
    .Y(_17151_));
 sky130_fd_sc_hd__o21ai_0 _38690_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[0] ),
    .A2(net2263),
    .B1(net2111),
    .Y(_17152_));
 sky130_fd_sc_hd__a31oi_1 _38691_ (.A1(_17149_),
    .A2(_17151_),
    .A3(net2263),
    .B1(_17152_),
    .Y(_04732_));
 sky130_fd_sc_hd__or2_2 _38692_ (.A(net1995),
    .B(_13679_),
    .X(_17153_));
 sky130_fd_sc_hd__nand2_1 _38693_ (.A(net1262),
    .B(net1995),
    .Y(_17154_));
 sky130_fd_sc_hd__o21ai_0 _38694_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[1] ),
    .A2(net2263),
    .B1(net2111),
    .Y(_17155_));
 sky130_fd_sc_hd__a31oi_1 _38695_ (.A1(_17153_),
    .A2(net2263),
    .A3(_17154_),
    .B1(_17155_),
    .Y(_04733_));
 sky130_fd_sc_hd__nand2_1 _38697_ (.A(_14258_),
    .B(net1858),
    .Y(_17157_));
 sky130_fd_sc_hd__o211ai_1 _38698_ (.A1(net1366),
    .A2(net1858),
    .B1(net2247),
    .C1(_17157_),
    .Y(_17158_));
 sky130_fd_sc_hd__o211ai_1 _38699_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[2] ),
    .A2(net2217),
    .B1(net2034),
    .C1(net3036),
    .Y(_17159_));
 sky130_fd_sc_hd__inv_2 _38700_ (.A(_17159_),
    .Y(_04734_));
 sky130_fd_sc_hd__a21oi_1 _38702_ (.A1(net1361),
    .A2(net1993),
    .B1(net1906),
    .Y(_17161_));
 sky130_fd_sc_hd__o21ai_2 _38703_ (.A1(net1993),
    .A2(_14374_),
    .B1(_17161_),
    .Y(_17162_));
 sky130_fd_sc_hd__o211ai_1 _38704_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[3] ),
    .A2(net2225),
    .B1(net2088),
    .C1(_17162_),
    .Y(_17163_));
 sky130_fd_sc_hd__inv_2 _38705_ (.A(_17163_),
    .Y(_04735_));
 sky130_fd_sc_hd__nand2_1 _38706_ (.A(_14408_),
    .B(net1858),
    .Y(_17164_));
 sky130_fd_sc_hd__o211ai_1 _38707_ (.A1(net1858),
    .A2(_05894_),
    .B1(net2247),
    .C1(_17164_),
    .Y(_17165_));
 sky130_fd_sc_hd__o211ai_1 _38708_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[4] ),
    .A2(net2240),
    .B1(net2070),
    .C1(_17165_),
    .Y(_17166_));
 sky130_fd_sc_hd__inv_2 _38709_ (.A(_17166_),
    .Y(_04736_));
 sky130_fd_sc_hd__nor2_1 _38710_ (.A(\inst$top.soc.cpu.sink__payload$12[21] ),
    .B(net1891),
    .Y(_17167_));
 sky130_fd_sc_hd__o21ai_0 _38711_ (.A1(\inst$top.soc.cpu.sink__payload$18[21] ),
    .A2(net2230),
    .B1(net2093),
    .Y(_17168_));
 sky130_fd_sc_hd__nor2_1 _38712_ (.A(_17167_),
    .B(_17168_),
    .Y(_04737_));
 sky130_fd_sc_hd__nand2_1 _38714_ (.A(_14439_),
    .B(net1858),
    .Y(_17170_));
 sky130_fd_sc_hd__a21oi_1 _38716_ (.A1(net1351),
    .A2(net1993),
    .B1(net1903),
    .Y(_17172_));
 sky130_fd_sc_hd__o21ai_0 _38717_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[5] ),
    .A2(net2247),
    .B1(net2080),
    .Y(_17173_));
 sky130_fd_sc_hd__a21oi_1 _38718_ (.A1(_17170_),
    .A2(_17172_),
    .B1(_17173_),
    .Y(_04738_));
 sky130_fd_sc_hd__nand2_1 _38719_ (.A(_14461_),
    .B(net1858),
    .Y(_17174_));
 sky130_fd_sc_hd__a21oi_1 _38721_ (.A1(net1350),
    .A2(net1996),
    .B1(net1906),
    .Y(_17176_));
 sky130_fd_sc_hd__o21ai_0 _38722_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[6] ),
    .A2(net2248),
    .B1(net2112),
    .Y(_17177_));
 sky130_fd_sc_hd__a21oi_1 _38723_ (.A1(_17174_),
    .A2(_17176_),
    .B1(_17177_),
    .Y(_04739_));
 sky130_fd_sc_hd__o21ai_0 _38724_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[7] ),
    .A2(net2242),
    .B1(net2105),
    .Y(_17178_));
 sky130_fd_sc_hd__a21oi_1 _38725_ (.A1(net1345),
    .A2(net1994),
    .B1(net1898),
    .Y(_17179_));
 sky130_fd_sc_hd__o21a_1 _38726_ (.A1(net1994),
    .A2(_14489_),
    .B1(_17179_),
    .X(_17180_));
 sky130_fd_sc_hd__nor2_1 _38727_ (.A(_17178_),
    .B(_17180_),
    .Y(_04740_));
 sky130_fd_sc_hd__nand2_1 _38728_ (.A(_14524_),
    .B(net1858),
    .Y(_17181_));
 sky130_fd_sc_hd__a21oi_1 _38729_ (.A1(net1341),
    .A2(net1996),
    .B1(net1903),
    .Y(_17182_));
 sky130_fd_sc_hd__o21ai_0 _38731_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[8] ),
    .A2(net2247),
    .B1(net2081),
    .Y(_17184_));
 sky130_fd_sc_hd__a21oi_1 _38732_ (.A1(_17181_),
    .A2(_17182_),
    .B1(_17184_),
    .Y(_04741_));
 sky130_fd_sc_hd__nand2_1 _38733_ (.A(_14555_),
    .B(net1857),
    .Y(_17185_));
 sky130_fd_sc_hd__a21oi_1 _38734_ (.A1(net1336),
    .A2(net1993),
    .B1(net1901),
    .Y(_17186_));
 sky130_fd_sc_hd__o21ai_0 _38735_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[9] ),
    .A2(net2247),
    .B1(net2079),
    .Y(_17187_));
 sky130_fd_sc_hd__a21oi_1 _38736_ (.A1(_17185_),
    .A2(_17186_),
    .B1(_17187_),
    .Y(_04742_));
 sky130_fd_sc_hd__nand2_1 _38737_ (.A(_13091_),
    .B(net1858),
    .Y(_17188_));
 sky130_fd_sc_hd__a21oi_1 _38738_ (.A1(net1331),
    .A2(net1996),
    .B1(net1906),
    .Y(_17189_));
 sky130_fd_sc_hd__o21ai_0 _38739_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[10] ),
    .A2(net2248),
    .B1(net2112),
    .Y(_17190_));
 sky130_fd_sc_hd__a21oi_1 _38740_ (.A1(_17188_),
    .A2(_17189_),
    .B1(_17190_),
    .Y(_04743_));
 sky130_fd_sc_hd__nand2_1 _38741_ (.A(_13128_),
    .B(net1858),
    .Y(_17191_));
 sky130_fd_sc_hd__a21oi_1 _38742_ (.A1(net1327),
    .A2(net1993),
    .B1(net1906),
    .Y(_17192_));
 sky130_fd_sc_hd__o21ai_0 _38743_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[11] ),
    .A2(net2247),
    .B1(net2112),
    .Y(_17193_));
 sky130_fd_sc_hd__a21oi_1 _38744_ (.A1(_17191_),
    .A2(_17192_),
    .B1(_17193_),
    .Y(_04744_));
 sky130_fd_sc_hd__nand2_1 _38745_ (.A(_13222_),
    .B(net1857),
    .Y(_17194_));
 sky130_fd_sc_hd__a21oi_1 _38746_ (.A1(net1322),
    .A2(net1993),
    .B1(net1897),
    .Y(_17195_));
 sky130_fd_sc_hd__o21ai_0 _38748_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[12] ),
    .A2(net2243),
    .B1(net2070),
    .Y(_17197_));
 sky130_fd_sc_hd__a21oi_1 _38749_ (.A1(_17194_),
    .A2(_17195_),
    .B1(_17197_),
    .Y(_04745_));
 sky130_fd_sc_hd__nand2_1 _38750_ (.A(_13284_),
    .B(net1859),
    .Y(_17198_));
 sky130_fd_sc_hd__a21oi_1 _38751_ (.A1(net1317),
    .A2(net1993),
    .B1(net1905),
    .Y(_17199_));
 sky130_fd_sc_hd__o21ai_0 _38752_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[13] ),
    .A2(net2248),
    .B1(net2111),
    .Y(_17200_));
 sky130_fd_sc_hd__a21oi_1 _38753_ (.A1(_17198_),
    .A2(_17199_),
    .B1(_17200_),
    .Y(_04746_));
 sky130_fd_sc_hd__nand2_1 _38754_ (.A(_13332_),
    .B(net1857),
    .Y(_17201_));
 sky130_fd_sc_hd__a21oi_1 _38755_ (.A1(net1312),
    .A2(net1993),
    .B1(net1897),
    .Y(_17202_));
 sky130_fd_sc_hd__o21ai_0 _38756_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[14] ),
    .A2(net2241),
    .B1(net2071),
    .Y(_17203_));
 sky130_fd_sc_hd__a21oi_1 _38757_ (.A1(_17201_),
    .A2(_17202_),
    .B1(_17203_),
    .Y(_04747_));
 sky130_fd_sc_hd__o21ai_0 _38758_ (.A1(\inst$top.soc.cpu.sink__payload$18[22] ),
    .A2(net2246),
    .B1(net2104),
    .Y(_17204_));
 sky130_fd_sc_hd__a21oi_1 _38759_ (.A1(_12304_),
    .A2(net2246),
    .B1(_17204_),
    .Y(_04748_));
 sky130_fd_sc_hd__nand2_1 _38760_ (.A(_13379_),
    .B(net1857),
    .Y(_17205_));
 sky130_fd_sc_hd__a21oi_1 _38762_ (.A1(net1308),
    .A2(net1993),
    .B1(net1895),
    .Y(_17207_));
 sky130_fd_sc_hd__o21ai_0 _38763_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[15] ),
    .A2(net2241),
    .B1(net2070),
    .Y(_17208_));
 sky130_fd_sc_hd__a21oi_1 _38764_ (.A1(_17205_),
    .A2(_17207_),
    .B1(_17208_),
    .Y(_04749_));
 sky130_fd_sc_hd__nand2_1 _38766_ (.A(_13452_),
    .B(net1860),
    .Y(_17210_));
 sky130_fd_sc_hd__a21oi_1 _38767_ (.A1(net1303),
    .A2(net1994),
    .B1(net1905),
    .Y(_17211_));
 sky130_fd_sc_hd__o21ai_0 _38768_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[16] ),
    .A2(net2263),
    .B1(net2111),
    .Y(_17212_));
 sky130_fd_sc_hd__a21oi_1 _38769_ (.A1(_17210_),
    .A2(_17211_),
    .B1(_17212_),
    .Y(_04750_));
 sky130_fd_sc_hd__nand2_1 _38770_ (.A(_13519_),
    .B(net1860),
    .Y(_17213_));
 sky130_fd_sc_hd__a21oi_1 _38771_ (.A1(net1299),
    .A2(net1994),
    .B1(net1905),
    .Y(_17214_));
 sky130_fd_sc_hd__o21ai_0 _38773_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[17] ),
    .A2(net2263),
    .B1(net2111),
    .Y(_17216_));
 sky130_fd_sc_hd__a21oi_1 _38774_ (.A1(_17213_),
    .A2(_17214_),
    .B1(_17216_),
    .Y(_04751_));
 sky130_fd_sc_hd__nand2_1 _38775_ (.A(_13569_),
    .B(net1859),
    .Y(_17217_));
 sky130_fd_sc_hd__a21oi_1 _38776_ (.A1(net1295),
    .A2(net1995),
    .B1(net1908),
    .Y(_17218_));
 sky130_fd_sc_hd__o21ai_0 _38777_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[18] ),
    .A2(net2263),
    .B1(net2113),
    .Y(_17219_));
 sky130_fd_sc_hd__a21oi_1 _38778_ (.A1(_17217_),
    .A2(_17218_),
    .B1(_17219_),
    .Y(_04752_));
 sky130_fd_sc_hd__nand2_1 _38779_ (.A(_13657_),
    .B(net1860),
    .Y(_17220_));
 sky130_fd_sc_hd__a21oi_1 _38780_ (.A1(net1289),
    .A2(net1995),
    .B1(net1908),
    .Y(_17221_));
 sky130_fd_sc_hd__o21ai_0 _38781_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[19] ),
    .A2(net2261),
    .B1(net2109),
    .Y(_17222_));
 sky130_fd_sc_hd__a21oi_1 _38782_ (.A1(_17220_),
    .A2(_17221_),
    .B1(_17222_),
    .Y(_04753_));
 sky130_fd_sc_hd__nand2_1 _38783_ (.A(_13699_),
    .B(net1857),
    .Y(_17223_));
 sky130_fd_sc_hd__a21oi_1 _38784_ (.A1(net1286),
    .A2(net1994),
    .B1(net1907),
    .Y(_17224_));
 sky130_fd_sc_hd__o21ai_0 _38785_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[20] ),
    .A2(net2261),
    .B1(net2109),
    .Y(_17225_));
 sky130_fd_sc_hd__a21oi_1 _38786_ (.A1(_17223_),
    .A2(_17224_),
    .B1(_17225_),
    .Y(_04754_));
 sky130_fd_sc_hd__nand2_1 _38787_ (.A(_13785_),
    .B(net1858),
    .Y(_17226_));
 sky130_fd_sc_hd__a21oi_1 _38788_ (.A1(net1281),
    .A2(net1993),
    .B1(net1906),
    .Y(_17227_));
 sky130_fd_sc_hd__o21ai_0 _38790_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[21] ),
    .A2(net2248),
    .B1(net2112),
    .Y(_17229_));
 sky130_fd_sc_hd__a21oi_1 _38791_ (.A1(_17226_),
    .A2(_17227_),
    .B1(_17229_),
    .Y(_04755_));
 sky130_fd_sc_hd__a21oi_1 _38792_ (.A1(net1260),
    .A2(net1996),
    .B1(net1908),
    .Y(_17230_));
 sky130_fd_sc_hd__nand2_1 _38793_ (.A(_13850_),
    .B(net1859),
    .Y(_17231_));
 sky130_fd_sc_hd__o21ai_0 _38794_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[22] ),
    .A2(net2264),
    .B1(net2113),
    .Y(_17232_));
 sky130_fd_sc_hd__a21oi_1 _38795_ (.A1(_17230_),
    .A2(_17231_),
    .B1(_17232_),
    .Y(_04756_));
 sky130_fd_sc_hd__nand2_1 _38796_ (.A(_13895_),
    .B(net1857),
    .Y(_17233_));
 sky130_fd_sc_hd__a21oi_1 _38797_ (.A1(net1276),
    .A2(net1994),
    .B1(net1908),
    .Y(_17234_));
 sky130_fd_sc_hd__o21ai_0 _38798_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[23] ),
    .A2(net2263),
    .B1(net2112),
    .Y(_17235_));
 sky130_fd_sc_hd__a21oi_1 _38799_ (.A1(_17233_),
    .A2(_17234_),
    .B1(_17235_),
    .Y(_04757_));
 sky130_fd_sc_hd__nand2_1 _38800_ (.A(_13940_),
    .B(net1857),
    .Y(_17236_));
 sky130_fd_sc_hd__a21oi_1 _38801_ (.A1(net1272),
    .A2(net1994),
    .B1(net1905),
    .Y(_17237_));
 sky130_fd_sc_hd__o21ai_0 _38802_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[24] ),
    .A2(net2248),
    .B1(net2111),
    .Y(_17238_));
 sky130_fd_sc_hd__a21oi_1 _38803_ (.A1(_17236_),
    .A2(_17237_),
    .B1(_17238_),
    .Y(_04758_));
 sky130_fd_sc_hd__o21ai_0 _38804_ (.A1(\inst$top.soc.cpu.sink__payload$18[23] ),
    .A2(net2243),
    .B1(net2104),
    .Y(_17239_));
 sky130_fd_sc_hd__a21oi_1 _38805_ (.A1(_05749_),
    .A2(net2243),
    .B1(_17239_),
    .Y(_04759_));
 sky130_fd_sc_hd__a21oi_1 _38806_ (.A1(net1256),
    .A2(net1996),
    .B1(net1908),
    .Y(_17240_));
 sky130_fd_sc_hd__nand2_1 _38807_ (.A(_13995_),
    .B(net1859),
    .Y(_17241_));
 sky130_fd_sc_hd__o21ai_0 _38808_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[25] ),
    .A2(net2263),
    .B1(net2112),
    .Y(_17242_));
 sky130_fd_sc_hd__a21oi_1 _38809_ (.A1(_17240_),
    .A2(_17241_),
    .B1(_17242_),
    .Y(_04760_));
 sky130_fd_sc_hd__a21oi_1 _38810_ (.A1(net1253),
    .A2(net1995),
    .B1(net1908),
    .Y(_17243_));
 sky130_fd_sc_hd__nand2_1 _38811_ (.A(_14051_),
    .B(net1859),
    .Y(_17244_));
 sky130_fd_sc_hd__o21ai_0 _38814_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[26] ),
    .A2(net2264),
    .B1(net2113),
    .Y(_17247_));
 sky130_fd_sc_hd__a21oi_1 _38815_ (.A1(_17243_),
    .A2(_17244_),
    .B1(_17247_),
    .Y(_04761_));
 sky130_fd_sc_hd__nand2_1 _38816_ (.A(_14111_),
    .B(net1857),
    .Y(_17248_));
 sky130_fd_sc_hd__a21oi_1 _38817_ (.A1(net1453),
    .A2(net1994),
    .B1(net1898),
    .Y(_17249_));
 sky130_fd_sc_hd__o21ai_0 _38818_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[27] ),
    .A2(net2260),
    .B1(net2109),
    .Y(_17250_));
 sky130_fd_sc_hd__a21oi_1 _38819_ (.A1(_17248_),
    .A2(_17249_),
    .B1(_17250_),
    .Y(_04762_));
 sky130_fd_sc_hd__a21oi_1 _38820_ (.A1(net1460),
    .A2(net1995),
    .B1(net1908),
    .Y(_17251_));
 sky130_fd_sc_hd__nand2_1 _38821_ (.A(_14156_),
    .B(net1859),
    .Y(_17252_));
 sky130_fd_sc_hd__o21ai_0 _38822_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[28] ),
    .A2(net2263),
    .B1(net2113),
    .Y(_17253_));
 sky130_fd_sc_hd__a21oi_1 _38823_ (.A1(_17251_),
    .A2(_17252_),
    .B1(_17253_),
    .Y(_04763_));
 sky130_fd_sc_hd__a21oi_1 _38824_ (.A1(net1468),
    .A2(net1995),
    .B1(net1905),
    .Y(_17254_));
 sky130_fd_sc_hd__nand2_1 _38825_ (.A(_14217_),
    .B(net1859),
    .Y(_17255_));
 sky130_fd_sc_hd__o21ai_0 _38826_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[29] ),
    .A2(net2248),
    .B1(net2111),
    .Y(_17256_));
 sky130_fd_sc_hd__a21oi_1 _38827_ (.A1(_17254_),
    .A2(_17255_),
    .B1(_17256_),
    .Y(_04764_));
 sky130_fd_sc_hd__nand2_1 _38828_ (.A(_14306_),
    .B(net1857),
    .Y(_17257_));
 sky130_fd_sc_hd__a21oi_1 _38829_ (.A1(net1475),
    .A2(net1994),
    .B1(net1907),
    .Y(_17258_));
 sky130_fd_sc_hd__o21ai_0 _38831_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[30] ),
    .A2(net2261),
    .B1(net2109),
    .Y(_17260_));
 sky130_fd_sc_hd__a21oi_1 _38832_ (.A1(_17257_),
    .A2(_17258_),
    .B1(_17260_),
    .Y(_04765_));
 sky130_fd_sc_hd__a21oi_1 _38833_ (.A1(net1482),
    .A2(net1995),
    .B1(net1907),
    .Y(_17261_));
 sky130_fd_sc_hd__nand2_1 _38834_ (.A(_14346_),
    .B(net1857),
    .Y(_17262_));
 sky130_fd_sc_hd__o21ai_0 _38835_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[31] ),
    .A2(net2262),
    .B1(net2110),
    .Y(_17263_));
 sky130_fd_sc_hd__a21oi_1 _38836_ (.A1(_17261_),
    .A2(_17262_),
    .B1(_17263_),
    .Y(_04766_));
 sky130_fd_sc_hd__o21ai_0 _38837_ (.A1(\inst$top.soc.cpu.d.sink__payload.mret ),
    .A2(net1901),
    .B1(net2078),
    .Y(_17264_));
 sky130_fd_sc_hd__a21oi_1 _38838_ (.A1(net2544),
    .A2(net1894),
    .B1(_17264_),
    .Y(_04767_));
 sky130_fd_sc_hd__o21ai_0 _38839_ (.A1(\inst$top.soc.cpu.sink__payload$18[24] ),
    .A2(net2244),
    .B1(net2107),
    .Y(_17265_));
 sky130_fd_sc_hd__a21oi_1 _38840_ (.A1(_05768_),
    .A2(net2244),
    .B1(_17265_),
    .Y(_04768_));
 sky130_fd_sc_hd__o21ai_0 _38841_ (.A1(\inst$top.soc.cpu.sink__payload$18[25] ),
    .A2(net2223),
    .B1(net2084),
    .Y(_17266_));
 sky130_fd_sc_hd__a21oi_1 _38842_ (.A1(_12384_),
    .A2(net2223),
    .B1(_17266_),
    .Y(_04769_));
 sky130_fd_sc_hd__o21ai_0 _38844_ (.A1(\inst$top.soc.cpu.sink__payload$18[26] ),
    .A2(net2244),
    .B1(net2106),
    .Y(_17268_));
 sky130_fd_sc_hd__a21oi_1 _38845_ (.A1(_12420_),
    .A2(net2245),
    .B1(_17268_),
    .Y(_04770_));
 sky130_fd_sc_hd__o21ai_0 _38847_ (.A1(\inst$top.soc.cpu.sink__payload$18[27] ),
    .A2(net2244),
    .B1(net2107),
    .Y(_17270_));
 sky130_fd_sc_hd__a21oi_1 _38848_ (.A1(_19947_),
    .A2(net2245),
    .B1(_17270_),
    .Y(_04771_));
 sky130_fd_sc_hd__o21ai_0 _38849_ (.A1(\inst$top.soc.cpu.sink__payload$18[28] ),
    .A2(net2244),
    .B1(net2107),
    .Y(_17271_));
 sky130_fd_sc_hd__a21oi_1 _38850_ (.A1(_12481_),
    .A2(net2245),
    .B1(_17271_),
    .Y(_04772_));
 sky130_fd_sc_hd__o21ai_0 _38851_ (.A1(\inst$top.soc.cpu.sink__payload$18[29] ),
    .A2(net2243),
    .B1(net2107),
    .Y(_17272_));
 sky130_fd_sc_hd__a21oi_1 _38852_ (.A1(_19920_),
    .A2(net2245),
    .B1(_17272_),
    .Y(_04773_));
 sky130_fd_sc_hd__o21ai_0 _38853_ (.A1(\inst$top.soc.cpu.sink__payload$18[2] ),
    .A2(net2217),
    .B1(net2033),
    .Y(_17273_));
 sky130_fd_sc_hd__a21oi_1 _38854_ (.A1(_20462_),
    .A2(net2217),
    .B1(_17273_),
    .Y(_04774_));
 sky130_fd_sc_hd__o21ai_0 _38855_ (.A1(\inst$top.soc.cpu.sink__payload$18[30] ),
    .A2(net2243),
    .B1(net2107),
    .Y(_17274_));
 sky130_fd_sc_hd__a21oi_1 _38856_ (.A1(_19900_),
    .A2(net2243),
    .B1(_17274_),
    .Y(_04775_));
 sky130_fd_sc_hd__o21ai_0 _38858_ (.A1(\inst$top.soc.cpu.sink__payload$18[31] ),
    .A2(net2216),
    .B1(net2031),
    .Y(_17276_));
 sky130_fd_sc_hd__a21oi_1 _38859_ (.A1(_19869_),
    .A2(net2216),
    .B1(_17276_),
    .Y(_04776_));
 sky130_fd_sc_hd__nor2_1 _38860_ (.A(\inst$top.soc.cpu.sink__payload$12[32] ),
    .B(net1889),
    .Y(_17277_));
 sky130_fd_sc_hd__o21ai_0 _38861_ (.A1(\inst$top.soc.cpu.sink__payload$18[32] ),
    .A2(net2228),
    .B1(net2044),
    .Y(_17278_));
 sky130_fd_sc_hd__nor2_1 _38862_ (.A(_17277_),
    .B(_17278_),
    .Y(_04777_));
 sky130_fd_sc_hd__nor2_1 _38863_ (.A(\inst$top.soc.cpu.sink__payload$12[33] ),
    .B(net1889),
    .Y(_17279_));
 sky130_fd_sc_hd__o21ai_0 _38865_ (.A1(\inst$top.soc.cpu.sink__payload$18[33] ),
    .A2(net2228),
    .B1(net2044),
    .Y(_17281_));
 sky130_fd_sc_hd__nor2_1 _38866_ (.A(_17279_),
    .B(_17281_),
    .Y(_04778_));
 sky130_fd_sc_hd__o21ai_0 _38869_ (.A1(\inst$top.soc.cpu.sink__payload$12[34] ),
    .A2(net1886),
    .B1(net2036),
    .Y(_17284_));
 sky130_fd_sc_hd__a21oi_1 _38870_ (.A1(_11842_),
    .A2(net1886),
    .B1(_17284_),
    .Y(_04779_));
 sky130_fd_sc_hd__nor2_1 _38871_ (.A(\inst$top.soc.cpu.sink__payload$12[35] ),
    .B(net1890),
    .Y(_17285_));
 sky130_fd_sc_hd__o21ai_0 _38872_ (.A1(\inst$top.soc.cpu.sink__payload$18[35] ),
    .A2(net2237),
    .B1(net2033),
    .Y(_17286_));
 sky130_fd_sc_hd__nor2_1 _38873_ (.A(_17285_),
    .B(_17286_),
    .Y(_04780_));
 sky130_fd_sc_hd__o21ai_0 _38874_ (.A1(\inst$top.soc.cpu.sink__payload$12[36] ),
    .A2(net1890),
    .B1(net2044),
    .Y(_17287_));
 sky130_fd_sc_hd__a21oi_1 _38875_ (.A1(_11864_),
    .A2(net1881),
    .B1(_17287_),
    .Y(_04781_));
 sky130_fd_sc_hd__o21ai_0 _38876_ (.A1(\inst$top.soc.cpu.sink__payload$12[37] ),
    .A2(net1888),
    .B1(net2042),
    .Y(_17288_));
 sky130_fd_sc_hd__a21oi_1 _38877_ (.A1(_11869_),
    .A2(net1888),
    .B1(_17288_),
    .Y(_04782_));
 sky130_fd_sc_hd__o21ai_0 _38878_ (.A1(\inst$top.soc.cpu.sink__payload$12[38] ),
    .A2(net1887),
    .B1(net2042),
    .Y(_17289_));
 sky130_fd_sc_hd__a21oi_1 _38879_ (.A1(_11874_),
    .A2(net1887),
    .B1(_17289_),
    .Y(_04783_));
 sky130_fd_sc_hd__nor2_1 _38880_ (.A(\inst$top.soc.cpu.sink__payload$12[3] ),
    .B(net1885),
    .Y(_17290_));
 sky130_fd_sc_hd__o21ai_0 _38881_ (.A1(\inst$top.soc.cpu.sink__payload$18[3] ),
    .A2(net2218),
    .B1(net2034),
    .Y(_17291_));
 sky130_fd_sc_hd__nor2_1 _38882_ (.A(_17290_),
    .B(_17291_),
    .Y(_04784_));
 sky130_fd_sc_hd__o21ai_0 _38884_ (.A1(\inst$top.soc.cpu.sink__payload$12[101] ),
    .A2(net1913),
    .B1(net2147),
    .Y(_17293_));
 sky130_fd_sc_hd__a21oi_1 _38885_ (.A1(_11750_),
    .A2(net1913),
    .B1(_17293_),
    .Y(_04785_));
 sky130_fd_sc_hd__o21ai_0 _38886_ (.A1(\inst$top.soc.cpu.sink__payload$18[48] ),
    .A2(net2229),
    .B1(net2045),
    .Y(_17294_));
 sky130_fd_sc_hd__a21oi_1 _38887_ (.A1(_20118_),
    .A2(net2228),
    .B1(_17294_),
    .Y(_04786_));
 sky130_fd_sc_hd__o21ai_0 _38888_ (.A1(\inst$top.soc.cpu.sink__payload$12[103] ),
    .A2(net1911),
    .B1(net2148),
    .Y(_17295_));
 sky130_fd_sc_hd__a21oi_1 _38889_ (.A1(_11762_),
    .A2(net1911),
    .B1(_17295_),
    .Y(_04787_));
 sky130_fd_sc_hd__nor2_1 _38890_ (.A(\inst$top.soc.cpu.sink__payload$12[4] ),
    .B(net1881),
    .Y(_17296_));
 sky130_fd_sc_hd__o21ai_0 _38891_ (.A1(\inst$top.soc.cpu.sink__payload$18[4] ),
    .A2(net2217),
    .B1(net2033),
    .Y(_17297_));
 sky130_fd_sc_hd__nor2_1 _38892_ (.A(_17296_),
    .B(_17297_),
    .Y(_04788_));
 sky130_fd_sc_hd__o21ai_0 _38893_ (.A1(\inst$top.soc.cpu.sink__payload$12[104] ),
    .A2(net1910),
    .B1(net2148),
    .Y(_17298_));
 sky130_fd_sc_hd__a21oi_1 _38894_ (.A1(_11768_),
    .A2(net1910),
    .B1(_17298_),
    .Y(_04789_));
 sky130_fd_sc_hd__o21ai_0 _38895_ (.A1(\inst$top.soc.cpu.sink__payload$12[105] ),
    .A2(net1911),
    .B1(net2148),
    .Y(_17299_));
 sky130_fd_sc_hd__a21oi_1 _38896_ (.A1(_11774_),
    .A2(net1911),
    .B1(_17299_),
    .Y(_04790_));
 sky130_fd_sc_hd__o21ai_0 _38897_ (.A1(\inst$top.soc.cpu.sink__payload$12[52] ),
    .A2(net1891),
    .B1(net2093),
    .Y(_17300_));
 sky130_fd_sc_hd__a21oi_1 _38898_ (.A1(_11784_),
    .A2(net1891),
    .B1(_17300_),
    .Y(_04791_));
 sky130_fd_sc_hd__o21ai_0 _38899_ (.A1(\inst$top.soc.cpu.sink__payload$12[53] ),
    .A2(net1903),
    .B1(net2080),
    .Y(_17301_));
 sky130_fd_sc_hd__a21oi_1 _38900_ (.A1(_11790_),
    .A2(net1903),
    .B1(_17301_),
    .Y(_04792_));
 sky130_fd_sc_hd__o21ai_1 _38903_ (.A1(\inst$top.soc.cpu.sink__payload$12[54] ),
    .A2(net1911),
    .B1(net2178),
    .Y(_17304_));
 sky130_fd_sc_hd__a21oi_1 _38904_ (.A1(_11796_),
    .A2(net1905),
    .B1(_17304_),
    .Y(_04793_));
 sky130_fd_sc_hd__o21ai_0 _38905_ (.A1(\inst$top.soc.cpu.sink__payload$12[55] ),
    .A2(net1897),
    .B1(net2107),
    .Y(_17305_));
 sky130_fd_sc_hd__a21oi_1 _38906_ (.A1(_11801_),
    .A2(net1897),
    .B1(_17305_),
    .Y(_04794_));
 sky130_fd_sc_hd__o21ai_0 _38907_ (.A1(\inst$top.soc.cpu.sink__payload$12[56] ),
    .A2(net1905),
    .B1(net2111),
    .Y(_17306_));
 sky130_fd_sc_hd__a21oi_1 _38908_ (.A1(_11806_),
    .A2(net1905),
    .B1(_17306_),
    .Y(_04795_));
 sky130_fd_sc_hd__o21ai_0 _38910_ (.A1(\inst$top.soc.cpu.sink__payload$12[57] ),
    .A2(net1882),
    .B1(net2031),
    .Y(_17308_));
 sky130_fd_sc_hd__a21oi_1 _38911_ (.A1(_11811_),
    .A2(net1882),
    .B1(_17308_),
    .Y(_04796_));
 sky130_fd_sc_hd__o21ai_0 _38912_ (.A1(\inst$top.soc.cpu.sink__payload$12[58] ),
    .A2(net1902),
    .B1(net2079),
    .Y(_17309_));
 sky130_fd_sc_hd__a21oi_1 _38913_ (.A1(_11818_),
    .A2(net1902),
    .B1(_17309_),
    .Y(_04797_));
 sky130_fd_sc_hd__o21ai_0 _38914_ (.A1(\inst$top.soc.cpu.sink__payload$12[59] ),
    .A2(net1901),
    .B1(net2078),
    .Y(_17310_));
 sky130_fd_sc_hd__a21oi_1 _38915_ (.A1(_11824_),
    .A2(net1901),
    .B1(_17310_),
    .Y(_04798_));
 sky130_fd_sc_hd__o21ai_0 _38916_ (.A1(\inst$top.soc.cpu.sink__payload$18[5] ),
    .A2(net2226),
    .B1(net2042),
    .Y(_17311_));
 sky130_fd_sc_hd__a21oi_1 _38917_ (.A1(_20566_),
    .A2(net2226),
    .B1(_17311_),
    .Y(_04799_));
 sky130_fd_sc_hd__o21ai_0 _38918_ (.A1(\inst$top.soc.cpu.sink__payload$12[60] ),
    .A2(net1902),
    .B1(net2078),
    .Y(_17312_));
 sky130_fd_sc_hd__a21oi_1 _38919_ (.A1(_11830_),
    .A2(net1901),
    .B1(_17312_),
    .Y(_04800_));
 sky130_fd_sc_hd__o21ai_0 _38920_ (.A1(\inst$top.soc.cpu.sink__payload$12[61] ),
    .A2(net1895),
    .B1(net2071),
    .Y(_17313_));
 sky130_fd_sc_hd__a21oi_1 _38921_ (.A1(_11836_),
    .A2(net1895),
    .B1(_17313_),
    .Y(_04801_));
 sky130_fd_sc_hd__o21ai_0 _38922_ (.A1(\inst$top.soc.cpu.sink__payload$12[62] ),
    .A2(net1901),
    .B1(net2071),
    .Y(_17314_));
 sky130_fd_sc_hd__a21oi_1 _38923_ (.A1(_11848_),
    .A2(net1897),
    .B1(_17314_),
    .Y(_04802_));
 sky130_fd_sc_hd__o21ai_0 _38924_ (.A1(\inst$top.soc.cpu.sink__payload$12[63] ),
    .A2(net1882),
    .B1(net2031),
    .Y(_17315_));
 sky130_fd_sc_hd__a21oi_1 _38925_ (.A1(_11853_),
    .A2(net1882),
    .B1(_17315_),
    .Y(_04803_));
 sky130_fd_sc_hd__o21ai_0 _38926_ (.A1(\inst$top.soc.cpu.sink__payload$18[6] ),
    .A2(net2226),
    .B1(net2042),
    .Y(_17316_));
 sky130_fd_sc_hd__a21oi_1 _38927_ (.A1(_20594_),
    .A2(net2226),
    .B1(_17316_),
    .Y(_04804_));
 sky130_fd_sc_hd__o21ai_0 _38929_ (.A1(\inst$top.soc.cpu.sink__payload$18[7] ),
    .A2(net2219),
    .B1(net2032),
    .Y(_17318_));
 sky130_fd_sc_hd__a21oi_1 _38930_ (.A1(_20623_),
    .A2(net2219),
    .B1(_17318_),
    .Y(_04805_));
 sky130_fd_sc_hd__o21ai_0 _38932_ (.A1(\inst$top.soc.cpu.sink__payload$18[8] ),
    .A2(net2239),
    .B1(net2068),
    .Y(_17320_));
 sky130_fd_sc_hd__a21oi_1 _38933_ (.A1(_20664_),
    .A2(net2239),
    .B1(_17320_),
    .Y(_04806_));
 sky130_fd_sc_hd__o21ai_2 _38934_ (.A1(\inst$top.soc.cpu.d.sink__payload.illegal ),
    .A2(net1901),
    .B1(net2079),
    .Y(_17321_));
 sky130_fd_sc_hd__a21oi_1 _38935_ (.A1(_20212_),
    .A2(net1887),
    .B1(_17321_),
    .Y(_04807_));
 sky130_fd_sc_hd__o21ai_0 _38936_ (.A1(_03083_),
    .A2(_13681_),
    .B1(_14886_),
    .Y(_17322_));
 sky130_fd_sc_hd__nor2_1 _38937_ (.A(_15001_),
    .B(net1913),
    .Y(_17323_));
 sky130_fd_sc_hd__o21ai_0 _38938_ (.A1(\inst$top.soc.cpu.d.sink__payload$6.loadstore_misaligned ),
    .A2(net2276),
    .B1(net2080),
    .Y(_17324_));
 sky130_fd_sc_hd__a21oi_1 _38939_ (.A1(_17322_),
    .A2(_17323_),
    .B1(_17324_),
    .Y(_04808_));
 sky130_fd_sc_hd__nor2_1 _38941_ (.A(\inst$top.soc.cpu.d.sink__payload.ecall ),
    .B(net1903),
    .Y(_17326_));
 sky130_fd_sc_hd__o21ai_0 _38943_ (.A1(\inst$top.soc.cpu.d.sink__payload$6.ecall ),
    .A2(net2247),
    .B1(net2079),
    .Y(_17328_));
 sky130_fd_sc_hd__nor2_1 _38944_ (.A(_17326_),
    .B(_17328_),
    .Y(_04809_));
 sky130_fd_sc_hd__nor2_2 _38945_ (.A(\inst$top.soc.cpu.d.sink__payload.ebreak ),
    .B(net1902),
    .Y(_17329_));
 sky130_fd_sc_hd__o21ai_0 _38946_ (.A1(\inst$top.soc.cpu.d.sink__payload$6.ebreak ),
    .A2(net2227),
    .B1(net2042),
    .Y(_17330_));
 sky130_fd_sc_hd__nor2_1 _38947_ (.A(_17329_),
    .B(_17330_),
    .Y(_04810_));
 sky130_fd_sc_hd__o21ai_0 _38948_ (.A1(\inst$top.soc.cpu.sink__payload$18[39] ),
    .A2(net2275),
    .B1(net2150),
    .Y(_17331_));
 sky130_fd_sc_hd__a21oi_1 _38949_ (.A1(_20321_),
    .A2(net2275),
    .B1(_17331_),
    .Y(_04811_));
 sky130_fd_sc_hd__o21ai_0 _38950_ (.A1(\inst$top.soc.cpu.sink__payload$18[9] ),
    .A2(net2228),
    .B1(net2044),
    .Y(_17332_));
 sky130_fd_sc_hd__a21oi_1 _38951_ (.A1(_20685_),
    .A2(net2228),
    .B1(_17332_),
    .Y(_04812_));
 sky130_fd_sc_hd__o21ai_0 _38952_ (.A1(\inst$top.soc.cpu.sink__payload$24[100] ),
    .A2(net2268),
    .B1(net2136),
    .Y(_17333_));
 sky130_fd_sc_hd__a21oi_1 _38953_ (.A1(_15072_),
    .A2(net2268),
    .B1(_17333_),
    .Y(_04813_));
 sky130_fd_sc_hd__o21ai_0 _38955_ (.A1(\inst$top.soc.cpu.sink__payload$24[101] ),
    .A2(net2265),
    .B1(net2130),
    .Y(_17335_));
 sky130_fd_sc_hd__a21oi_1 _38956_ (.A1(_15075_),
    .A2(net2265),
    .B1(_17335_),
    .Y(_04814_));
 sky130_fd_sc_hd__o21ai_0 _38957_ (.A1(\inst$top.soc.cpu.sink__payload$24[102] ),
    .A2(net2265),
    .B1(net2130),
    .Y(_17336_));
 sky130_fd_sc_hd__a21oi_1 _38958_ (.A1(_15079_),
    .A2(net2266),
    .B1(_17336_),
    .Y(_04815_));
 sky130_fd_sc_hd__o21ai_0 _38959_ (.A1(\inst$top.soc.cpu.sink__payload$24[103] ),
    .A2(net2272),
    .B1(net2138),
    .Y(_17337_));
 sky130_fd_sc_hd__a21oi_1 _38960_ (.A1(_15082_),
    .A2(net2271),
    .B1(_17337_),
    .Y(_04816_));
 sky130_fd_sc_hd__o21ai_0 _38961_ (.A1(\inst$top.soc.cpu.sink__payload$24[104] ),
    .A2(net2272),
    .B1(net2138),
    .Y(_17338_));
 sky130_fd_sc_hd__a21oi_1 _38962_ (.A1(_15088_),
    .A2(net2271),
    .B1(_17338_),
    .Y(_04817_));
 sky130_fd_sc_hd__o21ai_0 _38964_ (.A1(\inst$top.soc.cpu.sink__payload$24[105] ),
    .A2(net2270),
    .B1(net2150),
    .Y(_17340_));
 sky130_fd_sc_hd__a21oi_1 _38965_ (.A1(_15092_),
    .A2(net2270),
    .B1(_17340_),
    .Y(_04818_));
 sky130_fd_sc_hd__nor2_1 _38966_ (.A(\inst$top.soc.cpu.d.sink__payload$6.csr_we ),
    .B(net1895),
    .Y(_17341_));
 sky130_fd_sc_hd__o21ai_0 _38967_ (.A1(\inst$top.soc.cpu.d.sink__payload$16.csr_we ),
    .A2(net2238),
    .B1(net2065),
    .Y(_17342_));
 sky130_fd_sc_hd__nor2_1 _38968_ (.A(_17341_),
    .B(_17342_),
    .Y(_04819_));
 sky130_fd_sc_hd__nor2_1 _38969_ (.A(\inst$top.soc.cpu.exception.csr_bank.mie_m_select ),
    .B(\inst$top.soc.cpu.exception.csr_bank.mstatus_m_select ),
    .Y(_17343_));
 sky130_fd_sc_hd__nand3_1 _38970_ (.A(_17343_),
    .B(_11568_),
    .C(_11370_),
    .Y(_17344_));
 sky130_fd_sc_hd__o311ai_0 _38971_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mepc_m_select ),
    .A2(\inst$top.soc.cpu.exception.csr_bank.mtval_m_select ),
    .A3(_17344_),
    .B1(\inst$top.soc.cpu.csrf.bank_300_m_select ),
    .C1(net2220),
    .Y(_17345_));
 sky130_fd_sc_hd__nand2_1 _38972_ (.A(net1883),
    .B(\inst$top.soc.cpu.d.sink__payload$16.csr_rdy ),
    .Y(_17346_));
 sky130_fd_sc_hd__a21oi_1 _38973_ (.A1(_17345_),
    .A2(_17346_),
    .B1(net2957),
    .Y(_04820_));
 sky130_fd_sc_hd__nor2_1 _38974_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[0] ),
    .B(net1906),
    .Y(_17347_));
 sky130_fd_sc_hd__o21ai_0 _38975_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[0] ),
    .A2(net2264),
    .B1(net2113),
    .Y(_17348_));
 sky130_fd_sc_hd__nor2_1 _38976_ (.A(_17347_),
    .B(_17348_),
    .Y(_04821_));
 sky130_fd_sc_hd__nor2_1 _38977_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[1] ),
    .B(net1885),
    .Y(_17349_));
 sky130_fd_sc_hd__o21ai_0 _38978_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[1] ),
    .A2(net2254),
    .B1(net2087),
    .Y(_17350_));
 sky130_fd_sc_hd__nor2_1 _38979_ (.A(_17349_),
    .B(_17350_),
    .Y(_04822_));
 sky130_fd_sc_hd__nor2_1 _38980_ (.A(\inst$top.soc.cpu.sink__payload$18[10] ),
    .B(net1897),
    .Y(_17351_));
 sky130_fd_sc_hd__o21ai_0 _38981_ (.A1(\inst$top.soc.cpu.sink__payload$24[10] ),
    .A2(net2240),
    .B1(net2069),
    .Y(_17352_));
 sky130_fd_sc_hd__nor2_1 _38982_ (.A(_17351_),
    .B(_17352_),
    .Y(_04823_));
 sky130_fd_sc_hd__nor2_1 _38983_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[2] ),
    .B(net1885),
    .Y(_17353_));
 sky130_fd_sc_hd__o21ai_0 _38985_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[2] ),
    .A2(net2218),
    .B1(net2034),
    .Y(_17355_));
 sky130_fd_sc_hd__nor2_1 _38986_ (.A(_17353_),
    .B(_17355_),
    .Y(_04824_));
 sky130_fd_sc_hd__nor2_1 _38987_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[3] ),
    .B(net1885),
    .Y(_17356_));
 sky130_fd_sc_hd__o21ai_0 _38988_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[3] ),
    .A2(net2225),
    .B1(net2088),
    .Y(_17357_));
 sky130_fd_sc_hd__nor2_1 _38989_ (.A(_17356_),
    .B(_17357_),
    .Y(_04825_));
 sky130_fd_sc_hd__nor2_2 _38990_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[4] ),
    .B(net1897),
    .Y(_17358_));
 sky130_fd_sc_hd__o21ai_0 _38991_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[4] ),
    .A2(net2218),
    .B1(net2034),
    .Y(_17359_));
 sky130_fd_sc_hd__nor2_1 _38992_ (.A(_17358_),
    .B(_17359_),
    .Y(_04826_));
 sky130_fd_sc_hd__nor2_1 _38993_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[5] ),
    .B(net1901),
    .Y(_17360_));
 sky130_fd_sc_hd__o21ai_0 _38994_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[5] ),
    .A2(net2247),
    .B1(net2071),
    .Y(_17361_));
 sky130_fd_sc_hd__nor2_1 _38995_ (.A(_17360_),
    .B(_17361_),
    .Y(_04827_));
 sky130_fd_sc_hd__nor2_2 _38997_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[6] ),
    .B(net1906),
    .Y(_17363_));
 sky130_fd_sc_hd__o21ai_0 _38999_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[6] ),
    .A2(net2227),
    .B1(net2043),
    .Y(_17365_));
 sky130_fd_sc_hd__nor2_1 _39000_ (.A(_17363_),
    .B(_17365_),
    .Y(_04828_));
 sky130_fd_sc_hd__nor2_1 _39001_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[7] ),
    .B(net1900),
    .Y(_17366_));
 sky130_fd_sc_hd__o21ai_0 _39002_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[7] ),
    .A2(net2224),
    .B1(net2087),
    .Y(_17367_));
 sky130_fd_sc_hd__nor2_1 _39003_ (.A(_17366_),
    .B(_17367_),
    .Y(_04829_));
 sky130_fd_sc_hd__nor2_1 _39004_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[8] ),
    .B(net1904),
    .Y(_17368_));
 sky130_fd_sc_hd__o21ai_0 _39005_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[8] ),
    .A2(net2241),
    .B1(net2071),
    .Y(_17369_));
 sky130_fd_sc_hd__nor2_1 _39006_ (.A(_17368_),
    .B(_17369_),
    .Y(_04830_));
 sky130_fd_sc_hd__nor2_1 _39007_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[9] ),
    .B(net1894),
    .Y(_17370_));
 sky130_fd_sc_hd__o21ai_0 _39008_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[9] ),
    .A2(net2240),
    .B1(net2070),
    .Y(_17371_));
 sky130_fd_sc_hd__nor2_1 _39009_ (.A(_17370_),
    .B(_17371_),
    .Y(_04831_));
 sky130_fd_sc_hd__nor2_1 _39010_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[10] ),
    .B(net1897),
    .Y(_17372_));
 sky130_fd_sc_hd__o21ai_0 _39011_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[10] ),
    .A2(net2243),
    .B1(net2104),
    .Y(_17373_));
 sky130_fd_sc_hd__nor2_1 _39012_ (.A(_17372_),
    .B(_17373_),
    .Y(_04832_));
 sky130_fd_sc_hd__nor2_1 _39013_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[11] ),
    .B(net1892),
    .Y(_17374_));
 sky130_fd_sc_hd__o21ai_0 _39014_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[11] ),
    .A2(net2232),
    .B1(net2097),
    .Y(_17375_));
 sky130_fd_sc_hd__nor2_1 _39015_ (.A(_17374_),
    .B(_17375_),
    .Y(_04833_));
 sky130_fd_sc_hd__nor2_1 _39016_ (.A(\inst$top.soc.cpu.sink__payload$18[11] ),
    .B(net1891),
    .Y(_17376_));
 sky130_fd_sc_hd__o21ai_0 _39018_ (.A1(\inst$top.soc.cpu.sink__payload$24[11] ),
    .A2(net2230),
    .B1(net2093),
    .Y(_17378_));
 sky130_fd_sc_hd__nor2_1 _39019_ (.A(_17376_),
    .B(_17378_),
    .Y(_04834_));
 sky130_fd_sc_hd__nor2_1 _39020_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[12] ),
    .B(net1897),
    .Y(_17379_));
 sky130_fd_sc_hd__o21ai_0 _39021_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[12] ),
    .A2(net2243),
    .B1(net2070),
    .Y(_17380_));
 sky130_fd_sc_hd__nor2_1 _39022_ (.A(_17379_),
    .B(_17380_),
    .Y(_04835_));
 sky130_fd_sc_hd__nor2_1 _39023_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[13] ),
    .B(net1905),
    .Y(_17381_));
 sky130_fd_sc_hd__o21ai_0 _39024_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[13] ),
    .A2(net2248),
    .B1(net2111),
    .Y(_17382_));
 sky130_fd_sc_hd__nor2_1 _39025_ (.A(_17381_),
    .B(_17382_),
    .Y(_04836_));
 sky130_fd_sc_hd__nor2_1 _39026_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[14] ),
    .B(net1899),
    .Y(_17383_));
 sky130_fd_sc_hd__o21ai_0 _39027_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[14] ),
    .A2(net2240),
    .B1(net2070),
    .Y(_17384_));
 sky130_fd_sc_hd__nor2_1 _39028_ (.A(_17383_),
    .B(_17384_),
    .Y(_04837_));
 sky130_fd_sc_hd__nor2_1 _39030_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[15] ),
    .B(net1895),
    .Y(_17386_));
 sky130_fd_sc_hd__o21ai_0 _39032_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[15] ),
    .A2(net2240),
    .B1(net2070),
    .Y(_17388_));
 sky130_fd_sc_hd__nor2_1 _39033_ (.A(_17386_),
    .B(_17388_),
    .Y(_04838_));
 sky130_fd_sc_hd__nor2_1 _39034_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[16] ),
    .B(net1898),
    .Y(_17389_));
 sky130_fd_sc_hd__o21ai_0 _39035_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[16] ),
    .A2(net2260),
    .B1(net2106),
    .Y(_17390_));
 sky130_fd_sc_hd__nor2_1 _39036_ (.A(_17389_),
    .B(_17390_),
    .Y(_04839_));
 sky130_fd_sc_hd__nor2_1 _39037_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[17] ),
    .B(net1898),
    .Y(_17391_));
 sky130_fd_sc_hd__o21ai_0 _39038_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[17] ),
    .A2(net2260),
    .B1(net2109),
    .Y(_17392_));
 sky130_fd_sc_hd__nor2_1 _39039_ (.A(_17391_),
    .B(_17392_),
    .Y(_04840_));
 sky130_fd_sc_hd__nor2_1 _39040_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[18] ),
    .B(net1907),
    .Y(_17393_));
 sky130_fd_sc_hd__o21ai_0 _39041_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[18] ),
    .A2(net2262),
    .B1(net2110),
    .Y(_17394_));
 sky130_fd_sc_hd__nor2_1 _39042_ (.A(_17393_),
    .B(_17394_),
    .Y(_04841_));
 sky130_fd_sc_hd__nor2_1 _39043_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[19] ),
    .B(net1907),
    .Y(_17395_));
 sky130_fd_sc_hd__o21ai_0 _39044_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[19] ),
    .A2(net2261),
    .B1(net2109),
    .Y(_17396_));
 sky130_fd_sc_hd__nor2_1 _39045_ (.A(_17395_),
    .B(_17396_),
    .Y(_04842_));
 sky130_fd_sc_hd__nor2_1 _39046_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[20] ),
    .B(net1907),
    .Y(_17397_));
 sky130_fd_sc_hd__o21ai_0 _39047_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[20] ),
    .A2(net2262),
    .B1(net2110),
    .Y(_17398_));
 sky130_fd_sc_hd__nor2_1 _39048_ (.A(_17397_),
    .B(_17398_),
    .Y(_04843_));
 sky130_fd_sc_hd__nor2_1 _39049_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[21] ),
    .B(net1905),
    .Y(_17399_));
 sky130_fd_sc_hd__o21ai_0 _39051_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[21] ),
    .A2(net2245),
    .B1(net2108),
    .Y(_17401_));
 sky130_fd_sc_hd__nor2_1 _39052_ (.A(_17399_),
    .B(_17401_),
    .Y(_04844_));
 sky130_fd_sc_hd__nor2_1 _39053_ (.A(\inst$top.soc.cpu.sink__payload$18[12] ),
    .B(net1892),
    .Y(_17402_));
 sky130_fd_sc_hd__o21ai_0 _39054_ (.A1(\inst$top.soc.cpu.sink__payload$24[12] ),
    .A2(net2229),
    .B1(net2045),
    .Y(_17403_));
 sky130_fd_sc_hd__nor2_1 _39055_ (.A(_17402_),
    .B(_17403_),
    .Y(_04845_));
 sky130_fd_sc_hd__nor2_1 _39056_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[22] ),
    .B(net1907),
    .Y(_17404_));
 sky130_fd_sc_hd__o21ai_0 _39057_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[22] ),
    .A2(net2262),
    .B1(net2110),
    .Y(_17405_));
 sky130_fd_sc_hd__nor2_1 _39058_ (.A(_17404_),
    .B(_17405_),
    .Y(_04846_));
 sky130_fd_sc_hd__nor2_1 _39059_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[23] ),
    .B(net1907),
    .Y(_17406_));
 sky130_fd_sc_hd__o21ai_0 _39060_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[23] ),
    .A2(net2261),
    .B1(net2109),
    .Y(_17407_));
 sky130_fd_sc_hd__nor2_1 _39061_ (.A(_17406_),
    .B(_17407_),
    .Y(_04847_));
 sky130_fd_sc_hd__nor2_1 _39063_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[24] ),
    .B(net1898),
    .Y(_17409_));
 sky130_fd_sc_hd__o21ai_0 _39065_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[24] ),
    .A2(net2244),
    .B1(net2106),
    .Y(_17411_));
 sky130_fd_sc_hd__nor2_1 _39066_ (.A(_17409_),
    .B(_17411_),
    .Y(_04848_));
 sky130_fd_sc_hd__nor2_2 _39067_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[25] ),
    .B(net1908),
    .Y(_17412_));
 sky130_fd_sc_hd__o21ai_0 _39068_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[25] ),
    .A2(net2253),
    .B1(net2090),
    .Y(_17413_));
 sky130_fd_sc_hd__nor2_1 _39069_ (.A(_17412_),
    .B(_17413_),
    .Y(_04849_));
 sky130_fd_sc_hd__nor2_1 _39070_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[26] ),
    .B(net1907),
    .Y(_17414_));
 sky130_fd_sc_hd__o21ai_0 _39071_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[26] ),
    .A2(net2261),
    .B1(net2109),
    .Y(_17415_));
 sky130_fd_sc_hd__nor2_1 _39072_ (.A(_17414_),
    .B(_17415_),
    .Y(_04850_));
 sky130_fd_sc_hd__nor2_1 _39073_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[27] ),
    .B(net1898),
    .Y(_17416_));
 sky130_fd_sc_hd__o21ai_0 _39074_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[27] ),
    .A2(net2260),
    .B1(net2109),
    .Y(_17417_));
 sky130_fd_sc_hd__nor2_1 _39075_ (.A(_17416_),
    .B(_17417_),
    .Y(_04851_));
 sky130_fd_sc_hd__nor2_1 _39076_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[28] ),
    .B(net1898),
    .Y(_17418_));
 sky130_fd_sc_hd__o21ai_0 _39077_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[28] ),
    .A2(net2260),
    .B1(net2106),
    .Y(_17419_));
 sky130_fd_sc_hd__nor2_1 _39078_ (.A(_17418_),
    .B(_17419_),
    .Y(_04852_));
 sky130_fd_sc_hd__nor2_1 _39079_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[29] ),
    .B(net1906),
    .Y(_17420_));
 sky130_fd_sc_hd__o21ai_0 _39080_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[29] ),
    .A2(net2248),
    .B1(net2106),
    .Y(_17421_));
 sky130_fd_sc_hd__nor2_1 _39081_ (.A(_17420_),
    .B(_17421_),
    .Y(_04853_));
 sky130_fd_sc_hd__nor2_1 _39082_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[30] ),
    .B(net1907),
    .Y(_17422_));
 sky130_fd_sc_hd__o21ai_0 _39084_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[30] ),
    .A2(net2261),
    .B1(net2109),
    .Y(_17424_));
 sky130_fd_sc_hd__nor2_1 _39085_ (.A(_17422_),
    .B(_17424_),
    .Y(_04854_));
 sky130_fd_sc_hd__nor2_1 _39086_ (.A(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[31] ),
    .B(net1909),
    .Y(_17425_));
 sky130_fd_sc_hd__o21ai_0 _39087_ (.A1(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[31] ),
    .A2(net2253),
    .B1(net2090),
    .Y(_17426_));
 sky130_fd_sc_hd__nor2_1 _39088_ (.A(_17425_),
    .B(_17426_),
    .Y(_04855_));
 sky130_fd_sc_hd__nor2_1 _39089_ (.A(\inst$top.soc.cpu.sink__payload$18[13] ),
    .B(net1900),
    .Y(_17427_));
 sky130_fd_sc_hd__o21ai_0 _39090_ (.A1(\inst$top.soc.cpu.sink__payload$24[13] ),
    .A2(net2242),
    .B1(net2104),
    .Y(_17428_));
 sky130_fd_sc_hd__nor2_1 _39091_ (.A(_17427_),
    .B(_17428_),
    .Y(_04856_));
 sky130_fd_sc_hd__o21ai_0 _39092_ (.A1(\inst$top.soc.cpu.d.sink__payload$6.multiply ),
    .A2(net1915),
    .B1(net2154),
    .Y(_17429_));
 sky130_fd_sc_hd__a21oi_1 _39093_ (.A1(net2196),
    .A2(net1914),
    .B1(_17429_),
    .Y(_04857_));
 sky130_fd_sc_hd__nor2_1 _39094_ (.A(\inst$top.soc.cpu.sink__payload$18[14] ),
    .B(net1896),
    .Y(_17430_));
 sky130_fd_sc_hd__o21ai_0 _39095_ (.A1(\inst$top.soc.cpu.sink__payload$24[14] ),
    .A2(net2239),
    .B1(net2068),
    .Y(_17431_));
 sky130_fd_sc_hd__nor2_1 _39096_ (.A(_17430_),
    .B(_17431_),
    .Y(_04858_));
 sky130_fd_sc_hd__nor2_1 _39098_ (.A(\inst$top.soc.cpu.sink__payload$18[15] ),
    .B(net1894),
    .Y(_17433_));
 sky130_fd_sc_hd__o21ai_0 _39100_ (.A1(\inst$top.soc.cpu.sink__payload$24[15] ),
    .A2(net2241),
    .B1(net2071),
    .Y(_17435_));
 sky130_fd_sc_hd__nor2_1 _39101_ (.A(_17433_),
    .B(_17435_),
    .Y(_04859_));
 sky130_fd_sc_hd__nor2_1 _39102_ (.A(\inst$top.soc.cpu.sink__payload$18[16] ),
    .B(net1891),
    .Y(_17436_));
 sky130_fd_sc_hd__o21ai_0 _39103_ (.A1(\inst$top.soc.cpu.sink__payload$24[16] ),
    .A2(net2230),
    .B1(net2093),
    .Y(_17437_));
 sky130_fd_sc_hd__nor2_1 _39104_ (.A(_17436_),
    .B(_17437_),
    .Y(_04860_));
 sky130_fd_sc_hd__nor2_1 _39105_ (.A(\inst$top.soc.cpu.sink__payload$18[17] ),
    .B(net1892),
    .Y(_17438_));
 sky130_fd_sc_hd__o21ai_0 _39106_ (.A1(\inst$top.soc.cpu.sink__payload$24[17] ),
    .A2(net2257),
    .B1(net2096),
    .Y(_17439_));
 sky130_fd_sc_hd__nor2_1 _39107_ (.A(_17438_),
    .B(_17439_),
    .Y(_04861_));
 sky130_fd_sc_hd__nor2_1 _39108_ (.A(\inst$top.soc.cpu.sink__payload$18[18] ),
    .B(net1892),
    .Y(_17440_));
 sky130_fd_sc_hd__o21ai_0 _39109_ (.A1(\inst$top.soc.cpu.sink__payload$24[18] ),
    .A2(net2231),
    .B1(net2102),
    .Y(_17441_));
 sky130_fd_sc_hd__nor2_1 _39110_ (.A(_17440_),
    .B(_17441_),
    .Y(_04862_));
 sky130_fd_sc_hd__nor2_1 _39111_ (.A(\inst$top.soc.cpu.sink__payload$18[19] ),
    .B(net1892),
    .Y(_17442_));
 sky130_fd_sc_hd__o21ai_0 _39112_ (.A1(\inst$top.soc.cpu.sink__payload$24[19] ),
    .A2(net2231),
    .B1(net2094),
    .Y(_17443_));
 sky130_fd_sc_hd__nor2_1 _39113_ (.A(_17442_),
    .B(_17443_),
    .Y(_04863_));
 sky130_fd_sc_hd__nor2_1 _39114_ (.A(\inst$top.soc.cpu.sink__payload$18[20] ),
    .B(net1891),
    .Y(_17444_));
 sky130_fd_sc_hd__o21ai_0 _39115_ (.A1(\inst$top.soc.cpu.sink__payload$24[20] ),
    .A2(net2255),
    .B1(net2094),
    .Y(_17445_));
 sky130_fd_sc_hd__nor2_1 _39116_ (.A(_17444_),
    .B(_17445_),
    .Y(_04864_));
 sky130_fd_sc_hd__nor2_1 _39117_ (.A(\inst$top.soc.cpu.sink__payload$18[21] ),
    .B(net1891),
    .Y(_17446_));
 sky130_fd_sc_hd__o21ai_0 _39119_ (.A1(\inst$top.soc.cpu.sink__payload$24[21] ),
    .A2(net2230),
    .B1(net2094),
    .Y(_17448_));
 sky130_fd_sc_hd__nor2_1 _39120_ (.A(_17446_),
    .B(_17448_),
    .Y(_04865_));
 sky130_fd_sc_hd__nor2_1 _39121_ (.A(\inst$top.soc.cpu.sink__payload$18[22] ),
    .B(net1900),
    .Y(_17449_));
 sky130_fd_sc_hd__o21ai_0 _39122_ (.A1(\inst$top.soc.cpu.sink__payload$24[22] ),
    .A2(net2262),
    .B1(net2105),
    .Y(_17450_));
 sky130_fd_sc_hd__nor2_1 _39123_ (.A(_17449_),
    .B(_17450_),
    .Y(_04866_));
 sky130_fd_sc_hd__nor2_1 _39124_ (.A(\inst$top.soc.cpu.sink__payload$18[23] ),
    .B(net1897),
    .Y(_17451_));
 sky130_fd_sc_hd__o21ai_0 _39125_ (.A1(\inst$top.soc.cpu.sink__payload$24[23] ),
    .A2(net2262),
    .B1(net2105),
    .Y(_17452_));
 sky130_fd_sc_hd__nor2_1 _39126_ (.A(_17451_),
    .B(_17452_),
    .Y(_04867_));
 sky130_fd_sc_hd__nor2_1 _39127_ (.A(\inst$top.soc.cpu.sink__payload$18[24] ),
    .B(net1898),
    .Y(_17453_));
 sky130_fd_sc_hd__o21ai_0 _39128_ (.A1(\inst$top.soc.cpu.sink__payload$24[24] ),
    .A2(net2244),
    .B1(net2107),
    .Y(_17454_));
 sky130_fd_sc_hd__nor2_1 _39129_ (.A(_17453_),
    .B(_17454_),
    .Y(_04868_));
 sky130_fd_sc_hd__nor2_1 _39131_ (.A(\inst$top.soc.cpu.sink__payload$18[25] ),
    .B(net1885),
    .Y(_17456_));
 sky130_fd_sc_hd__o21ai_0 _39133_ (.A1(\inst$top.soc.cpu.sink__payload$24[25] ),
    .A2(net2252),
    .B1(net2086),
    .Y(_17458_));
 sky130_fd_sc_hd__nor2_1 _39134_ (.A(_17456_),
    .B(_17458_),
    .Y(_04869_));
 sky130_fd_sc_hd__nor2_1 _39135_ (.A(\inst$top.soc.cpu.sink__payload$18[26] ),
    .B(net1899),
    .Y(_17459_));
 sky130_fd_sc_hd__o21ai_0 _39136_ (.A1(\inst$top.soc.cpu.sink__payload$24[26] ),
    .A2(net2261),
    .B1(net2106),
    .Y(_17460_));
 sky130_fd_sc_hd__nor2_1 _39137_ (.A(_17459_),
    .B(_17460_),
    .Y(_04870_));
 sky130_fd_sc_hd__nor2_1 _39138_ (.A(\inst$top.soc.cpu.sink__payload$18[27] ),
    .B(net1898),
    .Y(_17461_));
 sky130_fd_sc_hd__o21ai_0 _39139_ (.A1(\inst$top.soc.cpu.sink__payload$24[27] ),
    .A2(net2244),
    .B1(net2106),
    .Y(_17462_));
 sky130_fd_sc_hd__nor2_1 _39140_ (.A(_17461_),
    .B(_17462_),
    .Y(_04871_));
 sky130_fd_sc_hd__nor2_1 _39141_ (.A(\inst$top.soc.cpu.sink__payload$18[28] ),
    .B(net1898),
    .Y(_17463_));
 sky130_fd_sc_hd__o21ai_0 _39142_ (.A1(\inst$top.soc.cpu.sink__payload$24[28] ),
    .A2(net2244),
    .B1(net2106),
    .Y(_17464_));
 sky130_fd_sc_hd__nor2_1 _39143_ (.A(_17463_),
    .B(_17464_),
    .Y(_04872_));
 sky130_fd_sc_hd__nor2_1 _39144_ (.A(\inst$top.soc.cpu.sink__payload$18[29] ),
    .B(net1899),
    .Y(_17465_));
 sky130_fd_sc_hd__o21ai_0 _39145_ (.A1(\inst$top.soc.cpu.sink__payload$24[29] ),
    .A2(net2243),
    .B1(net2107),
    .Y(_17466_));
 sky130_fd_sc_hd__nor2_1 _39146_ (.A(_17465_),
    .B(_17466_),
    .Y(_04873_));
 sky130_fd_sc_hd__nor2_1 _39147_ (.A(\inst$top.soc.cpu.sink__payload$18[2] ),
    .B(net1886),
    .Y(_17467_));
 sky130_fd_sc_hd__o21ai_0 _39148_ (.A1(\inst$top.soc.cpu.sink__payload$24[2] ),
    .A2(net2217),
    .B1(net2035),
    .Y(_17468_));
 sky130_fd_sc_hd__nor2_1 _39149_ (.A(_17467_),
    .B(_17468_),
    .Y(_04874_));
 sky130_fd_sc_hd__nor2_1 _39150_ (.A(\inst$top.soc.cpu.sink__payload$18[30] ),
    .B(net1899),
    .Y(_17469_));
 sky130_fd_sc_hd__o21ai_0 _39152_ (.A1(\inst$top.soc.cpu.sink__payload$24[30] ),
    .A2(net2243),
    .B1(net2107),
    .Y(_17471_));
 sky130_fd_sc_hd__nor2_1 _39153_ (.A(_17469_),
    .B(_17471_),
    .Y(_04875_));
 sky130_fd_sc_hd__nor2_1 _39154_ (.A(\inst$top.soc.cpu.sink__payload$18[31] ),
    .B(net1882),
    .Y(_17472_));
 sky130_fd_sc_hd__o21ai_0 _39155_ (.A1(\inst$top.soc.cpu.sink__payload$24[31] ),
    .A2(net2216),
    .B1(net2031),
    .Y(_17473_));
 sky130_fd_sc_hd__nor2_1 _39156_ (.A(_17472_),
    .B(_17473_),
    .Y(_04876_));
 sky130_fd_sc_hd__o21ai_0 _39158_ (.A1(\inst$top.soc.cpu.sink__payload$24[32] ),
    .A2(net2286),
    .B1(net2171),
    .Y(_17475_));
 sky130_fd_sc_hd__a21oi_1 _39159_ (.A1(_11880_),
    .A2(net2286),
    .B1(_17475_),
    .Y(_04877_));
 sky130_fd_sc_hd__o21ai_0 _39160_ (.A1(\inst$top.soc.cpu.sink__payload$24[33] ),
    .A2(net2286),
    .B1(net2171),
    .Y(_17476_));
 sky130_fd_sc_hd__a21oi_1 _39161_ (.A1(_11885_),
    .A2(net2286),
    .B1(_17476_),
    .Y(_04878_));
 sky130_fd_sc_hd__o21ai_0 _39162_ (.A1(\inst$top.soc.cpu.sink__payload$24[34] ),
    .A2(net2286),
    .B1(net2171),
    .Y(_17477_));
 sky130_fd_sc_hd__a21oi_1 _39163_ (.A1(_20267_),
    .A2(net2286),
    .B1(_17477_),
    .Y(_04879_));
 sky130_fd_sc_hd__o21ai_0 _39164_ (.A1(\inst$top.soc.cpu.sink__payload$24[35] ),
    .A2(net2286),
    .B1(net2171),
    .Y(_17478_));
 sky130_fd_sc_hd__a21oi_1 _39165_ (.A1(_11724_),
    .A2(net2286),
    .B1(_17478_),
    .Y(_04880_));
 sky130_fd_sc_hd__o21ai_0 _39166_ (.A1(\inst$top.soc.cpu.sink__payload$24[36] ),
    .A2(net2286),
    .B1(net2171),
    .Y(_17479_));
 sky130_fd_sc_hd__a21oi_1 _39167_ (.A1(_20271_),
    .A2(net2286),
    .B1(_17479_),
    .Y(_04881_));
 sky130_fd_sc_hd__nor2_1 _39168_ (.A(\inst$top.soc.cpu.d.sink__payload$6.rd_we ),
    .B(net1913),
    .Y(_17480_));
 sky130_fd_sc_hd__o21ai_0 _39169_ (.A1(\inst$top.soc.cpu.d.sink__payload$16.rd_we ),
    .A2(net2267),
    .B1(net2145),
    .Y(_17481_));
 sky130_fd_sc_hd__nor2_1 _39170_ (.A(_17480_),
    .B(_17481_),
    .Y(_04882_));
 sky130_fd_sc_hd__o21ai_0 _39172_ (.A1(\inst$top.soc.cpu.sink__payload$24[38] ),
    .A2(net2270),
    .B1(net2150),
    .Y(_17483_));
 sky130_fd_sc_hd__a21oi_1 _39173_ (.A1(_11735_),
    .A2(net2270),
    .B1(_17483_),
    .Y(_04883_));
 sky130_fd_sc_hd__o21ai_0 _39174_ (.A1(\inst$top.soc.cpu.sink__payload$24[39] ),
    .A2(net2265),
    .B1(net2144),
    .Y(_17484_));
 sky130_fd_sc_hd__a21oi_1 _39175_ (.A1(_11740_),
    .A2(net2265),
    .B1(_17484_),
    .Y(_04884_));
 sky130_fd_sc_hd__nor2_1 _39176_ (.A(\inst$top.soc.cpu.sink__payload$18[3] ),
    .B(net1885),
    .Y(_17485_));
 sky130_fd_sc_hd__o21ai_0 _39177_ (.A1(\inst$top.soc.cpu.sink__payload$24[3] ),
    .A2(net2225),
    .B1(net2034),
    .Y(_17486_));
 sky130_fd_sc_hd__nor2_1 _39178_ (.A(_17485_),
    .B(_17486_),
    .Y(_04885_));
 sky130_fd_sc_hd__o21ai_0 _39179_ (.A1(\inst$top.soc.cpu.sink__payload$24[40] ),
    .A2(net2265),
    .B1(net2144),
    .Y(_17487_));
 sky130_fd_sc_hd__a21oi_1 _39180_ (.A1(_11745_),
    .A2(net2265),
    .B1(_17487_),
    .Y(_04886_));
 sky130_fd_sc_hd__a21oi_1 _39181_ (.A1(net1915),
    .A2(_20409_),
    .B1(net2994),
    .Y(_17488_));
 sky130_fd_sc_hd__o21ai_0 _39182_ (.A1(net1915),
    .A2(_13006_),
    .B1(_17488_),
    .Y(_17489_));
 sky130_fd_sc_hd__inv_2 _39183_ (.A(_17489_),
    .Y(_04887_));
 sky130_fd_sc_hd__o21ai_0 _39185_ (.A1(net2822),
    .A2(net2270),
    .B1(net2150),
    .Y(_17491_));
 sky130_fd_sc_hd__a21oi_1 _39186_ (.A1(_13676_),
    .A2(net2270),
    .B1(_17491_),
    .Y(_04888_));
 sky130_fd_sc_hd__o21ai_0 _39187_ (.A1(\inst$top.soc.cpu.sink__payload$24[43] ),
    .A2(net2279),
    .B1(net2154),
    .Y(_17492_));
 sky130_fd_sc_hd__a21oi_1 _39188_ (.A1(_14249_),
    .A2(net2279),
    .B1(_17492_),
    .Y(_04889_));
 sky130_fd_sc_hd__o21ai_0 _39190_ (.A1(\inst$top.soc.cpu.sink__payload$24[44] ),
    .A2(net2278),
    .B1(net2157),
    .Y(_17494_));
 sky130_fd_sc_hd__a21oi_1 _39191_ (.A1(_14385_),
    .A2(net2278),
    .B1(_17494_),
    .Y(_04890_));
 sky130_fd_sc_hd__o21ai_0 _39192_ (.A1(\inst$top.soc.cpu.sink__payload$24[45] ),
    .A2(net2279),
    .B1(net2154),
    .Y(_17495_));
 sky130_fd_sc_hd__a21oi_1 _39193_ (.A1(_14399_),
    .A2(net2279),
    .B1(_17495_),
    .Y(_04891_));
 sky130_fd_sc_hd__o21ai_0 _39194_ (.A1(\inst$top.soc.cpu.sink__payload$24[46] ),
    .A2(net2280),
    .B1(net2157),
    .Y(_17496_));
 sky130_fd_sc_hd__a21oi_1 _39195_ (.A1(_14427_),
    .A2(net2281),
    .B1(_17496_),
    .Y(_04892_));
 sky130_fd_sc_hd__o21ai_0 _39196_ (.A1(\inst$top.soc.cpu.sink__payload$24[47] ),
    .A2(net2287),
    .B1(net2171),
    .Y(_17497_));
 sky130_fd_sc_hd__a21oi_1 _39197_ (.A1(_14458_),
    .A2(net2287),
    .B1(_17497_),
    .Y(_04893_));
 sky130_fd_sc_hd__o21ai_0 _39198_ (.A1(\inst$top.soc.cpu.sink__payload$24[48] ),
    .A2(net2274),
    .B1(net2151),
    .Y(_17498_));
 sky130_fd_sc_hd__a21oi_1 _39199_ (.A1(_14501_),
    .A2(net2274),
    .B1(_17498_),
    .Y(_04894_));
 sky130_fd_sc_hd__o21ai_0 _39201_ (.A1(\inst$top.soc.cpu.sink__payload$24[49] ),
    .A2(net2290),
    .B1(net2172),
    .Y(_17500_));
 sky130_fd_sc_hd__a21oi_1 _39202_ (.A1(_14516_),
    .A2(net2290),
    .B1(_17500_),
    .Y(_04895_));
 sky130_fd_sc_hd__nor2_1 _39203_ (.A(\inst$top.soc.cpu.sink__payload$18[4] ),
    .B(net1882),
    .Y(_17501_));
 sky130_fd_sc_hd__o21ai_0 _39204_ (.A1(\inst$top.soc.cpu.sink__payload$24[4] ),
    .A2(net2216),
    .B1(net2031),
    .Y(_17502_));
 sky130_fd_sc_hd__nor2_1 _39205_ (.A(_17501_),
    .B(_17502_),
    .Y(_04896_));
 sky130_fd_sc_hd__o21ai_0 _39206_ (.A1(\inst$top.soc.cpu.sink__payload$24[50] ),
    .A2(net2287),
    .B1(net2172),
    .Y(_17503_));
 sky130_fd_sc_hd__a21oi_1 _39207_ (.A1(_14544_),
    .A2(net2287),
    .B1(_17503_),
    .Y(_04897_));
 sky130_fd_sc_hd__o21ai_0 _39208_ (.A1(\inst$top.soc.cpu.sink__payload$24[51] ),
    .A2(net2280),
    .B1(net2154),
    .Y(_17504_));
 sky130_fd_sc_hd__a21oi_1 _39209_ (.A1(_13027_),
    .A2(net2280),
    .B1(_17504_),
    .Y(_04898_));
 sky130_fd_sc_hd__o21ai_0 _39211_ (.A1(\inst$top.soc.cpu.sink__payload$24[52] ),
    .A2(net2281),
    .B1(net2157),
    .Y(_17506_));
 sky130_fd_sc_hd__a21oi_1 _39212_ (.A1(_13113_),
    .A2(net2281),
    .B1(_17506_),
    .Y(_04899_));
 sky130_fd_sc_hd__o21ai_0 _39213_ (.A1(\inst$top.soc.cpu.sink__payload$24[53] ),
    .A2(net2290),
    .B1(net2174),
    .Y(_17507_));
 sky130_fd_sc_hd__a21oi_1 _39214_ (.A1(_13239_),
    .A2(net2290),
    .B1(_17507_),
    .Y(_04900_));
 sky130_fd_sc_hd__o21ai_0 _39216_ (.A1(\inst$top.soc.cpu.sink__payload$24[54] ),
    .A2(net2280),
    .B1(net2156),
    .Y(_17509_));
 sky130_fd_sc_hd__a21oi_1 _39217_ (.A1(_13255_),
    .A2(net2280),
    .B1(_17509_),
    .Y(_04901_));
 sky130_fd_sc_hd__o21ai_0 _39218_ (.A1(\inst$top.soc.cpu.sink__payload$24[55] ),
    .A2(net2287),
    .B1(net2153),
    .Y(_17510_));
 sky130_fd_sc_hd__nor2_1 _39219_ (.A(net1925),
    .B(_13348_),
    .Y(_17511_));
 sky130_fd_sc_hd__nor2_1 _39220_ (.A(_17510_),
    .B(_17511_),
    .Y(_04902_));
 sky130_fd_sc_hd__o21ai_0 _39221_ (.A1(\inst$top.soc.cpu.sink__payload$24[56] ),
    .A2(net2280),
    .B1(net2154),
    .Y(_17512_));
 sky130_fd_sc_hd__a21oi_1 _39222_ (.A1(_13396_),
    .A2(net2280),
    .B1(_17512_),
    .Y(_04903_));
 sky130_fd_sc_hd__o21ai_0 _39223_ (.A1(\inst$top.soc.cpu.sink__payload$24[57] ),
    .A2(net2281),
    .B1(net2157),
    .Y(_17513_));
 sky130_fd_sc_hd__a21oi_1 _39224_ (.A1(_13411_),
    .A2(net2281),
    .B1(_17513_),
    .Y(_04904_));
 sky130_fd_sc_hd__o21ai_0 _39225_ (.A1(\inst$top.soc.cpu.sink__payload$24[58] ),
    .A2(net2292),
    .B1(net2173),
    .Y(_17514_));
 sky130_fd_sc_hd__nor2_1 _39226_ (.A(net1925),
    .B(_13532_),
    .Y(_17515_));
 sky130_fd_sc_hd__nor2_1 _39227_ (.A(_17514_),
    .B(_17515_),
    .Y(_04905_));
 sky130_fd_sc_hd__o21ai_0 _39228_ (.A1(\inst$top.soc.cpu.sink__payload$24[59] ),
    .A2(net2274),
    .B1(net2151),
    .Y(_17516_));
 sky130_fd_sc_hd__a21oi_1 _39229_ (.A1(_13585_),
    .A2(net2274),
    .B1(_17516_),
    .Y(_04906_));
 sky130_fd_sc_hd__nor2_1 _39230_ (.A(\inst$top.soc.cpu.sink__payload$18[5] ),
    .B(net1887),
    .Y(_17517_));
 sky130_fd_sc_hd__o21ai_0 _39231_ (.A1(\inst$top.soc.cpu.sink__payload$24[5] ),
    .A2(net2226),
    .B1(net2042),
    .Y(_17518_));
 sky130_fd_sc_hd__nor2_1 _39232_ (.A(_17517_),
    .B(_17518_),
    .Y(_04907_));
 sky130_fd_sc_hd__o21ai_0 _39233_ (.A1(\inst$top.soc.cpu.sink__payload$24[60] ),
    .A2(net2289),
    .B1(net2156),
    .Y(_17519_));
 sky130_fd_sc_hd__a21oi_1 _39234_ (.A1(_13606_),
    .A2(net2289),
    .B1(_17519_),
    .Y(_04908_));
 sky130_fd_sc_hd__o21ai_0 _39235_ (.A1(\inst$top.soc.cpu.sink__payload$24[61] ),
    .A2(net2292),
    .B1(net2174),
    .Y(_17520_));
 sky130_fd_sc_hd__nor2_1 _39236_ (.A(net1925),
    .B(_13743_),
    .Y(_17521_));
 sky130_fd_sc_hd__nor2_1 _39237_ (.A(_17520_),
    .B(_17521_),
    .Y(_04909_));
 sky130_fd_sc_hd__o21ai_0 _39239_ (.A1(\inst$top.soc.cpu.sink__payload$24[62] ),
    .A2(net2292),
    .B1(net2174),
    .Y(_17523_));
 sky130_fd_sc_hd__a21oi_1 _39240_ (.A1(_13756_),
    .A2(net2292),
    .B1(_17523_),
    .Y(_04910_));
 sky130_fd_sc_hd__o21ai_0 _39241_ (.A1(\inst$top.soc.cpu.sink__payload$24[63] ),
    .A2(net2291),
    .B1(net2174),
    .Y(_17524_));
 sky130_fd_sc_hd__a21oi_1 _39242_ (.A1(_13811_),
    .A2(net2291),
    .B1(_17524_),
    .Y(_04911_));
 sky130_fd_sc_hd__o21ai_0 _39243_ (.A1(\inst$top.soc.cpu.sink__payload$24[64] ),
    .A2(net2291),
    .B1(net2174),
    .Y(_17525_));
 sky130_fd_sc_hd__nor2_1 _39244_ (.A(net1924),
    .B(_13909_),
    .Y(_17526_));
 sky130_fd_sc_hd__nor2_1 _39245_ (.A(_17525_),
    .B(_17526_),
    .Y(_04912_));
 sky130_fd_sc_hd__o21ai_0 _39246_ (.A1(\inst$top.soc.cpu.sink__payload$24[65] ),
    .A2(net2292),
    .B1(net2173),
    .Y(_17527_));
 sky130_fd_sc_hd__nor2_1 _39247_ (.A(net1925),
    .B(_13958_),
    .Y(_17528_));
 sky130_fd_sc_hd__nor2_1 _39248_ (.A(_17527_),
    .B(_17528_),
    .Y(_04913_));
 sky130_fd_sc_hd__o21ai_0 _39249_ (.A1(\inst$top.soc.cpu.sink__payload$24[66] ),
    .A2(net2280),
    .B1(net2157),
    .Y(_17529_));
 sky130_fd_sc_hd__nor2_1 _39250_ (.A(net1918),
    .B(_14008_),
    .Y(_17530_));
 sky130_fd_sc_hd__nor2_1 _39251_ (.A(_17529_),
    .B(_17530_),
    .Y(_04914_));
 sky130_fd_sc_hd__o21ai_0 _39252_ (.A1(\inst$top.soc.cpu.sink__payload$24[67] ),
    .A2(net2275),
    .B1(net2151),
    .Y(_17531_));
 sky130_fd_sc_hd__a21oi_1 _39253_ (.A1(_14021_),
    .A2(net2274),
    .B1(_17531_),
    .Y(_04915_));
 sky130_fd_sc_hd__o21ai_0 _39255_ (.A1(\inst$top.soc.cpu.sink__payload$24[68] ),
    .A2(net2274),
    .B1(net2153),
    .Y(_17533_));
 sky130_fd_sc_hd__a21oi_1 _39256_ (.A1(_14075_),
    .A2(net2274),
    .B1(_17533_),
    .Y(_04916_));
 sky130_fd_sc_hd__o21ai_0 _39257_ (.A1(\inst$top.soc.cpu.sink__payload$24[69] ),
    .A2(net2288),
    .B1(net2175),
    .Y(_17534_));
 sky130_fd_sc_hd__nor2_1 _39258_ (.A(net1925),
    .B(_14173_),
    .Y(_17535_));
 sky130_fd_sc_hd__nor2_1 _39259_ (.A(_17534_),
    .B(_17535_),
    .Y(_04917_));
 sky130_fd_sc_hd__nor2_1 _39260_ (.A(\inst$top.soc.cpu.sink__payload$18[6] ),
    .B(net1887),
    .Y(_17536_));
 sky130_fd_sc_hd__o21ai_0 _39261_ (.A1(\inst$top.soc.cpu.sink__payload$24[6] ),
    .A2(net2226),
    .B1(net2042),
    .Y(_17537_));
 sky130_fd_sc_hd__nor2_1 _39262_ (.A(_17536_),
    .B(_17537_),
    .Y(_04918_));
 sky130_fd_sc_hd__o21ai_0 _39263_ (.A1(\inst$top.soc.cpu.sink__payload$24[70] ),
    .A2(net2292),
    .B1(net2173),
    .Y(_17538_));
 sky130_fd_sc_hd__nor2_1 _39264_ (.A(net1924),
    .B(_14236_),
    .Y(_17539_));
 sky130_fd_sc_hd__nor2_1 _39265_ (.A(_17538_),
    .B(_17539_),
    .Y(_04919_));
 sky130_fd_sc_hd__o21ai_0 _39266_ (.A1(\inst$top.soc.cpu.sink__payload$24[71] ),
    .A2(net2274),
    .B1(net2156),
    .Y(_17540_));
 sky130_fd_sc_hd__a21oi_1 _39267_ (.A1(_14277_),
    .A2(net2274),
    .B1(_17540_),
    .Y(_04920_));
 sky130_fd_sc_hd__o21ai_0 _39269_ (.A1(\inst$top.soc.cpu.sink__payload$24[72] ),
    .A2(net2274),
    .B1(net2155),
    .Y(_17542_));
 sky130_fd_sc_hd__a21oi_1 _39270_ (.A1(_14359_),
    .A2(net2275),
    .B1(_17542_),
    .Y(_04921_));
 sky130_fd_sc_hd__o21ai_0 _39271_ (.A1(\inst$top.soc.cpu.d.sink__payload$16.load ),
    .A2(net2275),
    .B1(net2151),
    .Y(_17543_));
 sky130_fd_sc_hd__a21oi_1 _39272_ (.A1(_20187_),
    .A2(net2275),
    .B1(_17543_),
    .Y(_04922_));
 sky130_fd_sc_hd__o21ai_0 _39273_ (.A1(\inst$top.soc.cpu.sink__payload$24[74] ),
    .A2(net2266),
    .B1(net2130),
    .Y(_17544_));
 sky130_fd_sc_hd__a21oi_1 _39274_ (.A1(_15013_),
    .A2(net2266),
    .B1(_17544_),
    .Y(_04923_));
 sky130_fd_sc_hd__o21ai_0 _39275_ (.A1(\inst$top.soc.cpu.sink__payload$24[75] ),
    .A2(net2269),
    .B1(net2130),
    .Y(_17545_));
 sky130_fd_sc_hd__a21oi_1 _39276_ (.A1(_15049_),
    .A2(net2269),
    .B1(_17545_),
    .Y(_04924_));
 sky130_fd_sc_hd__o21ai_0 _39277_ (.A1(\inst$top.soc.cpu.sink__payload$24[76] ),
    .A2(net2267),
    .B1(net2127),
    .Y(_17546_));
 sky130_fd_sc_hd__a21oi_1 _39278_ (.A1(_15085_),
    .A2(net2267),
    .B1(_17546_),
    .Y(_04925_));
 sky130_fd_sc_hd__o21ai_0 _39280_ (.A1(\inst$top.soc.cpu.sink__payload$24[77] ),
    .A2(net2265),
    .B1(net2130),
    .Y(_17548_));
 sky130_fd_sc_hd__a21oi_1 _39281_ (.A1(_15095_),
    .A2(net2265),
    .B1(_17548_),
    .Y(_04926_));
 sky130_fd_sc_hd__o21ai_0 _39282_ (.A1(\inst$top.soc.cpu.sink__payload$24[78] ),
    .A2(net2269),
    .B1(net2136),
    .Y(_17549_));
 sky130_fd_sc_hd__a21oi_1 _39283_ (.A1(_15098_),
    .A2(net2269),
    .B1(_17549_),
    .Y(_04927_));
 sky130_fd_sc_hd__o21ai_0 _39284_ (.A1(\inst$top.soc.cpu.sink__payload$24[79] ),
    .A2(net2269),
    .B1(net2136),
    .Y(_17550_));
 sky130_fd_sc_hd__a21oi_1 _39285_ (.A1(_15101_),
    .A2(net2268),
    .B1(_17550_),
    .Y(_04928_));
 sky130_fd_sc_hd__nor2_1 _39286_ (.A(\inst$top.soc.cpu.sink__payload$18[7] ),
    .B(net1883),
    .Y(_17551_));
 sky130_fd_sc_hd__o21ai_0 _39287_ (.A1(\inst$top.soc.cpu.sink__payload$24[7] ),
    .A2(net2219),
    .B1(net2032),
    .Y(_17552_));
 sky130_fd_sc_hd__nor2_1 _39288_ (.A(_17551_),
    .B(_17552_),
    .Y(_04929_));
 sky130_fd_sc_hd__o21ai_0 _39290_ (.A1(\inst$top.soc.cpu.sink__payload$24[80] ),
    .A2(net2273),
    .B1(net2138),
    .Y(_17554_));
 sky130_fd_sc_hd__a21oi_1 _39291_ (.A1(_15104_),
    .A2(net2273),
    .B1(_17554_),
    .Y(_04930_));
 sky130_fd_sc_hd__o21ai_0 _39292_ (.A1(\inst$top.soc.cpu.sink__payload$24[81] ),
    .A2(net2269),
    .B1(net2136),
    .Y(_17555_));
 sky130_fd_sc_hd__a21oi_1 _39293_ (.A1(_15107_),
    .A2(net2268),
    .B1(_17555_),
    .Y(_04931_));
 sky130_fd_sc_hd__o21ai_0 _39295_ (.A1(\inst$top.soc.cpu.sink__payload$24[82] ),
    .A2(net2265),
    .B1(net2144),
    .Y(_17557_));
 sky130_fd_sc_hd__a21oi_1 _39296_ (.A1(_15110_),
    .A2(net2266),
    .B1(_17557_),
    .Y(_04932_));
 sky130_fd_sc_hd__o21ai_0 _39297_ (.A1(\inst$top.soc.cpu.sink__payload$24[83] ),
    .A2(net2273),
    .B1(net2136),
    .Y(_17558_));
 sky130_fd_sc_hd__a21oi_1 _39298_ (.A1(_15113_),
    .A2(net2273),
    .B1(_17558_),
    .Y(_04933_));
 sky130_fd_sc_hd__o21ai_0 _39299_ (.A1(\inst$top.soc.cpu.sink__payload$24[84] ),
    .A2(net2266),
    .B1(net2130),
    .Y(_17559_));
 sky130_fd_sc_hd__a21oi_1 _39300_ (.A1(_15016_),
    .A2(net2266),
    .B1(_17559_),
    .Y(_04934_));
 sky130_fd_sc_hd__o21ai_0 _39301_ (.A1(\inst$top.soc.cpu.sink__payload$24[85] ),
    .A2(net2270),
    .B1(net2136),
    .Y(_17560_));
 sky130_fd_sc_hd__a21oi_1 _39302_ (.A1(_15019_),
    .A2(net2270),
    .B1(_17560_),
    .Y(_04935_));
 sky130_fd_sc_hd__o21ai_0 _39303_ (.A1(\inst$top.soc.cpu.sink__payload$24[86] ),
    .A2(net2270),
    .B1(net2130),
    .Y(_17561_));
 sky130_fd_sc_hd__a21oi_1 _39304_ (.A1(_15022_),
    .A2(net2269),
    .B1(_17561_),
    .Y(_04936_));
 sky130_fd_sc_hd__o21ai_0 _39306_ (.A1(\inst$top.soc.cpu.sink__payload$24[87] ),
    .A2(net2272),
    .B1(net2138),
    .Y(_17563_));
 sky130_fd_sc_hd__a21oi_1 _39307_ (.A1(_15026_),
    .A2(net2272),
    .B1(_17563_),
    .Y(_04937_));
 sky130_fd_sc_hd__o21ai_0 _39308_ (.A1(\inst$top.soc.cpu.sink__payload$24[88] ),
    .A2(net2272),
    .B1(net2138),
    .Y(_17564_));
 sky130_fd_sc_hd__a21oi_1 _39309_ (.A1(_15029_),
    .A2(net2272),
    .B1(_17564_),
    .Y(_04938_));
 sky130_fd_sc_hd__o21ai_0 _39310_ (.A1(\inst$top.soc.cpu.sink__payload$24[89] ),
    .A2(net2268),
    .B1(net2136),
    .Y(_17565_));
 sky130_fd_sc_hd__a21oi_1 _39311_ (.A1(_15032_),
    .A2(net2268),
    .B1(_17565_),
    .Y(_04939_));
 sky130_fd_sc_hd__nor2_1 _39312_ (.A(\inst$top.soc.cpu.sink__payload$18[8] ),
    .B(net1896),
    .Y(_17566_));
 sky130_fd_sc_hd__o21ai_0 _39313_ (.A1(\inst$top.soc.cpu.sink__payload$24[8] ),
    .A2(net2228),
    .B1(net2044),
    .Y(_17567_));
 sky130_fd_sc_hd__nor2_1 _39314_ (.A(_17566_),
    .B(_17567_),
    .Y(_04940_));
 sky130_fd_sc_hd__o21ai_0 _39317_ (.A1(\inst$top.soc.cpu.sink__payload$24[90] ),
    .A2(net2271),
    .B1(net2139),
    .Y(_17570_));
 sky130_fd_sc_hd__a21oi_1 _39318_ (.A1(_15035_),
    .A2(net2271),
    .B1(_17570_),
    .Y(_04941_));
 sky130_fd_sc_hd__o21ai_0 _39319_ (.A1(\inst$top.soc.cpu.sink__payload$24[91] ),
    .A2(net2288),
    .B1(net2138),
    .Y(_17571_));
 sky130_fd_sc_hd__a21oi_1 _39320_ (.A1(_15039_),
    .A2(net2288),
    .B1(_17571_),
    .Y(_04942_));
 sky130_fd_sc_hd__o21ai_0 _39321_ (.A1(\inst$top.soc.cpu.sink__payload$24[92] ),
    .A2(net2268),
    .B1(net2137),
    .Y(_17572_));
 sky130_fd_sc_hd__a21oi_1 _39322_ (.A1(_15042_),
    .A2(net2268),
    .B1(_17572_),
    .Y(_04943_));
 sky130_fd_sc_hd__o21ai_0 _39323_ (.A1(\inst$top.soc.cpu.sink__payload$24[93] ),
    .A2(net2288),
    .B1(net2138),
    .Y(_17573_));
 sky130_fd_sc_hd__a21oi_1 _39324_ (.A1(_15046_),
    .A2(net2288),
    .B1(_17573_),
    .Y(_04944_));
 sky130_fd_sc_hd__o21ai_0 _39325_ (.A1(\inst$top.soc.cpu.sink__payload$24[94] ),
    .A2(net2273),
    .B1(net2137),
    .Y(_17574_));
 sky130_fd_sc_hd__a21oi_1 _39326_ (.A1(_15052_),
    .A2(net2273),
    .B1(_17574_),
    .Y(_04945_));
 sky130_fd_sc_hd__o21ai_0 _39327_ (.A1(\inst$top.soc.cpu.sink__payload$24[95] ),
    .A2(net2271),
    .B1(net2138),
    .Y(_17575_));
 sky130_fd_sc_hd__a21oi_1 _39328_ (.A1(_15055_),
    .A2(net2271),
    .B1(_17575_),
    .Y(_04946_));
 sky130_fd_sc_hd__o21ai_0 _39329_ (.A1(\inst$top.soc.cpu.sink__payload$24[96] ),
    .A2(net2271),
    .B1(net2138),
    .Y(_17576_));
 sky130_fd_sc_hd__a21oi_1 _39330_ (.A1(_15059_),
    .A2(net2271),
    .B1(_17576_),
    .Y(_04947_));
 sky130_fd_sc_hd__o21ai_0 _39331_ (.A1(\inst$top.soc.cpu.sink__payload$24[97] ),
    .A2(net2268),
    .B1(net2136),
    .Y(_17577_));
 sky130_fd_sc_hd__a21oi_1 _39332_ (.A1(_15062_),
    .A2(net2268),
    .B1(_17577_),
    .Y(_04948_));
 sky130_fd_sc_hd__o21ai_0 _39333_ (.A1(\inst$top.soc.cpu.sink__payload$24[98] ),
    .A2(net2271),
    .B1(net2138),
    .Y(_17578_));
 sky130_fd_sc_hd__a21oi_1 _39334_ (.A1(_15065_),
    .A2(net2271),
    .B1(_17578_),
    .Y(_04949_));
 sky130_fd_sc_hd__o21ai_0 _39335_ (.A1(\inst$top.soc.cpu.sink__payload$24[99] ),
    .A2(net2273),
    .B1(net2136),
    .Y(_17579_));
 sky130_fd_sc_hd__a21oi_1 _39336_ (.A1(_15068_),
    .A2(net2273),
    .B1(_17579_),
    .Y(_04950_));
 sky130_fd_sc_hd__nor2_1 _39337_ (.A(\inst$top.soc.cpu.sink__payload$18[9] ),
    .B(net1889),
    .Y(_17580_));
 sky130_fd_sc_hd__o21ai_0 _39338_ (.A1(\inst$top.soc.cpu.sink__payload$24[9] ),
    .A2(net2228),
    .B1(net2044),
    .Y(_17581_));
 sky130_fd_sc_hd__nor2_1 _39339_ (.A(_17580_),
    .B(_17581_),
    .Y(_04951_));
 sky130_fd_sc_hd__nor2_1 _39340_ (.A(\inst$top.soc.cpu.sink__payload$6[10] ),
    .B(net676),
    .Y(_17582_));
 sky130_fd_sc_hd__o21ai_1 _39342_ (.A1(\inst$top.soc.cpu.sink__payload[10] ),
    .A2(net630),
    .B1(net2067),
    .Y(_17584_));
 sky130_fd_sc_hd__nor2_4 _39343_ (.A(_17582_),
    .B(_17584_),
    .Y(_04952_));
 sky130_fd_sc_hd__nor2_1 _39344_ (.A(\inst$top.soc.cpu.sink__payload$6[11] ),
    .B(net669),
    .Y(_17585_));
 sky130_fd_sc_hd__o21ai_1 _39345_ (.A1(\inst$top.soc.cpu.sink__payload[11] ),
    .A2(net629),
    .B1(net2038),
    .Y(_17586_));
 sky130_fd_sc_hd__nor2_4 _39346_ (.A(_17585_),
    .B(_17586_),
    .Y(_04953_));
 sky130_fd_sc_hd__nor2_1 _39347_ (.A(\inst$top.soc.cpu.sink__payload$6[12] ),
    .B(net675),
    .Y(_17587_));
 sky130_fd_sc_hd__o21ai_1 _39349_ (.A1(\inst$top.soc.cpu.sink__payload[12] ),
    .A2(net629),
    .B1(net2039),
    .Y(_17589_));
 sky130_fd_sc_hd__nor2_4 _39350_ (.A(_17587_),
    .B(_17589_),
    .Y(_04954_));
 sky130_fd_sc_hd__nor2_1 _39351_ (.A(\inst$top.soc.cpu.sink__payload$6[13] ),
    .B(net676),
    .Y(_17590_));
 sky130_fd_sc_hd__o21ai_1 _39352_ (.A1(\inst$top.soc.cpu.sink__payload[13] ),
    .A2(net630),
    .B1(net2039),
    .Y(_17591_));
 sky130_fd_sc_hd__nor2_4 _39353_ (.A(_17590_),
    .B(_17591_),
    .Y(_04955_));
 sky130_fd_sc_hd__nor2_1 _39354_ (.A(\inst$top.soc.cpu.sink__payload$6[14] ),
    .B(net675),
    .Y(_17592_));
 sky130_fd_sc_hd__o21ai_1 _39355_ (.A1(\inst$top.soc.cpu.sink__payload[14] ),
    .A2(net627),
    .B1(net2039),
    .Y(_17593_));
 sky130_fd_sc_hd__nor2_4 _39356_ (.A(_17592_),
    .B(_17593_),
    .Y(_04956_));
 sky130_fd_sc_hd__nor2_1 _39357_ (.A(\inst$top.soc.cpu.sink__payload$6[15] ),
    .B(net675),
    .Y(_17594_));
 sky130_fd_sc_hd__o21ai_1 _39358_ (.A1(\inst$top.soc.cpu.sink__payload[15] ),
    .A2(net628),
    .B1(net2067),
    .Y(_17595_));
 sky130_fd_sc_hd__nor2_4 _39359_ (.A(_17594_),
    .B(_17595_),
    .Y(_04957_));
 sky130_fd_sc_hd__nor2_1 _39360_ (.A(\inst$top.soc.cpu.sink__payload$6[16] ),
    .B(net676),
    .Y(_17596_));
 sky130_fd_sc_hd__o21ai_1 _39361_ (.A1(\inst$top.soc.cpu.sink__payload[16] ),
    .A2(net627),
    .B1(net2039),
    .Y(_17597_));
 sky130_fd_sc_hd__nor2_4 _39362_ (.A(_17596_),
    .B(_17597_),
    .Y(_04958_));
 sky130_fd_sc_hd__nor2_1 _39363_ (.A(\inst$top.soc.cpu.sink__payload$6[17] ),
    .B(net676),
    .Y(_17598_));
 sky130_fd_sc_hd__o21ai_1 _39364_ (.A1(\inst$top.soc.cpu.sink__payload[17] ),
    .A2(net627),
    .B1(net2039),
    .Y(_17599_));
 sky130_fd_sc_hd__nor2_4 _39365_ (.A(_17598_),
    .B(_17599_),
    .Y(_04959_));
 sky130_fd_sc_hd__nor2_1 _39366_ (.A(\inst$top.soc.cpu.sink__payload$6[18] ),
    .B(net670),
    .Y(_17600_));
 sky130_fd_sc_hd__o21ai_1 _39367_ (.A1(\inst$top.soc.cpu.sink__payload[18] ),
    .A2(net622),
    .B1(net2037),
    .Y(_17601_));
 sky130_fd_sc_hd__nor2_4 _39368_ (.A(_17600_),
    .B(_17601_),
    .Y(_04960_));
 sky130_fd_sc_hd__nor2_1 _39370_ (.A(\inst$top.soc.cpu.sink__payload$6[19] ),
    .B(net675),
    .Y(_17603_));
 sky130_fd_sc_hd__o21ai_1 _39371_ (.A1(\inst$top.soc.cpu.sink__payload[19] ),
    .A2(net631),
    .B1(net2039),
    .Y(_17604_));
 sky130_fd_sc_hd__nor2_4 _39372_ (.A(_17603_),
    .B(_17604_),
    .Y(_04961_));
 sky130_fd_sc_hd__nor2_1 _39373_ (.A(\inst$top.soc.cpu.sink__payload$6[20] ),
    .B(net670),
    .Y(_17605_));
 sky130_fd_sc_hd__o21ai_1 _39375_ (.A1(\inst$top.soc.cpu.sink__payload[20] ),
    .A2(net622),
    .B1(net2037),
    .Y(_17607_));
 sky130_fd_sc_hd__nor2_4 _39376_ (.A(_17605_),
    .B(_17607_),
    .Y(_04962_));
 sky130_fd_sc_hd__nor2_1 _39377_ (.A(\inst$top.soc.cpu.sink__payload$6[21] ),
    .B(net670),
    .Y(_17608_));
 sky130_fd_sc_hd__o21ai_1 _39378_ (.A1(\inst$top.soc.cpu.sink__payload[21] ),
    .A2(net626),
    .B1(net2037),
    .Y(_17609_));
 sky130_fd_sc_hd__nor2_4 _39379_ (.A(_17608_),
    .B(_17609_),
    .Y(_04963_));
 sky130_fd_sc_hd__nor2_1 _39380_ (.A(\inst$top.soc.cpu.sink__payload$6[22] ),
    .B(net677),
    .Y(_17610_));
 sky130_fd_sc_hd__o21ai_0 _39382_ (.A1(\inst$top.soc.cpu.sink__payload[22] ),
    .A2(net636),
    .B1(net2067),
    .Y(_17612_));
 sky130_fd_sc_hd__nor2_2 _39383_ (.A(_17610_),
    .B(_17612_),
    .Y(_04964_));
 sky130_fd_sc_hd__nor2_1 _39384_ (.A(\inst$top.soc.cpu.sink__payload$6[23] ),
    .B(net677),
    .Y(_17613_));
 sky130_fd_sc_hd__o21ai_0 _39385_ (.A1(\inst$top.soc.cpu.sink__payload[23] ),
    .A2(net636),
    .B1(net2067),
    .Y(_17614_));
 sky130_fd_sc_hd__nor2_2 _39386_ (.A(_17613_),
    .B(_17614_),
    .Y(_04965_));
 sky130_fd_sc_hd__nor2_1 _39387_ (.A(\inst$top.soc.cpu.sink__payload$6[24] ),
    .B(net677),
    .Y(_17615_));
 sky130_fd_sc_hd__o21ai_0 _39388_ (.A1(\inst$top.soc.cpu.sink__payload[24] ),
    .A2(net636),
    .B1(net2050),
    .Y(_17616_));
 sky130_fd_sc_hd__nor2_2 _39389_ (.A(_17615_),
    .B(_17616_),
    .Y(_04966_));
 sky130_fd_sc_hd__nor2_1 _39390_ (.A(\inst$top.soc.cpu.sink__payload$6[25] ),
    .B(net676),
    .Y(_17617_));
 sky130_fd_sc_hd__o21ai_0 _39391_ (.A1(\inst$top.soc.cpu.sink__payload[25] ),
    .A2(net628),
    .B1(net2067),
    .Y(_17618_));
 sky130_fd_sc_hd__nor2_2 _39392_ (.A(_17617_),
    .B(_17618_),
    .Y(_04967_));
 sky130_fd_sc_hd__nor2_1 _39393_ (.A(\inst$top.soc.cpu.sink__payload$6[26] ),
    .B(net682),
    .Y(_17619_));
 sky130_fd_sc_hd__o21ai_0 _39394_ (.A1(\inst$top.soc.cpu.sink__payload[26] ),
    .A2(net638),
    .B1(net2073),
    .Y(_17620_));
 sky130_fd_sc_hd__nor2_2 _39395_ (.A(_17619_),
    .B(_17620_),
    .Y(_04968_));
 sky130_fd_sc_hd__nor2_1 _39396_ (.A(\inst$top.soc.cpu.sink__payload$6[27] ),
    .B(net682),
    .Y(_17621_));
 sky130_fd_sc_hd__o21ai_0 _39397_ (.A1(\inst$top.soc.cpu.sink__payload[27] ),
    .A2(net638),
    .B1(net2073),
    .Y(_17622_));
 sky130_fd_sc_hd__nor2_2 _39398_ (.A(_17621_),
    .B(_17622_),
    .Y(_04969_));
 sky130_fd_sc_hd__nor2_1 _39399_ (.A(\inst$top.soc.cpu.sink__payload$6[28] ),
    .B(net682),
    .Y(_17623_));
 sky130_fd_sc_hd__o21ai_0 _39400_ (.A1(\inst$top.soc.cpu.sink__payload[28] ),
    .A2(net636),
    .B1(net2066),
    .Y(_17624_));
 sky130_fd_sc_hd__nor2_2 _39401_ (.A(_17623_),
    .B(_17624_),
    .Y(_04970_));
 sky130_fd_sc_hd__nor2_1 _39403_ (.A(\inst$top.soc.cpu.sink__payload$6[29] ),
    .B(net677),
    .Y(_17626_));
 sky130_fd_sc_hd__o21ai_0 _39404_ (.A1(\inst$top.soc.cpu.sink__payload[29] ),
    .A2(net635),
    .B1(net2066),
    .Y(_17627_));
 sky130_fd_sc_hd__nor2_2 _39405_ (.A(_17626_),
    .B(_17627_),
    .Y(_04971_));
 sky130_fd_sc_hd__nor2_1 _39406_ (.A(\inst$top.soc.cpu.sink__payload$6[2] ),
    .B(net667),
    .Y(_17628_));
 sky130_fd_sc_hd__o21ai_0 _39408_ (.A1(\inst$top.soc.cpu.sink__payload[2] ),
    .A2(net624),
    .B1(net2030),
    .Y(_17630_));
 sky130_fd_sc_hd__nor2_2 _39409_ (.A(_17628_),
    .B(_17630_),
    .Y(_04972_));
 sky130_fd_sc_hd__nor2_1 _39410_ (.A(\inst$top.soc.cpu.sink__payload$6[30] ),
    .B(net677),
    .Y(_17631_));
 sky130_fd_sc_hd__o21ai_0 _39411_ (.A1(\inst$top.soc.cpu.sink__payload[30] ),
    .A2(net635),
    .B1(net2050),
    .Y(_17632_));
 sky130_fd_sc_hd__nor2_2 _39412_ (.A(_17631_),
    .B(_17632_),
    .Y(_04973_));
 sky130_fd_sc_hd__nor2_1 _39413_ (.A(\inst$top.soc.cpu.sink__payload$6[31] ),
    .B(net670),
    .Y(_17633_));
 sky130_fd_sc_hd__o21ai_0 _39415_ (.A1(\inst$top.soc.cpu.sink__payload[31] ),
    .A2(net621),
    .B1(net2030),
    .Y(_17635_));
 sky130_fd_sc_hd__nor2_2 _39416_ (.A(_17633_),
    .B(_17635_),
    .Y(_04974_));
 sky130_fd_sc_hd__nor2_1 _39417_ (.A(\inst$top.soc.cpu.sink__payload$6[32] ),
    .B(net685),
    .Y(_17636_));
 sky130_fd_sc_hd__o21ai_0 _39418_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[0] ),
    .A2(net638),
    .B1(net2060),
    .Y(_17637_));
 sky130_fd_sc_hd__nor2_2 _39419_ (.A(_17636_),
    .B(_17637_),
    .Y(_04975_));
 sky130_fd_sc_hd__nor2_1 _39420_ (.A(\inst$top.soc.cpu.sink__payload$6[33] ),
    .B(net685),
    .Y(_17638_));
 sky130_fd_sc_hd__o21ai_0 _39421_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[1] ),
    .A2(net638),
    .B1(net2060),
    .Y(_17639_));
 sky130_fd_sc_hd__nor2_2 _39422_ (.A(_17638_),
    .B(_17639_),
    .Y(_04976_));
 sky130_fd_sc_hd__nor2_1 _39423_ (.A(\inst$top.soc.cpu.sink__payload$6[34] ),
    .B(net682),
    .Y(_17640_));
 sky130_fd_sc_hd__o21ai_0 _39424_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[2] ),
    .A2(net638),
    .B1(net2060),
    .Y(_17641_));
 sky130_fd_sc_hd__nor2_2 _39425_ (.A(_17640_),
    .B(_17641_),
    .Y(_04977_));
 sky130_fd_sc_hd__nor2_1 _39426_ (.A(\inst$top.soc.cpu.sink__payload$6[35] ),
    .B(net686),
    .Y(_17642_));
 sky130_fd_sc_hd__o21ai_0 _39427_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[3] ),
    .A2(net639),
    .B1(net2076),
    .Y(_17643_));
 sky130_fd_sc_hd__nor2_2 _39428_ (.A(_17642_),
    .B(_17643_),
    .Y(_04978_));
 sky130_fd_sc_hd__nor2_1 _39429_ (.A(\inst$top.soc.cpu.sink__payload$6[36] ),
    .B(net686),
    .Y(_17644_));
 sky130_fd_sc_hd__o21ai_0 _39430_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[4] ),
    .A2(net639),
    .B1(net2062),
    .Y(_17645_));
 sky130_fd_sc_hd__nor2_2 _39431_ (.A(_17644_),
    .B(_17645_),
    .Y(_04979_));
 sky130_fd_sc_hd__nor2_1 _39432_ (.A(\inst$top.soc.cpu.sink__payload$6[37] ),
    .B(net686),
    .Y(_17646_));
 sky130_fd_sc_hd__o21ai_0 _39433_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[5] ),
    .A2(net639),
    .B1(net2062),
    .Y(_17647_));
 sky130_fd_sc_hd__nor2_2 _39434_ (.A(_17646_),
    .B(_17647_),
    .Y(_04980_));
 sky130_fd_sc_hd__nor2_1 _39436_ (.A(\inst$top.soc.cpu.sink__payload$6[38] ),
    .B(net689),
    .Y(_17649_));
 sky130_fd_sc_hd__o21ai_0 _39437_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[6] ),
    .A2(net649),
    .B1(net2062),
    .Y(_17650_));
 sky130_fd_sc_hd__nor2_2 _39438_ (.A(_17649_),
    .B(_17650_),
    .Y(_04981_));
 sky130_fd_sc_hd__nor2_1 _39439_ (.A(\inst$top.soc.cpu.sink__payload$6[39] ),
    .B(net697),
    .Y(_17651_));
 sky130_fd_sc_hd__o21ai_0 _39441_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[7] ),
    .A2(net651),
    .B1(net2131),
    .Y(_17653_));
 sky130_fd_sc_hd__nor2_2 _39442_ (.A(_17651_),
    .B(_17653_),
    .Y(_04982_));
 sky130_fd_sc_hd__nor2_1 _39443_ (.A(\inst$top.soc.cpu.sink__payload$6[3] ),
    .B(net667),
    .Y(_17654_));
 sky130_fd_sc_hd__o21ai_0 _39444_ (.A1(\inst$top.soc.cpu.sink__payload[3] ),
    .A2(net623),
    .B1(net2029),
    .Y(_17655_));
 sky130_fd_sc_hd__nor2_2 _39445_ (.A(_17654_),
    .B(_17655_),
    .Y(_04983_));
 sky130_fd_sc_hd__nor2_1 _39446_ (.A(\inst$top.soc.cpu.sink__payload$6[40] ),
    .B(net697),
    .Y(_17656_));
 sky130_fd_sc_hd__o21ai_0 _39448_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[8] ),
    .A2(net651),
    .B1(net2130),
    .Y(_17658_));
 sky130_fd_sc_hd__nor2_2 _39449_ (.A(_17656_),
    .B(_17658_),
    .Y(_04984_));
 sky130_fd_sc_hd__nor2_1 _39450_ (.A(\inst$top.soc.cpu.sink__payload$6[41] ),
    .B(net695),
    .Y(_17659_));
 sky130_fd_sc_hd__o21ai_0 _39451_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[9] ),
    .A2(net651),
    .B1(net2143),
    .Y(_17660_));
 sky130_fd_sc_hd__nor2_2 _39452_ (.A(_17659_),
    .B(_17660_),
    .Y(_04985_));
 sky130_fd_sc_hd__nor2_1 _39453_ (.A(\inst$top.soc.cpu.sink__payload$6[42] ),
    .B(net695),
    .Y(_17661_));
 sky130_fd_sc_hd__o21ai_0 _39454_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[10] ),
    .A2(net649),
    .B1(net2128),
    .Y(_17662_));
 sky130_fd_sc_hd__nor2_2 _39455_ (.A(_17661_),
    .B(_17662_),
    .Y(_04986_));
 sky130_fd_sc_hd__nor2_1 _39456_ (.A(\inst$top.soc.cpu.sink__payload$6[43] ),
    .B(net697),
    .Y(_17663_));
 sky130_fd_sc_hd__o21ai_0 _39457_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[11] ),
    .A2(net651),
    .B1(net2144),
    .Y(_17664_));
 sky130_fd_sc_hd__nor2_2 _39458_ (.A(_17663_),
    .B(_17664_),
    .Y(_04987_));
 sky130_fd_sc_hd__nor2_1 _39459_ (.A(\inst$top.soc.cpu.sink__payload$6[44] ),
    .B(net695),
    .Y(_17665_));
 sky130_fd_sc_hd__o21ai_0 _39460_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[12] ),
    .A2(net649),
    .B1(net2128),
    .Y(_17666_));
 sky130_fd_sc_hd__nor2_2 _39461_ (.A(_17665_),
    .B(_17666_),
    .Y(_04988_));
 sky130_fd_sc_hd__nor2_1 _39462_ (.A(\inst$top.soc.cpu.sink__payload$6[45] ),
    .B(net695),
    .Y(_17667_));
 sky130_fd_sc_hd__o21ai_0 _39463_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[13] ),
    .A2(net649),
    .B1(net2127),
    .Y(_17668_));
 sky130_fd_sc_hd__nor2_2 _39464_ (.A(_17667_),
    .B(_17668_),
    .Y(_04989_));
 sky130_fd_sc_hd__nor2_1 _39465_ (.A(net2820),
    .B(net686),
    .Y(_17669_));
 sky130_fd_sc_hd__o21ai_0 _39466_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[14] ),
    .A2(net649),
    .B1(net2063),
    .Y(_17670_));
 sky130_fd_sc_hd__nor2_2 _39467_ (.A(_17669_),
    .B(_17670_),
    .Y(_04990_));
 sky130_fd_sc_hd__nor2_1 _39469_ (.A(net2767),
    .B(net697),
    .Y(_17672_));
 sky130_fd_sc_hd__o21ai_0 _39470_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[15] ),
    .A2(net651),
    .B1(net2137),
    .Y(_17673_));
 sky130_fd_sc_hd__nor2_2 _39471_ (.A(_17672_),
    .B(_17673_),
    .Y(_04991_));
 sky130_fd_sc_hd__nor2_1 _39472_ (.A(net2724),
    .B(net708),
    .Y(_17674_));
 sky130_fd_sc_hd__o21ai_0 _39474_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[16] ),
    .A2(net656),
    .B1(net2139),
    .Y(_17676_));
 sky130_fd_sc_hd__nor2_2 _39475_ (.A(_17674_),
    .B(_17676_),
    .Y(_04992_));
 sky130_fd_sc_hd__nor2_1 _39476_ (.A(net2703),
    .B(net706),
    .Y(_17677_));
 sky130_fd_sc_hd__o21ai_0 _39477_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[17] ),
    .A2(net656),
    .B1(net2139),
    .Y(_17678_));
 sky130_fd_sc_hd__nor2_2 _39478_ (.A(_17677_),
    .B(_17678_),
    .Y(_04993_));
 sky130_fd_sc_hd__nor2_1 _39479_ (.A(\inst$top.soc.cpu.sink__payload$6[4] ),
    .B(net666),
    .Y(_17679_));
 sky130_fd_sc_hd__o21ai_0 _39481_ (.A1(\inst$top.soc.cpu.sink__payload[4] ),
    .A2(net624),
    .B1(net2029),
    .Y(_17681_));
 sky130_fd_sc_hd__nor2_2 _39482_ (.A(_17679_),
    .B(_17681_),
    .Y(_04994_));
 sky130_fd_sc_hd__nor2_1 _39483_ (.A(net2696),
    .B(net697),
    .Y(_17682_));
 sky130_fd_sc_hd__o21ai_0 _39484_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[18] ),
    .A2(net651),
    .B1(net2129),
    .Y(_17683_));
 sky130_fd_sc_hd__nor2_2 _39485_ (.A(_17682_),
    .B(_17683_),
    .Y(_04995_));
 sky130_fd_sc_hd__nor2_1 _39486_ (.A(net2690),
    .B(net697),
    .Y(_17684_));
 sky130_fd_sc_hd__o21ai_0 _39487_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[19] ),
    .A2(net651),
    .B1(net2136),
    .Y(_17685_));
 sky130_fd_sc_hd__nor2_2 _39488_ (.A(_17684_),
    .B(_17685_),
    .Y(_04996_));
 sky130_fd_sc_hd__nor2_1 _39489_ (.A(net2686),
    .B(net697),
    .Y(_17686_));
 sky130_fd_sc_hd__o21ai_0 _39490_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[20] ),
    .A2(net651),
    .B1(net2129),
    .Y(_17687_));
 sky130_fd_sc_hd__nor2_2 _39491_ (.A(_17686_),
    .B(_17687_),
    .Y(_04997_));
 sky130_fd_sc_hd__nor2_1 _39492_ (.A(net2620),
    .B(net697),
    .Y(_17688_));
 sky130_fd_sc_hd__o21ai_0 _39493_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[21] ),
    .A2(net651),
    .B1(net2137),
    .Y(_17689_));
 sky130_fd_sc_hd__nor2_2 _39494_ (.A(_17688_),
    .B(_17689_),
    .Y(_04998_));
 sky130_fd_sc_hd__nor2_1 _39495_ (.A(net2608),
    .B(net708),
    .Y(_17690_));
 sky130_fd_sc_hd__o21ai_0 _39496_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[22] ),
    .A2(net656),
    .B1(net2139),
    .Y(_17691_));
 sky130_fd_sc_hd__nor2_2 _39497_ (.A(_17690_),
    .B(_17691_),
    .Y(_04999_));
 sky130_fd_sc_hd__nor2_1 _39498_ (.A(net2597),
    .B(net689),
    .Y(_17692_));
 sky130_fd_sc_hd__o21ai_0 _39499_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[23] ),
    .A2(net649),
    .B1(net2127),
    .Y(_17693_));
 sky130_fd_sc_hd__nor2_2 _39500_ (.A(_17692_),
    .B(_17693_),
    .Y(_05000_));
 sky130_fd_sc_hd__nor2_1 _39502_ (.A(net2590),
    .B(net685),
    .Y(_17695_));
 sky130_fd_sc_hd__o21ai_0 _39503_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[24] ),
    .A2(net638),
    .B1(net2060),
    .Y(_17696_));
 sky130_fd_sc_hd__nor2_2 _39504_ (.A(_17695_),
    .B(_17696_),
    .Y(_05001_));
 sky130_fd_sc_hd__nor2_1 _39505_ (.A(\inst$top.soc.cpu.sink__payload$6[57] ),
    .B(net686),
    .Y(_17697_));
 sky130_fd_sc_hd__o21ai_0 _39507_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[25] ),
    .A2(net639),
    .B1(net2062),
    .Y(_17699_));
 sky130_fd_sc_hd__nor2_2 _39508_ (.A(_17697_),
    .B(_17699_),
    .Y(_05002_));
 sky130_fd_sc_hd__nor2_1 _39509_ (.A(\inst$top.soc.cpu.sink__payload$6[58] ),
    .B(net686),
    .Y(_17700_));
 sky130_fd_sc_hd__o21ai_0 _39510_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[26] ),
    .A2(net639),
    .B1(net2062),
    .Y(_17701_));
 sky130_fd_sc_hd__nor2_2 _39511_ (.A(_17700_),
    .B(_17701_),
    .Y(_05003_));
 sky130_fd_sc_hd__nor2_1 _39512_ (.A(\inst$top.soc.cpu.sink__payload$6[59] ),
    .B(net685),
    .Y(_17702_));
 sky130_fd_sc_hd__o21ai_0 _39514_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[27] ),
    .A2(net640),
    .B1(net2060),
    .Y(_17704_));
 sky130_fd_sc_hd__nor2_2 _39515_ (.A(_17702_),
    .B(_17704_),
    .Y(_05004_));
 sky130_fd_sc_hd__nor2_1 _39516_ (.A(\inst$top.soc.cpu.sink__payload$6[5] ),
    .B(net669),
    .Y(_17705_));
 sky130_fd_sc_hd__o21ai_0 _39517_ (.A1(\inst$top.soc.cpu.sink__payload[5] ),
    .A2(net625),
    .B1(net2038),
    .Y(_17706_));
 sky130_fd_sc_hd__nor2_2 _39518_ (.A(_17705_),
    .B(_17706_),
    .Y(_05005_));
 sky130_fd_sc_hd__nor2_1 _39519_ (.A(\inst$top.soc.cpu.sink__payload$6[60] ),
    .B(net686),
    .Y(_17707_));
 sky130_fd_sc_hd__o21ai_0 _39520_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[28] ),
    .A2(net640),
    .B1(net2062),
    .Y(_17708_));
 sky130_fd_sc_hd__nor2_2 _39521_ (.A(_17707_),
    .B(_17708_),
    .Y(_05006_));
 sky130_fd_sc_hd__nor2_1 _39522_ (.A(\inst$top.soc.cpu.sink__payload$6[61] ),
    .B(net689),
    .Y(_17709_));
 sky130_fd_sc_hd__o21ai_0 _39523_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[29] ),
    .A2(net639),
    .B1(net2063),
    .Y(_17710_));
 sky130_fd_sc_hd__nor2_2 _39524_ (.A(_17709_),
    .B(_17710_),
    .Y(_05007_));
 sky130_fd_sc_hd__nor2_1 _39525_ (.A(\inst$top.soc.cpu.sink__payload$6[62] ),
    .B(net686),
    .Y(_17711_));
 sky130_fd_sc_hd__o21ai_0 _39526_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[30] ),
    .A2(net640),
    .B1(net2062),
    .Y(_17712_));
 sky130_fd_sc_hd__nor2_2 _39527_ (.A(_17711_),
    .B(_17712_),
    .Y(_05008_));
 sky130_fd_sc_hd__nor2_1 _39528_ (.A(\inst$top.soc.cpu.sink__payload$6[63] ),
    .B(net689),
    .Y(_17713_));
 sky130_fd_sc_hd__o21ai_0 _39529_ (.A1(\inst$top.soc.cpu.fetch.ibus_rdata[31] ),
    .A2(net649),
    .B1(net2077),
    .Y(_17714_));
 sky130_fd_sc_hd__nor2_2 _39530_ (.A(_17713_),
    .B(_17714_),
    .Y(_05009_));
 sky130_fd_sc_hd__nor2_1 _39531_ (.A(\inst$top.soc.cpu.sink__payload$6[6] ),
    .B(net668),
    .Y(_17715_));
 sky130_fd_sc_hd__o21ai_0 _39532_ (.A1(\inst$top.soc.cpu.sink__payload[6] ),
    .A2(net625),
    .B1(net2038),
    .Y(_17716_));
 sky130_fd_sc_hd__nor2_2 _39533_ (.A(_17715_),
    .B(_17716_),
    .Y(_05010_));
 sky130_fd_sc_hd__nor2_1 _39534_ (.A(\inst$top.soc.cpu.sink__payload$6[7] ),
    .B(net668),
    .Y(_17717_));
 sky130_fd_sc_hd__o21ai_0 _39535_ (.A1(\inst$top.soc.cpu.sink__payload[7] ),
    .A2(net625),
    .B1(net2038),
    .Y(_17718_));
 sky130_fd_sc_hd__nor2_2 _39536_ (.A(_17717_),
    .B(_17718_),
    .Y(_05011_));
 sky130_fd_sc_hd__nor2_1 _39537_ (.A(\inst$top.soc.cpu.sink__payload$6[8] ),
    .B(net675),
    .Y(_17719_));
 sky130_fd_sc_hd__o21ai_0 _39539_ (.A1(\inst$top.soc.cpu.sink__payload[8] ),
    .A2(net630),
    .B1(net2040),
    .Y(_17721_));
 sky130_fd_sc_hd__nor2_2 _39540_ (.A(_17719_),
    .B(_17721_),
    .Y(_05012_));
 sky130_fd_sc_hd__nor2_1 _39541_ (.A(\inst$top.soc.cpu.sink__payload$6[9] ),
    .B(net675),
    .Y(_17722_));
 sky130_fd_sc_hd__o21ai_0 _39542_ (.A1(\inst$top.soc.cpu.sink__payload[9] ),
    .A2(net630),
    .B1(net2040),
    .Y(_17723_));
 sky130_fd_sc_hd__nor2_2 _39543_ (.A(_17722_),
    .B(_17723_),
    .Y(_05013_));
 sky130_fd_sc_hd__nand2_1 _39545_ (.A(net631),
    .B(\inst$top.soc.cpu.sink__payload[10] ),
    .Y(_17725_));
 sky130_fd_sc_hd__nand3_1 _39547_ (.A(_17725_),
    .B(_12673_),
    .C(net2041),
    .Y(_05014_));
 sky130_fd_sc_hd__nand2_1 _39548_ (.A(net632),
    .B(\inst$top.soc.cpu.sink__payload[11] ),
    .Y(_17727_));
 sky130_fd_sc_hd__nand3_1 _39549_ (.A(_17727_),
    .B(_12689_),
    .C(net2037),
    .Y(_05015_));
 sky130_fd_sc_hd__nand2_1 _39550_ (.A(net629),
    .B(\inst$top.soc.cpu.sink__payload[12] ),
    .Y(_17728_));
 sky130_fd_sc_hd__nand3_1 _39551_ (.A(_17728_),
    .B(_12001_),
    .C(net2039),
    .Y(_05016_));
 sky130_fd_sc_hd__nand2_1 _39552_ (.A(net631),
    .B(\inst$top.soc.cpu.sink__payload[13] ),
    .Y(_17729_));
 sky130_fd_sc_hd__nand3_1 _39553_ (.A(_17729_),
    .B(_12043_),
    .C(net2041),
    .Y(_05017_));
 sky130_fd_sc_hd__nand2_1 _39554_ (.A(net627),
    .B(\inst$top.soc.cpu.sink__payload[14] ),
    .Y(_17730_));
 sky130_fd_sc_hd__nand3_1 _39555_ (.A(_17730_),
    .B(_12064_),
    .C(net2039),
    .Y(_05018_));
 sky130_fd_sc_hd__nand2_1 _39556_ (.A(net628),
    .B(\inst$top.soc.cpu.sink__payload[15] ),
    .Y(_17731_));
 sky130_fd_sc_hd__nand3_1 _39557_ (.A(_17731_),
    .B(_12100_),
    .C(net2067),
    .Y(_05019_));
 sky130_fd_sc_hd__nand2_1 _39558_ (.A(net626),
    .B(\inst$top.soc.cpu.sink__payload[16] ),
    .Y(_17732_));
 sky130_fd_sc_hd__nand3_1 _39559_ (.A(_12126_),
    .B(net2027),
    .C(_17732_),
    .Y(_05020_));
 sky130_fd_sc_hd__nand2_1 _39560_ (.A(net627),
    .B(\inst$top.soc.cpu.sink__payload[17] ),
    .Y(_17733_));
 sky130_fd_sc_hd__nand3_1 _39561_ (.A(_17733_),
    .B(_12156_),
    .C(net2028),
    .Y(_05021_));
 sky130_fd_sc_hd__nand2_1 _39562_ (.A(net622),
    .B(\inst$top.soc.cpu.sink__payload[18] ),
    .Y(_17734_));
 sky130_fd_sc_hd__nand3_1 _39563_ (.A(_17734_),
    .B(_12178_),
    .C(net2037),
    .Y(_05022_));
 sky130_fd_sc_hd__nand2_1 _39564_ (.A(net626),
    .B(\inst$top.soc.cpu.sink__payload[19] ),
    .Y(_17735_));
 sky130_fd_sc_hd__nand3_1 _39565_ (.A(_12213_),
    .B(net2039),
    .C(_17735_),
    .Y(_05023_));
 sky130_fd_sc_hd__nand2_1 _39566_ (.A(net622),
    .B(\inst$top.soc.cpu.sink__payload[20] ),
    .Y(_17736_));
 sky130_fd_sc_hd__a21oi_2 _39567_ (.A1(_17736_),
    .A2(_12251_),
    .B1(net2943),
    .Y(_05024_));
 sky130_fd_sc_hd__nand2_1 _39568_ (.A(net626),
    .B(\inst$top.soc.cpu.sink__payload[21] ),
    .Y(_17737_));
 sky130_fd_sc_hd__a21oi_2 _39569_ (.A1(_17737_),
    .A2(_12273_),
    .B1(net2943),
    .Y(_05025_));
 sky130_fd_sc_hd__nand2_1 _39570_ (.A(net636),
    .B(\inst$top.soc.cpu.sink__payload[22] ),
    .Y(_17738_));
 sky130_fd_sc_hd__a21oi_2 _39571_ (.A1(_17738_),
    .A2(_12311_),
    .B1(net2945),
    .Y(_05026_));
 sky130_fd_sc_hd__nand2_1 _39572_ (.A(net636),
    .B(\inst$top.soc.cpu.sink__payload[23] ),
    .Y(_17739_));
 sky130_fd_sc_hd__a21oi_4 _39573_ (.A1(_12337_),
    .A2(_17739_),
    .B1(net2945),
    .Y(_05027_));
 sky130_fd_sc_hd__nand2_1 _39574_ (.A(net636),
    .B(\inst$top.soc.cpu.sink__payload[24] ),
    .Y(_17740_));
 sky130_fd_sc_hd__a21oi_4 _39575_ (.A1(_12361_),
    .A2(_17740_),
    .B1(net2945),
    .Y(_05028_));
 sky130_fd_sc_hd__nand2_1 _39576_ (.A(net627),
    .B(\inst$top.soc.cpu.sink__payload[25] ),
    .Y(_17741_));
 sky130_fd_sc_hd__a21oi_4 _39578_ (.A1(_12391_),
    .A2(_17741_),
    .B1(net2945),
    .Y(_05029_));
 sky130_fd_sc_hd__nand2_1 _39579_ (.A(net635),
    .B(\inst$top.soc.cpu.sink__payload[26] ),
    .Y(_17743_));
 sky130_fd_sc_hd__a21oi_4 _39580_ (.A1(_12427_),
    .A2(_17743_),
    .B1(net2951),
    .Y(_05030_));
 sky130_fd_sc_hd__nand2_1 _39581_ (.A(net638),
    .B(\inst$top.soc.cpu.sink__payload[27] ),
    .Y(_17744_));
 sky130_fd_sc_hd__a21oi_4 _39582_ (.A1(_12464_),
    .A2(_17744_),
    .B1(net2948),
    .Y(_05031_));
 sky130_fd_sc_hd__nand2_1 _39583_ (.A(net635),
    .B(\inst$top.soc.cpu.sink__payload[28] ),
    .Y(_17745_));
 sky130_fd_sc_hd__a21oi_4 _39584_ (.A1(_12488_),
    .A2(_17745_),
    .B1(net2946),
    .Y(_05032_));
 sky130_fd_sc_hd__nand2_1 _39585_ (.A(net635),
    .B(\inst$top.soc.cpu.sink__payload[29] ),
    .Y(_17746_));
 sky130_fd_sc_hd__a21oi_4 _39586_ (.A1(_12513_),
    .A2(_17746_),
    .B1(net2946),
    .Y(_05033_));
 sky130_fd_sc_hd__nand2_1 _39587_ (.A(net623),
    .B(\inst$top.soc.cpu.sink__payload[2] ),
    .Y(_17747_));
 sky130_fd_sc_hd__nand3_1 _39588_ (.A(_17747_),
    .B(_11952_),
    .C(net2030),
    .Y(_05034_));
 sky130_fd_sc_hd__nand2_1 _39589_ (.A(net635),
    .B(\inst$top.soc.cpu.sink__payload[30] ),
    .Y(_17748_));
 sky130_fd_sc_hd__a21oi_4 _39590_ (.A1(_12538_),
    .A2(_17748_),
    .B1(net2946),
    .Y(_05035_));
 sky130_fd_sc_hd__nand2_1 _39591_ (.A(net621),
    .B(\inst$top.soc.cpu.sink__payload[31] ),
    .Y(_17749_));
 sky130_fd_sc_hd__a21oi_4 _39592_ (.A1(_12567_),
    .A2(_17749_),
    .B1(net2938),
    .Y(_05036_));
 sky130_fd_sc_hd__nand2_1 _39593_ (.A(net623),
    .B(\inst$top.soc.cpu.sink__payload[3] ),
    .Y(_17750_));
 sky130_fd_sc_hd__nand3_1 _39594_ (.A(_17750_),
    .B(_12287_),
    .C(net2030),
    .Y(_05037_));
 sky130_fd_sc_hd__nand2_1 _39595_ (.A(net623),
    .B(\inst$top.soc.cpu.sink__payload[4] ),
    .Y(_17751_));
 sky130_fd_sc_hd__nand3_1 _39596_ (.A(_17751_),
    .B(_12585_),
    .C(net2030),
    .Y(_05038_));
 sky130_fd_sc_hd__nand2_1 _39597_ (.A(net625),
    .B(\inst$top.soc.cpu.sink__payload[5] ),
    .Y(_17752_));
 sky130_fd_sc_hd__nand3_1 _39598_ (.A(_12598_),
    .B(net2038),
    .C(_17752_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand2_1 _39599_ (.A(net625),
    .B(\inst$top.soc.cpu.sink__payload[6] ),
    .Y(_17753_));
 sky130_fd_sc_hd__nand3_1 _39600_ (.A(_12612_),
    .B(net2038),
    .C(_17753_),
    .Y(_05040_));
 sky130_fd_sc_hd__nand2_1 _39601_ (.A(net625),
    .B(\inst$top.soc.cpu.sink__payload[7] ),
    .Y(_17754_));
 sky130_fd_sc_hd__nand3_1 _39602_ (.A(_12626_),
    .B(net2037),
    .C(_17754_),
    .Y(_05041_));
 sky130_fd_sc_hd__nand2_1 _39603_ (.A(net629),
    .B(\inst$top.soc.cpu.sink__payload[8] ),
    .Y(_17755_));
 sky130_fd_sc_hd__nand3_1 _39604_ (.A(_12641_),
    .B(net2040),
    .C(_17755_),
    .Y(_05042_));
 sky130_fd_sc_hd__nand2_1 _39605_ (.A(net629),
    .B(\inst$top.soc.cpu.sink__payload[9] ),
    .Y(_17756_));
 sky130_fd_sc_hd__nand3_1 _39606_ (.A(_12655_),
    .B(net2040),
    .C(_17756_),
    .Y(_05043_));
 sky130_fd_sc_hd__o21ai_0 _39608_ (.A1(\inst$top.soc.cpu.x.source__valid ),
    .A2(net2267),
    .B1(net2145),
    .Y(_17758_));
 sky130_fd_sc_hd__a21oi_1 _39609_ (.A1(_20231_),
    .A2(net2267),
    .B1(_17758_),
    .Y(_05044_));
 sky130_fd_sc_hd__inv_1 _39610_ (.A(net2585),
    .Y(_17759_));
 sky130_fd_sc_hd__o21ai_0 _39611_ (.A1(\inst$top.soc.gpio_0._gpio.w_data ),
    .A2(_17759_),
    .B1(net2168),
    .Y(_17760_));
 sky130_fd_sc_hd__a21oi_1 _39612_ (.A1(_02871_),
    .A2(_17759_),
    .B1(_17760_),
    .Y(_05045_));
 sky130_fd_sc_hd__inv_1 _39613_ (.A(\inst$top.soc.gpio_0._gpio.w_data$16 ),
    .Y(_17761_));
 sky130_fd_sc_hd__o21ai_0 _39616_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__0._storage[1] ),
    .A2(net2585),
    .B1(net2168),
    .Y(_17764_));
 sky130_fd_sc_hd__a21oi_1 _39617_ (.A1(_17761_),
    .A2(net2585),
    .B1(_17764_),
    .Y(_05046_));
 sky130_fd_sc_hd__o21ai_0 _39618_ (.A1(\inst$top.soc.gpio_0._gpio.w_data$26 ),
    .A2(_17759_),
    .B1(net2167),
    .Y(_17765_));
 sky130_fd_sc_hd__a21oi_1 _39619_ (.A1(_02893_),
    .A2(_17759_),
    .B1(_17765_),
    .Y(_05047_));
 sky130_fd_sc_hd__inv_1 _39620_ (.A(\inst$top.soc.gpio_0._gpio.w_data$29 ),
    .Y(_17766_));
 sky130_fd_sc_hd__o21ai_0 _39621_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__1._storage[1] ),
    .A2(net2585),
    .B1(net2167),
    .Y(_17767_));
 sky130_fd_sc_hd__a21oi_1 _39622_ (.A1(_17766_),
    .A2(net2585),
    .B1(_17767_),
    .Y(_05048_));
 sky130_fd_sc_hd__inv_1 _39623_ (.A(\inst$top.soc.gpio_0._gpio.w_data$38 ),
    .Y(_17768_));
 sky130_fd_sc_hd__o21ai_0 _39624_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__2._storage[0] ),
    .A2(net2586),
    .B1(net2163),
    .Y(_17769_));
 sky130_fd_sc_hd__a21oi_1 _39625_ (.A1(_17768_),
    .A2(net2586),
    .B1(_17769_),
    .Y(_05049_));
 sky130_fd_sc_hd__inv_1 _39626_ (.A(\inst$top.soc.gpio_0._gpio.w_data$41 ),
    .Y(_17770_));
 sky130_fd_sc_hd__o21ai_0 _39627_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__2._storage[1] ),
    .A2(net2586),
    .B1(net2163),
    .Y(_17771_));
 sky130_fd_sc_hd__a21oi_1 _39628_ (.A1(_17770_),
    .A2(net2586),
    .B1(_17771_),
    .Y(_05050_));
 sky130_fd_sc_hd__o21ai_0 _39629_ (.A1(\inst$top.soc.gpio_0._gpio.w_data$50 ),
    .A2(_17759_),
    .B1(net2167),
    .Y(_17772_));
 sky130_fd_sc_hd__a21oi_1 _39630_ (.A1(_02896_),
    .A2(_17759_),
    .B1(_17772_),
    .Y(_05051_));
 sky130_fd_sc_hd__inv_1 _39631_ (.A(\inst$top.soc.gpio_0._gpio.w_data$53 ),
    .Y(_17773_));
 sky130_fd_sc_hd__o21ai_0 _39632_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__3._storage[1] ),
    .A2(net2585),
    .B1(net2167),
    .Y(_17774_));
 sky130_fd_sc_hd__a21oi_1 _39633_ (.A1(_17773_),
    .A2(net2585),
    .B1(_17774_),
    .Y(_05052_));
 sky130_fd_sc_hd__inv_1 _39634_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__0.port__w_data ),
    .Y(_17775_));
 sky130_fd_sc_hd__o21ai_0 _39635_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__4._storage[0] ),
    .A2(net2585),
    .B1(net2168),
    .Y(_17776_));
 sky130_fd_sc_hd__a21oi_1 _39636_ (.A1(_17775_),
    .A2(net2584),
    .B1(_17776_),
    .Y(_05053_));
 sky130_fd_sc_hd__inv_1 _39637_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__1.port__w_data ),
    .Y(_17777_));
 sky130_fd_sc_hd__o21ai_0 _39639_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__4._storage[1] ),
    .A2(net2585),
    .B1(net2169),
    .Y(_17779_));
 sky130_fd_sc_hd__a21oi_1 _39640_ (.A1(_17777_),
    .A2(net2584),
    .B1(_17779_),
    .Y(_05054_));
 sky130_fd_sc_hd__inv_1 _39641_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__2.port__w_data ),
    .Y(_17780_));
 sky130_fd_sc_hd__o21ai_0 _39642_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__5._storage[0] ),
    .A2(net2586),
    .B1(net2163),
    .Y(_17781_));
 sky130_fd_sc_hd__a21oi_1 _39643_ (.A1(_17780_),
    .A2(net2586),
    .B1(_17781_),
    .Y(_05055_));
 sky130_fd_sc_hd__inv_1 _39644_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__3.port__w_data ),
    .Y(_17782_));
 sky130_fd_sc_hd__o21ai_0 _39645_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__5._storage[1] ),
    .A2(net2586),
    .B1(net2167),
    .Y(_17783_));
 sky130_fd_sc_hd__a21oi_1 _39646_ (.A1(_17782_),
    .A2(net2586),
    .B1(_17783_),
    .Y(_05056_));
 sky130_fd_sc_hd__inv_1 _39647_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__4.port__w_data ),
    .Y(_17784_));
 sky130_fd_sc_hd__o21ai_0 _39648_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__6._storage[0] ),
    .A2(net2584),
    .B1(net2169),
    .Y(_17785_));
 sky130_fd_sc_hd__a21oi_1 _39649_ (.A1(_17784_),
    .A2(net2584),
    .B1(_17785_),
    .Y(_05057_));
 sky130_fd_sc_hd__inv_1 _39650_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__5.port__w_data ),
    .Y(_17786_));
 sky130_fd_sc_hd__o21ai_0 _39651_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__6._storage[1] ),
    .A2(net2584),
    .B1(net2168),
    .Y(_17787_));
 sky130_fd_sc_hd__a21oi_1 _39652_ (.A1(_17786_),
    .A2(net2584),
    .B1(_17787_),
    .Y(_05058_));
 sky130_fd_sc_hd__inv_1 _39653_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__6.port__w_data ),
    .Y(_17788_));
 sky130_fd_sc_hd__o21ai_0 _39654_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__7._storage[0] ),
    .A2(net2584),
    .B1(net2168),
    .Y(_17789_));
 sky130_fd_sc_hd__a21oi_1 _39655_ (.A1(_17788_),
    .A2(net2584),
    .B1(_17789_),
    .Y(_05059_));
 sky130_fd_sc_hd__inv_1 _39656_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__7.port__w_data ),
    .Y(_17790_));
 sky130_fd_sc_hd__o21ai_0 _39657_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__7._storage[1] ),
    .A2(net2584),
    .B1(net2168),
    .Y(_17791_));
 sky130_fd_sc_hd__a21oi_1 _39658_ (.A1(_17790_),
    .A2(net2584),
    .B1(_17791_),
    .Y(_05060_));
 sky130_fd_sc_hd__inv_1 _39659_ (.A(net2587),
    .Y(_17792_));
 sky130_fd_sc_hd__nor3_1 _39660_ (.A(\inst$top.soc.gpio_0._gpio.w_data ),
    .B(_17792_),
    .C(_17761_),
    .Y(_17793_));
 sky130_fd_sc_hd__inv_1 _39663_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__0._storage ),
    .Y(_17796_));
 sky130_fd_sc_hd__nand2_1 _39664_ (.A(net2589),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__0.port__w_data ),
    .Y(_17797_));
 sky130_fd_sc_hd__o21ai_0 _39665_ (.A1(net2589),
    .A2(_17796_),
    .B1(_17797_),
    .Y(_17798_));
 sky130_fd_sc_hd__a31oi_1 _39666_ (.A1(\inst$top.soc.gpio_0._gpio.w_data ),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb$21 ),
    .A3(_17761_),
    .B1(_17798_),
    .Y(_17799_));
 sky130_fd_sc_hd__nor3_1 _39667_ (.A(net3002),
    .B(_17793_),
    .C(_17799_),
    .Y(_05061_));
 sky130_fd_sc_hd__nor3_1 _39668_ (.A(\inst$top.soc.gpio_0._gpio.w_data$26 ),
    .B(_17792_),
    .C(_17766_),
    .Y(_17800_));
 sky130_fd_sc_hd__inv_1 _39669_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__1._storage ),
    .Y(_17801_));
 sky130_fd_sc_hd__nand2_1 _39670_ (.A(net2589),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__1.port__w_data ),
    .Y(_17802_));
 sky130_fd_sc_hd__o21ai_0 _39671_ (.A1(net2589),
    .A2(_17801_),
    .B1(_17802_),
    .Y(_17803_));
 sky130_fd_sc_hd__a31oi_1 _39672_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb$21 ),
    .A2(\inst$top.soc.gpio_0._gpio.w_data$26 ),
    .A3(_17766_),
    .B1(_17803_),
    .Y(_17804_));
 sky130_fd_sc_hd__nor3_1 _39673_ (.A(net3002),
    .B(_17800_),
    .C(_17804_),
    .Y(_05062_));
 sky130_fd_sc_hd__inv_1 _39674_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__2._storage ),
    .Y(_17805_));
 sky130_fd_sc_hd__nand2_1 _39675_ (.A(net2588),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__2.port__w_data ),
    .Y(_17806_));
 sky130_fd_sc_hd__o21ai_0 _39676_ (.A1(net2588),
    .A2(_17805_),
    .B1(_17806_),
    .Y(_17807_));
 sky130_fd_sc_hd__a31oi_1 _39677_ (.A1(net2587),
    .A2(\inst$top.soc.gpio_0._gpio.w_data$38 ),
    .A3(_17770_),
    .B1(_17807_),
    .Y(_17808_));
 sky130_fd_sc_hd__a311oi_1 _39678_ (.A1(net2587),
    .A2(_17768_),
    .A3(\inst$top.soc.gpio_0._gpio.w_data$41 ),
    .B1(net2997),
    .C1(_17808_),
    .Y(_05063_));
 sky130_fd_sc_hd__nor3_1 _39679_ (.A(\inst$top.soc.gpio_0._gpio.w_data$50 ),
    .B(_17792_),
    .C(_17773_),
    .Y(_17809_));
 sky130_fd_sc_hd__inv_1 _39680_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__3._storage ),
    .Y(_17810_));
 sky130_fd_sc_hd__nand2_1 _39681_ (.A(net2588),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__3.port__w_data ),
    .Y(_17811_));
 sky130_fd_sc_hd__o21ai_0 _39682_ (.A1(net2588),
    .A2(_17810_),
    .B1(_17811_),
    .Y(_17812_));
 sky130_fd_sc_hd__a31oi_1 _39683_ (.A1(net2587),
    .A2(\inst$top.soc.gpio_0._gpio.w_data$50 ),
    .A3(_17773_),
    .B1(_17812_),
    .Y(_17813_));
 sky130_fd_sc_hd__nor3_1 _39684_ (.A(net3001),
    .B(_17809_),
    .C(_17813_),
    .Y(_05064_));
 sky130_fd_sc_hd__inv_1 _39685_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__4._storage ),
    .Y(_17814_));
 sky130_fd_sc_hd__nand2_1 _39686_ (.A(net2588),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__4.port__w_data ),
    .Y(_17815_));
 sky130_fd_sc_hd__o21ai_0 _39687_ (.A1(net2589),
    .A2(_17814_),
    .B1(_17815_),
    .Y(_17816_));
 sky130_fd_sc_hd__a31oi_1 _39688_ (.A1(net2587),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__0.port__w_data ),
    .A3(_17777_),
    .B1(_17816_),
    .Y(_17817_));
 sky130_fd_sc_hd__a311oi_1 _39689_ (.A1(net2587),
    .A2(_17775_),
    .A3(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__1.port__w_data ),
    .B1(net3002),
    .C1(_17817_),
    .Y(_05065_));
 sky130_fd_sc_hd__inv_1 _39690_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__5._storage ),
    .Y(_17818_));
 sky130_fd_sc_hd__nand2_1 _39691_ (.A(net2588),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__5.port__w_data ),
    .Y(_17819_));
 sky130_fd_sc_hd__o21ai_0 _39692_ (.A1(net2588),
    .A2(_17818_),
    .B1(_17819_),
    .Y(_17820_));
 sky130_fd_sc_hd__a31oi_1 _39693_ (.A1(net2587),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__2.port__w_data ),
    .A3(_17782_),
    .B1(_17820_),
    .Y(_17821_));
 sky130_fd_sc_hd__a311oi_1 _39694_ (.A1(net2587),
    .A2(_17780_),
    .A3(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__3.port__w_data ),
    .B1(net3001),
    .C1(_17821_),
    .Y(_05066_));
 sky130_fd_sc_hd__inv_1 _39695_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__6._storage ),
    .Y(_17822_));
 sky130_fd_sc_hd__nand2_1 _39696_ (.A(net2588),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__6.port__w_data ),
    .Y(_17823_));
 sky130_fd_sc_hd__o21ai_0 _39697_ (.A1(net2588),
    .A2(_17822_),
    .B1(_17823_),
    .Y(_17824_));
 sky130_fd_sc_hd__a31oi_1 _39698_ (.A1(net2587),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__4.port__w_data ),
    .A3(_17786_),
    .B1(_17824_),
    .Y(_17825_));
 sky130_fd_sc_hd__a311oi_1 _39699_ (.A1(net2587),
    .A2(_17784_),
    .A3(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__5.port__w_data ),
    .B1(net3002),
    .C1(_17825_),
    .Y(_05067_));
 sky130_fd_sc_hd__o221ai_1 _39700_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__7._storage ),
    .A2(net2589),
    .B1(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__6.port__w_data ),
    .B2(_17792_),
    .C1(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__7.port__w_data ),
    .Y(_17826_));
 sky130_fd_sc_hd__inv_1 _39701_ (.A(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__7._storage ),
    .Y(_17827_));
 sky130_fd_sc_hd__o22ai_1 _39702_ (.A1(net2588),
    .A2(_17827_),
    .B1(_17792_),
    .B2(_17788_),
    .Y(_17828_));
 sky130_fd_sc_hd__nand2_1 _39703_ (.A(_17828_),
    .B(_17790_),
    .Y(_17829_));
 sky130_fd_sc_hd__a21oi_1 _39704_ (.A1(_17826_),
    .A2(_17829_),
    .B1(net3002),
    .Y(_05068_));
 sky130_fd_sc_hd__nor2_2 _39705_ (.A(\inst$top.soc.bus__addr[2] ),
    .B(\inst$top.soc.bus__addr[3] ),
    .Y(_17830_));
 sky130_fd_sc_hd__nand2_1 _39706_ (.A(\inst$top.soc.wb_to_csr.cycle[0] ),
    .B(\inst$top.soc.wb_to_csr.cycle[1] ),
    .Y(_17831_));
 sky130_fd_sc_hd__nor2_1 _39707_ (.A(net2989),
    .B(_17831_),
    .Y(_17832_));
 sky130_fd_sc_hd__nand2_1 _39708_ (.A(_17830_),
    .B(_17832_),
    .Y(_17833_));
 sky130_fd_sc_hd__inv_1 _39709_ (.A(_09300_),
    .Y(_17834_));
 sky130_fd_sc_hd__nor3_1 _39710_ (.A(_09277_),
    .B(_09298_),
    .C(_17834_),
    .Y(_17835_));
 sky130_fd_sc_hd__inv_1 _39711_ (.A(_17835_),
    .Y(_17836_));
 sky130_fd_sc_hd__nor2_1 _39712_ (.A(\inst$top.soc.bus__adr[4] ),
    .B(\inst$top.soc.bus__adr[3] ),
    .Y(_17837_));
 sky130_fd_sc_hd__inv_1 _39713_ (.A(_17837_),
    .Y(_17838_));
 sky130_fd_sc_hd__nand2_1 _39714_ (.A(_09293_),
    .B(_09332_),
    .Y(_17839_));
 sky130_fd_sc_hd__nor4_1 _39715_ (.A(_17838_),
    .B(_09288_),
    .C(_09326_),
    .D(_17839_),
    .Y(_17840_));
 sky130_fd_sc_hd__nor2_1 _39716_ (.A(\inst$top.soc.bus__adr[5] ),
    .B(\inst$top.soc.bus__adr[6] ),
    .Y(_17841_));
 sky130_fd_sc_hd__inv_1 _39717_ (.A(_17841_),
    .Y(_17842_));
 sky130_fd_sc_hd__nor3_1 _39718_ (.A(\inst$top.soc.bus__adr[7] ),
    .B(\inst$top.soc.bus__adr[2] ),
    .C(_17842_),
    .Y(_17843_));
 sky130_fd_sc_hd__nand2_1 _39719_ (.A(_17840_),
    .B(_17843_),
    .Y(_17844_));
 sky130_fd_sc_hd__nor3_2 _39720_ (.A(_09270_),
    .B(_17836_),
    .C(_17844_),
    .Y(_17845_));
 sky130_fd_sc_hd__nor2_1 _39721_ (.A(\inst$top.soc.wb_to_csr.cycle[2] ),
    .B(_17831_),
    .Y(_17846_));
 sky130_fd_sc_hd__inv_1 _39722_ (.A(_17846_),
    .Y(_17847_));
 sky130_fd_sc_hd__a21oi_1 _39723_ (.A1(net2563),
    .A2(_09350_),
    .B1(_17847_),
    .Y(_17848_));
 sky130_fd_sc_hd__inv_1 _39724_ (.A(\inst$top.soc.wb_to_csr.cycle[0] ),
    .Y(_17849_));
 sky130_fd_sc_hd__nor2_2 _39725_ (.A(\inst$top.soc.wb_to_csr.cycle[1] ),
    .B(_17849_),
    .Y(_17850_));
 sky130_fd_sc_hd__inv_1 _39726_ (.A(_17850_),
    .Y(_17851_));
 sky130_fd_sc_hd__nor2_1 _39727_ (.A(\inst$top.soc.wb_to_csr.cycle[2] ),
    .B(_17851_),
    .Y(_17852_));
 sky130_fd_sc_hd__o21ai_0 _39728_ (.A1(net2557),
    .A2(\inst$top.soc.cpu.loadstore.dbus__sel[1] ),
    .B1(_17852_),
    .Y(_17853_));
 sky130_fd_sc_hd__inv_1 _39729_ (.A(\inst$top.soc.wb_to_csr.cycle[1] ),
    .Y(_17854_));
 sky130_fd_sc_hd__nor2_2 _39730_ (.A(\inst$top.soc.wb_to_csr.cycle[0] ),
    .B(_17854_),
    .Y(_17855_));
 sky130_fd_sc_hd__inv_1 _39731_ (.A(_17855_),
    .Y(_17856_));
 sky130_fd_sc_hd__nor2_2 _39732_ (.A(\inst$top.soc.wb_to_csr.cycle[2] ),
    .B(_17856_),
    .Y(_17857_));
 sky130_fd_sc_hd__o21ai_0 _39733_ (.A1(net2557),
    .A2(\inst$top.soc.cpu.loadstore.dbus__sel[2] ),
    .B1(_17857_),
    .Y(_17858_));
 sky130_fd_sc_hd__nor2_2 _39734_ (.A(\inst$top.soc.wb_to_csr.cycle[0] ),
    .B(\inst$top.soc.wb_to_csr.cycle[1] ),
    .Y(_17859_));
 sky130_fd_sc_hd__o22ai_1 _39735_ (.A1(\inst$top.soc.cpu.loadstore.dbus__sel[0] ),
    .A2(net2557),
    .B1(\inst$top.soc.wb_to_csr.cycle[2] ),
    .B2(_17859_),
    .Y(_17860_));
 sky130_fd_sc_hd__nand3_1 _39736_ (.A(_17853_),
    .B(_17858_),
    .C(_17860_),
    .Y(_17861_));
 sky130_fd_sc_hd__nor2_1 _39737_ (.A(_17848_),
    .B(_17861_),
    .Y(_17862_));
 sky130_fd_sc_hd__nor2_2 _39738_ (.A(_09345_),
    .B(net1085),
    .Y(_17863_));
 sky130_fd_sc_hd__inv_1 _39739_ (.A(\inst$top.soc.wb_to_csr.cycle[2] ),
    .Y(_17864_));
 sky130_fd_sc_hd__nand2_1 _39740_ (.A(_17863_),
    .B(_17864_),
    .Y(_17865_));
 sky130_fd_sc_hd__nor3_1 _39741_ (.A(_09256_),
    .B(_17862_),
    .C(_17865_),
    .Y(_17866_));
 sky130_fd_sc_hd__nand2_1 _39742_ (.A(_17845_),
    .B(_17866_),
    .Y(_17867_));
 sky130_fd_sc_hd__nor2_1 _39743_ (.A(_17833_),
    .B(_17867_),
    .Y(_05069_));
 sky130_fd_sc_hd__inv_1 _39744_ (.A(\inst$top.soc.bus__addr[2] ),
    .Y(_17868_));
 sky130_fd_sc_hd__nor2_1 _39745_ (.A(_17868_),
    .B(\inst$top.soc.bus__addr[3] ),
    .Y(_17869_));
 sky130_fd_sc_hd__inv_1 _39746_ (.A(_17869_),
    .Y(_17870_));
 sky130_fd_sc_hd__nor2_1 _39747_ (.A(_17851_),
    .B(_17870_),
    .Y(_17871_));
 sky130_fd_sc_hd__nand2_1 _39748_ (.A(_17871_),
    .B(net2137),
    .Y(_17872_));
 sky130_fd_sc_hd__nor2_1 _39749_ (.A(_17872_),
    .B(_17867_),
    .Y(_05070_));
 sky130_fd_sc_hd__nand3_1 _39750_ (.A(_17830_),
    .B(net2137),
    .C(_17850_),
    .Y(_17873_));
 sky130_fd_sc_hd__nor2_1 _39751_ (.A(_17873_),
    .B(_17867_),
    .Y(_05071_));
 sky130_fd_sc_hd__clkinv_1 _39752_ (.A(_17830_),
    .Y(_17874_));
 sky130_fd_sc_hd__nor2_1 _39753_ (.A(_17862_),
    .B(_17865_),
    .Y(_17875_));
 sky130_fd_sc_hd__nand2_1 _39754_ (.A(_17875_),
    .B(_09256_),
    .Y(_17876_));
 sky130_fd_sc_hd__nor2_1 _39755_ (.A(_17874_),
    .B(_17876_),
    .Y(_17877_));
 sky130_fd_sc_hd__nand3_1 _39756_ (.A(_17845_),
    .B(_17849_),
    .C(_17877_),
    .Y(_17878_));
 sky130_fd_sc_hd__nor2_1 _39757_ (.A(_17856_),
    .B(_17874_),
    .Y(_17879_));
 sky130_fd_sc_hd__inv_1 _39758_ (.A(_17879_),
    .Y(_17880_));
 sky130_fd_sc_hd__nor3_1 _39759_ (.A(_09270_),
    .B(_17836_),
    .C(_17844_),
    .Y(_17881_));
 sky130_fd_sc_hd__clkinv_1 _39760_ (.A(_17876_),
    .Y(_17882_));
 sky130_fd_sc_hd__nand2_1 _39761_ (.A(_17881_),
    .B(_17882_),
    .Y(_17883_));
 sky130_fd_sc_hd__nor2_1 _39762_ (.A(_17880_),
    .B(_17883_),
    .Y(_17884_));
 sky130_fd_sc_hd__inv_1 _39763_ (.A(_17859_),
    .Y(_17885_));
 sky130_fd_sc_hd__nor2_1 _39764_ (.A(_17885_),
    .B(_17874_),
    .Y(_17886_));
 sky130_fd_sc_hd__inv_1 _39765_ (.A(_17886_),
    .Y(_17887_));
 sky130_fd_sc_hd__nor2_2 _39766_ (.A(_17887_),
    .B(_17883_),
    .Y(_17888_));
 sky130_fd_sc_hd__inv_1 _39767_ (.A(_17888_),
    .Y(_17889_));
 sky130_fd_sc_hd__nor2_1 _39768_ (.A(_02871_),
    .B(_17889_),
    .Y(_17890_));
 sky130_fd_sc_hd__a221oi_1 _39769_ (.A1(_17878_),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[0] ),
    .B1(\inst$top.soc.gpio_0._gpio.r_data ),
    .B2(_17884_),
    .C1(_17890_),
    .Y(_17891_));
 sky130_fd_sc_hd__nor2_2 _39770_ (.A(net3001),
    .B(_17891_),
    .Y(_05072_));
 sky130_fd_sc_hd__nand2_1 _39771_ (.A(_17884_),
    .B(\inst$top.soc.gpio_0._gpio.r_data$23 ),
    .Y(_17892_));
 sky130_fd_sc_hd__nand2_1 _39772_ (.A(_17888_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__0._storage[1] ),
    .Y(_17893_));
 sky130_fd_sc_hd__nand2_1 _39773_ (.A(_17878_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[1] ),
    .Y(_17894_));
 sky130_fd_sc_hd__a31oi_1 _39774_ (.A1(_17892_),
    .A2(_17893_),
    .A3(_17894_),
    .B1(net3001),
    .Y(_05073_));
 sky130_fd_sc_hd__nor2_1 _39775_ (.A(_02893_),
    .B(_17889_),
    .Y(_17895_));
 sky130_fd_sc_hd__a221oi_1 _39776_ (.A1(_17878_),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[2] ),
    .B1(\inst$top.soc.gpio_0._gpio.r_data$35 ),
    .B2(_17884_),
    .C1(_17895_),
    .Y(_17896_));
 sky130_fd_sc_hd__nor2_2 _39777_ (.A(net3001),
    .B(_17896_),
    .Y(_05074_));
 sky130_fd_sc_hd__nand2_1 _39778_ (.A(_17884_),
    .B(\inst$top.soc.gpio_0._gpio.r_data$47 ),
    .Y(_17897_));
 sky130_fd_sc_hd__nand2_1 _39779_ (.A(_17888_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__1._storage[1] ),
    .Y(_17898_));
 sky130_fd_sc_hd__nand2_1 _39780_ (.A(_17878_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[3] ),
    .Y(_17899_));
 sky130_fd_sc_hd__a31oi_1 _39781_ (.A1(_17897_),
    .A2(_17898_),
    .A3(_17899_),
    .B1(net3001),
    .Y(_05075_));
 sky130_fd_sc_hd__nor2_1 _39782_ (.A(_02868_),
    .B(_17889_),
    .Y(_17900_));
 sky130_fd_sc_hd__a221oi_1 _39783_ (.A1(_17878_),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[4] ),
    .B1(\inst$top.soc.gpio_0._gpio.r_data$59 ),
    .B2(_17884_),
    .C1(_17900_),
    .Y(_17901_));
 sky130_fd_sc_hd__nor2_2 _39784_ (.A(net2997),
    .B(_17901_),
    .Y(_05076_));
 sky130_fd_sc_hd__nand2_1 _39785_ (.A(_17884_),
    .B(\inst$top.soc.gpio_0._gpio.r_data$71 ),
    .Y(_17902_));
 sky130_fd_sc_hd__nand2_1 _39786_ (.A(_17888_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__2._storage[1] ),
    .Y(_17903_));
 sky130_fd_sc_hd__nand2_1 _39787_ (.A(_17878_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[5] ),
    .Y(_17904_));
 sky130_fd_sc_hd__a31oi_1 _39788_ (.A1(_17902_),
    .A2(_17903_),
    .A3(_17904_),
    .B1(net2997),
    .Y(_05077_));
 sky130_fd_sc_hd__nor2_1 _39789_ (.A(_02896_),
    .B(_17889_),
    .Y(_17905_));
 sky130_fd_sc_hd__a221oi_1 _39790_ (.A1(_17878_),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[6] ),
    .B1(\inst$top.soc.gpio_0._gpio.r_data$83 ),
    .B2(_17884_),
    .C1(_17905_),
    .Y(_17906_));
 sky130_fd_sc_hd__nor2_2 _39791_ (.A(net3001),
    .B(_17906_),
    .Y(_05078_));
 sky130_fd_sc_hd__nand2_1 _39792_ (.A(_17884_),
    .B(\inst$top.soc.gpio_0._gpio.r_data$95 ),
    .Y(_17907_));
 sky130_fd_sc_hd__nand2_1 _39793_ (.A(_17888_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__3._storage[1] ),
    .Y(_17908_));
 sky130_fd_sc_hd__nand2_1 _39794_ (.A(_17878_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[7] ),
    .Y(_17909_));
 sky130_fd_sc_hd__a31oi_1 _39795_ (.A1(_17907_),
    .A2(_17908_),
    .A3(_17909_),
    .B1(net3001),
    .Y(_05079_));
 sky130_fd_sc_hd__nor2_1 _39796_ (.A(net2997),
    .B(_17878_),
    .Y(_05080_));
 sky130_fd_sc_hd__nor2_1 _39798_ (.A(_17831_),
    .B(_17874_),
    .Y(_17911_));
 sky130_fd_sc_hd__o211ai_1 _39799_ (.A1(_17911_),
    .A2(_17886_),
    .B1(_17882_),
    .C1(_17845_),
    .Y(_17912_));
 sky130_fd_sc_hd__nand3_1 _39800_ (.A(_17881_),
    .B(_17911_),
    .C(_17882_),
    .Y(_17913_));
 sky130_fd_sc_hd__o22ai_1 _39801_ (.A1(_17796_),
    .A2(_17913_),
    .B1(_02908_),
    .B2(_17889_),
    .Y(_17914_));
 sky130_fd_sc_hd__a21oi_1 _39802_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[0] ),
    .A2(_17912_),
    .B1(_17914_),
    .Y(_17915_));
 sky130_fd_sc_hd__nor2_2 _39803_ (.A(net2998),
    .B(_17915_),
    .Y(_05081_));
 sky130_fd_sc_hd__nor2_1 _39804_ (.A(_17801_),
    .B(_17913_),
    .Y(_17916_));
 sky130_fd_sc_hd__a221oi_1 _39805_ (.A1(_17888_),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__4._storage[1] ),
    .B1(_17912_),
    .B2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[1] ),
    .C1(_17916_),
    .Y(_17917_));
 sky130_fd_sc_hd__nor2_1 _39806_ (.A(net3002),
    .B(_17917_),
    .Y(_05082_));
 sky130_fd_sc_hd__o22ai_1 _39807_ (.A1(_17805_),
    .A2(_17913_),
    .B1(_02905_),
    .B2(_17889_),
    .Y(_17918_));
 sky130_fd_sc_hd__a21oi_1 _39808_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[2] ),
    .A2(_17912_),
    .B1(_17918_),
    .Y(_17919_));
 sky130_fd_sc_hd__nor2_2 _39809_ (.A(net2998),
    .B(_17919_),
    .Y(_05083_));
 sky130_fd_sc_hd__nor2_1 _39810_ (.A(_17810_),
    .B(_17913_),
    .Y(_17920_));
 sky130_fd_sc_hd__a221oi_1 _39811_ (.A1(_17888_),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__5._storage[1] ),
    .B1(_17912_),
    .B2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[3] ),
    .C1(_17920_),
    .Y(_17921_));
 sky130_fd_sc_hd__nor2_1 _39812_ (.A(net3001),
    .B(_17921_),
    .Y(_05084_));
 sky130_fd_sc_hd__o22ai_1 _39813_ (.A1(_17814_),
    .A2(_17913_),
    .B1(_02902_),
    .B2(_17889_),
    .Y(_17922_));
 sky130_fd_sc_hd__a21oi_1 _39814_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[4] ),
    .A2(_17912_),
    .B1(_17922_),
    .Y(_17923_));
 sky130_fd_sc_hd__nor2_2 _39815_ (.A(net2997),
    .B(_17923_),
    .Y(_05085_));
 sky130_fd_sc_hd__nor2_1 _39816_ (.A(_17818_),
    .B(_17913_),
    .Y(_17924_));
 sky130_fd_sc_hd__a221oi_1 _39817_ (.A1(_17888_),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__6._storage[1] ),
    .B1(_17912_),
    .B2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[5] ),
    .C1(_17924_),
    .Y(_17925_));
 sky130_fd_sc_hd__nor2_1 _39818_ (.A(net2997),
    .B(_17925_),
    .Y(_05086_));
 sky130_fd_sc_hd__o22ai_1 _39819_ (.A1(_17822_),
    .A2(_17913_),
    .B1(_02899_),
    .B2(_17889_),
    .Y(_17926_));
 sky130_fd_sc_hd__a21oi_1 _39820_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[6] ),
    .A2(_17912_),
    .B1(_17926_),
    .Y(_17927_));
 sky130_fd_sc_hd__nor2_2 _39821_ (.A(net2997),
    .B(_17927_),
    .Y(_05087_));
 sky130_fd_sc_hd__nor2_1 _39822_ (.A(_17827_),
    .B(_17913_),
    .Y(_17928_));
 sky130_fd_sc_hd__a221oi_1 _39823_ (.A1(_17888_),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__7._storage[1] ),
    .B1(_17912_),
    .B2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[7] ),
    .C1(_17928_),
    .Y(_17929_));
 sky130_fd_sc_hd__nor2_1 _39824_ (.A(net3001),
    .B(_17929_),
    .Y(_05088_));
 sky130_fd_sc_hd__nand2_1 _39825_ (.A(_17845_),
    .B(_17882_),
    .Y(_17930_));
 sky130_fd_sc_hd__nor4_2 _39826_ (.A(_17849_),
    .B(net2989),
    .C(_17874_),
    .D(_17930_),
    .Y(_05089_));
 sky130_fd_sc_hd__nor2_1 _39827_ (.A(_17885_),
    .B(\inst$top.soc.bus__addr[3] ),
    .Y(_17931_));
 sky130_fd_sc_hd__inv_1 _39828_ (.A(_17931_),
    .Y(_17932_));
 sky130_fd_sc_hd__nor2_1 _39829_ (.A(_17932_),
    .B(_17867_),
    .Y(_17933_));
 sky130_fd_sc_hd__nor2_1 _39831_ (.A(\inst$top.soc.wb_to_csr.cycle[2] ),
    .B(_17885_),
    .Y(_17935_));
 sky130_fd_sc_hd__inv_1 _39832_ (.A(_17935_),
    .Y(_17936_));
 sky130_fd_sc_hd__nand2_1 _39833_ (.A(_17857_),
    .B(\inst$top.soc.bus__dat_w[16] ),
    .Y(_17937_));
 sky130_fd_sc_hd__o21ai_0 _39834_ (.A1(_07435_),
    .A2(_17936_),
    .B1(_17937_),
    .Y(_17938_));
 sky130_fd_sc_hd__inv_1 _39835_ (.A(_17852_),
    .Y(_17939_));
 sky130_fd_sc_hd__o22ai_1 _39836_ (.A1(_07430_),
    .A2(_17847_),
    .B1(_07434_),
    .B2(_17939_),
    .Y(_17940_));
 sky130_fd_sc_hd__o21ai_4 _39837_ (.A1(_17938_),
    .A2(_17940_),
    .B1(_17863_),
    .Y(_17941_));
 sky130_fd_sc_hd__o21ai_0 _39839_ (.A1(\inst$top.soc.gpio_0._gpio.w_data ),
    .A2(net845),
    .B1(net2168),
    .Y(_17943_));
 sky130_fd_sc_hd__a21oi_2 _39840_ (.A1(net845),
    .A2(net900),
    .B1(_17943_),
    .Y(_05090_));
 sky130_fd_sc_hd__nand2_1 _39841_ (.A(_17857_),
    .B(\inst$top.soc.bus__dat_w[17] ),
    .Y(_17944_));
 sky130_fd_sc_hd__o21ai_0 _39842_ (.A1(_07436_),
    .A2(_17847_),
    .B1(_17944_),
    .Y(_17945_));
 sky130_fd_sc_hd__o22ai_1 _39843_ (.A1(_07439_),
    .A2(_17936_),
    .B1(_07438_),
    .B2(_17939_),
    .Y(_17946_));
 sky130_fd_sc_hd__inv_1 _39844_ (.A(_17865_),
    .Y(_17947_));
 sky130_fd_sc_hd__o21ai_4 _39845_ (.A1(_17945_),
    .A2(_17946_),
    .B1(_17947_),
    .Y(_17948_));
 sky130_fd_sc_hd__o21ai_0 _39847_ (.A1(\inst$top.soc.gpio_0._gpio.w_data$16 ),
    .A2(net844),
    .B1(net2168),
    .Y(_17950_));
 sky130_fd_sc_hd__a21oi_2 _39848_ (.A1(net844),
    .A2(net868),
    .B1(_17950_),
    .Y(_05091_));
 sky130_fd_sc_hd__nand2_1 _39849_ (.A(_17857_),
    .B(\inst$top.soc.bus__dat_w[18] ),
    .Y(_17951_));
 sky130_fd_sc_hd__o21ai_0 _39850_ (.A1(_07443_),
    .A2(_17936_),
    .B1(_17951_),
    .Y(_17952_));
 sky130_fd_sc_hd__o22ai_1 _39851_ (.A1(_07440_),
    .A2(_17847_),
    .B1(_07442_),
    .B2(_17939_),
    .Y(_17953_));
 sky130_fd_sc_hd__o21ai_4 _39852_ (.A1(_17952_),
    .A2(_17953_),
    .B1(_17863_),
    .Y(_17954_));
 sky130_fd_sc_hd__o21ai_0 _39854_ (.A1(\inst$top.soc.gpio_0._gpio.w_data$26 ),
    .A2(net844),
    .B1(net2167),
    .Y(_17956_));
 sky130_fd_sc_hd__a21oi_1 _39855_ (.A1(net844),
    .A2(_17954_),
    .B1(_17956_),
    .Y(_05092_));
 sky130_fd_sc_hd__nand2_1 _39856_ (.A(_17857_),
    .B(\inst$top.soc.bus__dat_w[19] ),
    .Y(_17957_));
 sky130_fd_sc_hd__o21ai_0 _39857_ (.A1(_07447_),
    .A2(_17936_),
    .B1(_17957_),
    .Y(_17958_));
 sky130_fd_sc_hd__o22ai_1 _39858_ (.A1(_07444_),
    .A2(_17847_),
    .B1(_07446_),
    .B2(_17939_),
    .Y(_17959_));
 sky130_fd_sc_hd__o21ai_4 _39859_ (.A1(_17958_),
    .A2(_17959_),
    .B1(_17863_),
    .Y(_17960_));
 sky130_fd_sc_hd__o21ai_0 _39862_ (.A1(\inst$top.soc.gpio_0._gpio.w_data$29 ),
    .A2(net844),
    .B1(net2170),
    .Y(_17963_));
 sky130_fd_sc_hd__a21oi_1 _39863_ (.A1(net844),
    .A2(_17960_),
    .B1(_17963_),
    .Y(_05093_));
 sky130_fd_sc_hd__nand2_1 _39864_ (.A(_17857_),
    .B(\inst$top.soc.bus__dat_w[20] ),
    .Y(_17964_));
 sky130_fd_sc_hd__o21ai_0 _39865_ (.A1(_07448_),
    .A2(_17847_),
    .B1(_17964_),
    .Y(_17965_));
 sky130_fd_sc_hd__o22ai_1 _39866_ (.A1(_07451_),
    .A2(_17936_),
    .B1(_07450_),
    .B2(_17939_),
    .Y(_17966_));
 sky130_fd_sc_hd__o21ai_4 _39867_ (.A1(_17965_),
    .A2(_17966_),
    .B1(_17947_),
    .Y(_17967_));
 sky130_fd_sc_hd__o21ai_0 _39869_ (.A1(\inst$top.soc.gpio_0._gpio.w_data$38 ),
    .A2(net845),
    .B1(net2163),
    .Y(_17969_));
 sky130_fd_sc_hd__a21oi_1 _39870_ (.A1(net845),
    .A2(net867),
    .B1(_17969_),
    .Y(_05094_));
 sky130_fd_sc_hd__a22oi_1 _39871_ (.A1(\inst$top.soc.bus__dat_w[29] ),
    .A2(_17846_),
    .B1(_17857_),
    .B2(\inst$top.soc.bus__dat_w[21] ),
    .Y(_17970_));
 sky130_fd_sc_hd__o221ai_1 _39872_ (.A1(_07455_),
    .A2(_17936_),
    .B1(_07454_),
    .B2(_17939_),
    .C1(_17970_),
    .Y(_17971_));
 sky130_fd_sc_hd__nand2_1 _39873_ (.A(_17971_),
    .B(_17947_),
    .Y(_17972_));
 sky130_fd_sc_hd__o21ai_0 _39874_ (.A1(\inst$top.soc.gpio_0._gpio.w_data$41 ),
    .A2(net845),
    .B1(net2163),
    .Y(_17973_));
 sky130_fd_sc_hd__a21oi_1 _39875_ (.A1(net845),
    .A2(_17972_),
    .B1(_17973_),
    .Y(_05095_));
 sky130_fd_sc_hd__nand2_1 _39876_ (.A(_17857_),
    .B(\inst$top.soc.bus__dat_w[22] ),
    .Y(_17974_));
 sky130_fd_sc_hd__o21ai_0 _39877_ (.A1(_07456_),
    .A2(_17847_),
    .B1(_17974_),
    .Y(_17975_));
 sky130_fd_sc_hd__o22ai_1 _39878_ (.A1(_07459_),
    .A2(_17936_),
    .B1(_07458_),
    .B2(_17939_),
    .Y(_17976_));
 sky130_fd_sc_hd__o21ai_4 _39879_ (.A1(_17975_),
    .A2(_17976_),
    .B1(_17947_),
    .Y(_17977_));
 sky130_fd_sc_hd__o21ai_0 _39881_ (.A1(\inst$top.soc.gpio_0._gpio.w_data$50 ),
    .A2(net844),
    .B1(net2167),
    .Y(_17979_));
 sky130_fd_sc_hd__a21oi_1 _39882_ (.A1(net844),
    .A2(_17977_),
    .B1(_17979_),
    .Y(_05096_));
 sky130_fd_sc_hd__a22oi_1 _39883_ (.A1(\inst$top.soc.bus__dat_w[31] ),
    .A2(_17846_),
    .B1(_17857_),
    .B2(\inst$top.soc.bus__dat_w[23] ),
    .Y(_17980_));
 sky130_fd_sc_hd__o221ai_1 _39884_ (.A1(_07463_),
    .A2(_17936_),
    .B1(_07462_),
    .B2(_17939_),
    .C1(_17980_),
    .Y(_17981_));
 sky130_fd_sc_hd__nand2_1 _39885_ (.A(_17981_),
    .B(_17947_),
    .Y(_17982_));
 sky130_fd_sc_hd__o21ai_0 _39886_ (.A1(\inst$top.soc.gpio_0._gpio.w_data$53 ),
    .A2(net844),
    .B1(net2167),
    .Y(_17983_));
 sky130_fd_sc_hd__a21oi_1 _39887_ (.A1(net844),
    .A2(_17982_),
    .B1(_17983_),
    .Y(_05097_));
 sky130_fd_sc_hd__inv_1 _39888_ (.A(_17871_),
    .Y(_17984_));
 sky130_fd_sc_hd__o21ai_0 _39889_ (.A1(_17849_),
    .A2(_17874_),
    .B1(_17984_),
    .Y(_17985_));
 sky130_fd_sc_hd__nand3_1 _39890_ (.A(_17845_),
    .B(_17866_),
    .C(_17985_),
    .Y(_17986_));
 sky130_fd_sc_hd__inv_1 _39891_ (.A(_17986_),
    .Y(_17987_));
 sky130_fd_sc_hd__o21ai_0 _39893_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__0.port__w_data ),
    .A2(net843),
    .B1(net2169),
    .Y(_17989_));
 sky130_fd_sc_hd__a21oi_1 _39894_ (.A1(net900),
    .A2(net843),
    .B1(_17989_),
    .Y(_05098_));
 sky130_fd_sc_hd__o21ai_0 _39895_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__1.port__w_data ),
    .A2(net843),
    .B1(net2168),
    .Y(_17990_));
 sky130_fd_sc_hd__a21oi_1 _39896_ (.A1(net868),
    .A2(net843),
    .B1(_17990_),
    .Y(_05099_));
 sky130_fd_sc_hd__o21ai_0 _39897_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__2.port__w_data ),
    .A2(net842),
    .B1(net2163),
    .Y(_17991_));
 sky130_fd_sc_hd__a21oi_1 _39898_ (.A1(_17954_),
    .A2(net842),
    .B1(_17991_),
    .Y(_05100_));
 sky130_fd_sc_hd__o21ai_0 _39899_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__3.port__w_data ),
    .A2(net842),
    .B1(net2167),
    .Y(_17992_));
 sky130_fd_sc_hd__a21oi_1 _39900_ (.A1(_17960_),
    .A2(net842),
    .B1(_17992_),
    .Y(_05101_));
 sky130_fd_sc_hd__o21ai_0 _39901_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__4.port__w_data ),
    .A2(net842),
    .B1(net2169),
    .Y(_17993_));
 sky130_fd_sc_hd__a21oi_1 _39902_ (.A1(net867),
    .A2(net843),
    .B1(_17993_),
    .Y(_05102_));
 sky130_fd_sc_hd__o21ai_0 _39904_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__5.port__w_data ),
    .A2(net842),
    .B1(net2167),
    .Y(_17995_));
 sky130_fd_sc_hd__a21oi_1 _39905_ (.A1(_17972_),
    .A2(net842),
    .B1(_17995_),
    .Y(_05103_));
 sky130_fd_sc_hd__o21ai_0 _39906_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__6.port__w_data ),
    .A2(net842),
    .B1(net2169),
    .Y(_17996_));
 sky130_fd_sc_hd__a21oi_1 _39907_ (.A1(_17977_),
    .A2(net843),
    .B1(_17996_),
    .Y(_05104_));
 sky130_fd_sc_hd__o21ai_0 _39908_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__7.port__w_data ),
    .A2(net842),
    .B1(net2168),
    .Y(_17997_));
 sky130_fd_sc_hd__a21oi_1 _39909_ (.A1(_17982_),
    .A2(net842),
    .B1(_17997_),
    .Y(_05105_));
 sky130_fd_sc_hd__inv_1 _39910_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__0.port__w_data ),
    .Y(_17998_));
 sky130_fd_sc_hd__o21ai_0 _39912_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__0._storage[0] ),
    .A2(net2582),
    .B1(net2165),
    .Y(_18000_));
 sky130_fd_sc_hd__a21oi_1 _39913_ (.A1(_17998_),
    .A2(net2582),
    .B1(_18000_),
    .Y(_05106_));
 sky130_fd_sc_hd__inv_1 _39914_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__1.port__w_data ),
    .Y(_18001_));
 sky130_fd_sc_hd__o21ai_0 _39915_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__0._storage[1] ),
    .A2(net2582),
    .B1(net2165),
    .Y(_18002_));
 sky130_fd_sc_hd__a21oi_1 _39916_ (.A1(_18001_),
    .A2(net2582),
    .B1(_18002_),
    .Y(_05107_));
 sky130_fd_sc_hd__inv_1 _39917_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__2.port__w_data ),
    .Y(_18003_));
 sky130_fd_sc_hd__o21ai_0 _39918_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__1._storage[0] ),
    .A2(net2582),
    .B1(net2165),
    .Y(_18004_));
 sky130_fd_sc_hd__a21oi_1 _39919_ (.A1(_18003_),
    .A2(net2582),
    .B1(_18004_),
    .Y(_05108_));
 sky130_fd_sc_hd__inv_1 _39920_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__3.port__w_data ),
    .Y(_18005_));
 sky130_fd_sc_hd__o21ai_0 _39921_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__1._storage[1] ),
    .A2(net2582),
    .B1(net2164),
    .Y(_18006_));
 sky130_fd_sc_hd__a21oi_1 _39922_ (.A1(_18005_),
    .A2(net2582),
    .B1(_18006_),
    .Y(_05109_));
 sky130_fd_sc_hd__inv_1 _39923_ (.A(\inst$top.soc.gpio_open_drain._gpio.w_data$38 ),
    .Y(_18007_));
 sky130_fd_sc_hd__o21ai_0 _39924_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__2._storage[0] ),
    .A2(net2582),
    .B1(net2164),
    .Y(_18008_));
 sky130_fd_sc_hd__a21oi_1 _39925_ (.A1(_18007_),
    .A2(net2583),
    .B1(_18008_),
    .Y(_05110_));
 sky130_fd_sc_hd__inv_1 _39926_ (.A(\inst$top.soc.gpio_open_drain._gpio.w_data$41 ),
    .Y(_18009_));
 sky130_fd_sc_hd__o21ai_0 _39927_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__2._storage[1] ),
    .A2(net2582),
    .B1(net2164),
    .Y(_18010_));
 sky130_fd_sc_hd__a21oi_1 _39928_ (.A1(_18009_),
    .A2(net2583),
    .B1(_18010_),
    .Y(_05111_));
 sky130_fd_sc_hd__inv_1 _39929_ (.A(\inst$top.soc.gpio_open_drain._gpio.w_data$50 ),
    .Y(_18011_));
 sky130_fd_sc_hd__o21ai_0 _39930_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__3._storage[0] ),
    .A2(net2583),
    .B1(net2164),
    .Y(_18012_));
 sky130_fd_sc_hd__a21oi_1 _39931_ (.A1(_18011_),
    .A2(net2583),
    .B1(_18012_),
    .Y(_05112_));
 sky130_fd_sc_hd__inv_1 _39932_ (.A(\inst$top.soc.gpio_open_drain._gpio.w_data$53 ),
    .Y(_18013_));
 sky130_fd_sc_hd__o21ai_0 _39934_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__3._storage[1] ),
    .A2(net2583),
    .B1(net2165),
    .Y(_18015_));
 sky130_fd_sc_hd__a21oi_1 _39935_ (.A1(_18013_),
    .A2(net2583),
    .B1(_18015_),
    .Y(_05113_));
 sky130_fd_sc_hd__nand2_1 _39936_ (.A(_17998_),
    .B(_18001_),
    .Y(_18016_));
 sky130_fd_sc_hd__nand2_1 _39937_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__0.port__w_data ),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__1.port__w_data ),
    .Y(_18017_));
 sky130_fd_sc_hd__a31oi_1 _39938_ (.A1(_18016_),
    .A2(_18017_),
    .A3(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$15 ),
    .B1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$14 ),
    .Y(_18018_));
 sky130_fd_sc_hd__inv_1 _39939_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__0._storage ),
    .Y(_18019_));
 sky130_fd_sc_hd__nor2_1 _39940_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__0.port__w_data ),
    .B(_18018_),
    .Y(_18020_));
 sky130_fd_sc_hd__a211oi_1 _39941_ (.A1(_18018_),
    .A2(_18019_),
    .B1(net3000),
    .C1(_18020_),
    .Y(_05114_));
 sky130_fd_sc_hd__inv_1 _39942_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__1._storage ),
    .Y(_18021_));
 sky130_fd_sc_hd__nand2_1 _39943_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__1.port__w_data ),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$14 ),
    .Y(_18022_));
 sky130_fd_sc_hd__o21ai_0 _39944_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$14 ),
    .A2(_18021_),
    .B1(_18022_),
    .Y(_18023_));
 sky130_fd_sc_hd__a31oi_1 _39945_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$15 ),
    .A2(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__2.port__w_data ),
    .A3(_18005_),
    .B1(_18023_),
    .Y(_18024_));
 sky130_fd_sc_hd__a311oi_1 _39946_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$15 ),
    .A2(_18003_),
    .A3(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__3.port__w_data ),
    .B1(net3000),
    .C1(_18024_),
    .Y(_05115_));
 sky130_fd_sc_hd__inv_1 _39947_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__2._storage ),
    .Y(_18025_));
 sky130_fd_sc_hd__nand2_1 _39948_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$14 ),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__2.port__w_data ),
    .Y(_18026_));
 sky130_fd_sc_hd__o21ai_0 _39949_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$14 ),
    .A2(_18025_),
    .B1(_18026_),
    .Y(_18027_));
 sky130_fd_sc_hd__a31oi_1 _39950_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$15 ),
    .A2(\inst$top.soc.gpio_open_drain._gpio.w_data$38 ),
    .A3(_18009_),
    .B1(_18027_),
    .Y(_18028_));
 sky130_fd_sc_hd__a311oi_1 _39951_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$15 ),
    .A2(_18007_),
    .A3(\inst$top.soc.gpio_open_drain._gpio.w_data$41 ),
    .B1(net3000),
    .C1(_18028_),
    .Y(_05116_));
 sky130_fd_sc_hd__inv_1 _39952_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__3._storage ),
    .Y(_18029_));
 sky130_fd_sc_hd__nand2_1 _39953_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$14 ),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__3.port__w_data ),
    .Y(_18030_));
 sky130_fd_sc_hd__o21ai_0 _39954_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$14 ),
    .A2(_18029_),
    .B1(_18030_),
    .Y(_18031_));
 sky130_fd_sc_hd__a31oi_1 _39955_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$15 ),
    .A2(\inst$top.soc.gpio_open_drain._gpio.w_data$50 ),
    .A3(_18013_),
    .B1(_18031_),
    .Y(_18032_));
 sky130_fd_sc_hd__a311oi_1 _39956_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$15 ),
    .A2(_18011_),
    .A3(\inst$top.soc.gpio_open_drain._gpio.w_data$53 ),
    .B1(net3000),
    .C1(_18032_),
    .Y(_05117_));
 sky130_fd_sc_hd__inv_1 _39957_ (.A(_09261_),
    .Y(_18033_));
 sky130_fd_sc_hd__nand3_1 _39958_ (.A(_17835_),
    .B(_18033_),
    .C(_09259_),
    .Y(_18034_));
 sky130_fd_sc_hd__inv_1 _39959_ (.A(_09269_),
    .Y(_18035_));
 sky130_fd_sc_hd__inv_1 _39960_ (.A(_09318_),
    .Y(_18036_));
 sky130_fd_sc_hd__nor4_1 _39961_ (.A(\inst$top.soc.bus__adr[2] ),
    .B(_18035_),
    .C(_18036_),
    .D(_09333_),
    .Y(_18037_));
 sky130_fd_sc_hd__nor2_1 _39962_ (.A(_17838_),
    .B(_17842_),
    .Y(_18038_));
 sky130_fd_sc_hd__nor3_1 _39963_ (.A(\inst$top.soc.bus__adr[7] ),
    .B(_09321_),
    .C(_09324_),
    .Y(_18039_));
 sky130_fd_sc_hd__nand4_1 _39964_ (.A(_18037_),
    .B(_09295_),
    .C(_18038_),
    .D(_18039_),
    .Y(_18040_));
 sky130_fd_sc_hd__nor2_1 _39965_ (.A(_18034_),
    .B(_18040_),
    .Y(_18041_));
 sky130_fd_sc_hd__nand2_1 _39966_ (.A(_18041_),
    .B(_17866_),
    .Y(_18042_));
 sky130_fd_sc_hd__nor3_2 _39967_ (.A(net2989),
    .B(_17880_),
    .C(_18042_),
    .Y(_05118_));
 sky130_fd_sc_hd__nor2_1 _39968_ (.A(_17833_),
    .B(_18042_),
    .Y(_05119_));
 sky130_fd_sc_hd__nor2_1 _39969_ (.A(net2989),
    .B(_17887_),
    .Y(_18043_));
 sky130_fd_sc_hd__clkinv_1 _39970_ (.A(_18043_),
    .Y(_18044_));
 sky130_fd_sc_hd__nor2_1 _39971_ (.A(_18044_),
    .B(_18042_),
    .Y(_05120_));
 sky130_fd_sc_hd__nor4_4 _39972_ (.A(_17874_),
    .B(_17876_),
    .C(_18034_),
    .D(_18040_),
    .Y(_18045_));
 sky130_fd_sc_hd__nand2_1 _39973_ (.A(_18045_),
    .B(_17859_),
    .Y(_18046_));
 sky130_fd_sc_hd__nand3_1 _39974_ (.A(_18045_),
    .B(\inst$top.soc.gpio_open_drain._gpio.r_data ),
    .C(_17850_),
    .Y(_18047_));
 sky130_fd_sc_hd__nand2_1 _39975_ (.A(_18045_),
    .B(_17831_),
    .Y(_18048_));
 sky130_fd_sc_hd__a21oi_1 _39977_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__0._storage ),
    .A2(_17855_),
    .B1(_18048_),
    .Y(_18050_));
 sky130_fd_sc_hd__o211ai_1 _39978_ (.A1(_02887_),
    .A2(_18046_),
    .B1(_18047_),
    .C1(_18050_),
    .Y(_18051_));
 sky130_fd_sc_hd__inv_1 _39979_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[0] ),
    .Y(_18052_));
 sky130_fd_sc_hd__a21oi_1 _39980_ (.A1(net829),
    .A2(_18052_),
    .B1(net2999),
    .Y(_18053_));
 sky130_fd_sc_hd__nand2_1 _39981_ (.A(_18051_),
    .B(_18053_),
    .Y(_18054_));
 sky130_fd_sc_hd__inv_2 _39982_ (.A(_18054_),
    .Y(_05121_));
 sky130_fd_sc_hd__a21oi_1 _39983_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__1._storage ),
    .A2(_17855_),
    .B1(net829),
    .Y(_18055_));
 sky130_fd_sc_hd__nand3_1 _39984_ (.A(_18045_),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__0._storage[1] ),
    .C(_17859_),
    .Y(_18056_));
 sky130_fd_sc_hd__nand3_1 _39985_ (.A(_18045_),
    .B(\inst$top.soc.gpio_open_drain._gpio.r_data$23 ),
    .C(_17850_),
    .Y(_18057_));
 sky130_fd_sc_hd__a21oi_1 _39986_ (.A1(_18045_),
    .A2(_17831_),
    .B1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[1] ),
    .Y(_18058_));
 sky130_fd_sc_hd__a311o_1 _39987_ (.A1(_18055_),
    .A2(_18056_),
    .A3(_18057_),
    .B1(net3000),
    .C1(_18058_),
    .X(_18059_));
 sky130_fd_sc_hd__inv_2 _39988_ (.A(_18059_),
    .Y(_05122_));
 sky130_fd_sc_hd__nand3_1 _39989_ (.A(_18045_),
    .B(\inst$top.soc.gpio_open_drain._gpio.r_data$35 ),
    .C(_17850_),
    .Y(_18060_));
 sky130_fd_sc_hd__a21oi_1 _39990_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__2._storage ),
    .A2(_17855_),
    .B1(net829),
    .Y(_18061_));
 sky130_fd_sc_hd__o211ai_1 _39991_ (.A1(_02884_),
    .A2(_18046_),
    .B1(_18060_),
    .C1(_18061_),
    .Y(_18062_));
 sky130_fd_sc_hd__inv_1 _39992_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[2] ),
    .Y(_18063_));
 sky130_fd_sc_hd__a21oi_1 _39993_ (.A1(net829),
    .A2(_18063_),
    .B1(net2999),
    .Y(_18064_));
 sky130_fd_sc_hd__nand2_1 _39994_ (.A(_18062_),
    .B(_18064_),
    .Y(_18065_));
 sky130_fd_sc_hd__inv_2 _39995_ (.A(_18065_),
    .Y(_05123_));
 sky130_fd_sc_hd__a21oi_1 _39996_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__3._storage ),
    .A2(_17855_),
    .B1(net829),
    .Y(_18066_));
 sky130_fd_sc_hd__nand3_1 _39997_ (.A(_18045_),
    .B(\inst$top.soc.gpio_open_drain._gpio.r_data$47 ),
    .C(_17850_),
    .Y(_18067_));
 sky130_fd_sc_hd__nand3_1 _39998_ (.A(_18045_),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__1._storage[1] ),
    .C(_17859_),
    .Y(_18068_));
 sky130_fd_sc_hd__a21oi_1 _39999_ (.A1(_18045_),
    .A2(_17831_),
    .B1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[3] ),
    .Y(_18069_));
 sky130_fd_sc_hd__a311o_1 _40000_ (.A1(_18066_),
    .A2(_18067_),
    .A3(_18068_),
    .B1(net3000),
    .C1(_18069_),
    .X(_18070_));
 sky130_fd_sc_hd__inv_2 _40001_ (.A(_18070_),
    .Y(_05124_));
 sky130_fd_sc_hd__nand2_1 _40002_ (.A(net829),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[4] ),
    .Y(_18071_));
 sky130_fd_sc_hd__nand4_1 _40003_ (.A(_17835_),
    .B(_09269_),
    .C(_18033_),
    .D(_09259_),
    .Y(_18072_));
 sky130_fd_sc_hd__nor4_2 _40004_ (.A(_17887_),
    .B(_18072_),
    .C(_17876_),
    .D(_17844_),
    .Y(_18073_));
 sky130_fd_sc_hd__nand2_1 _40005_ (.A(net841),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__2._storage[0] ),
    .Y(_18074_));
 sky130_fd_sc_hd__a21oi_2 _40006_ (.A1(_18071_),
    .A2(_18074_),
    .B1(net2999),
    .Y(_05125_));
 sky130_fd_sc_hd__nand2_1 _40007_ (.A(net829),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[5] ),
    .Y(_18075_));
 sky130_fd_sc_hd__nand2_1 _40008_ (.A(net841),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__2._storage[1] ),
    .Y(_18076_));
 sky130_fd_sc_hd__a21oi_2 _40009_ (.A1(_18075_),
    .A2(_18076_),
    .B1(net2999),
    .Y(_05126_));
 sky130_fd_sc_hd__nand2_1 _40010_ (.A(net829),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[6] ),
    .Y(_18077_));
 sky130_fd_sc_hd__nand2_1 _40011_ (.A(net841),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__3._storage[0] ),
    .Y(_18078_));
 sky130_fd_sc_hd__a21oi_2 _40013_ (.A1(_18077_),
    .A2(_18078_),
    .B1(net3000),
    .Y(_05127_));
 sky130_fd_sc_hd__nand2_1 _40014_ (.A(net829),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[7] ),
    .Y(_18080_));
 sky130_fd_sc_hd__nand2_1 _40015_ (.A(net841),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__3._storage[1] ),
    .Y(_18081_));
 sky130_fd_sc_hd__a21oi_2 _40016_ (.A1(_18080_),
    .A2(_18081_),
    .B1(net3000),
    .Y(_05128_));
 sky130_fd_sc_hd__nor2_2 _40017_ (.A(net2999),
    .B(net829),
    .Y(_05129_));
 sky130_fd_sc_hd__nor3_1 _40018_ (.A(_17850_),
    .B(_17874_),
    .C(_18042_),
    .Y(_18082_));
 sky130_fd_sc_hd__o21ai_0 _40020_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__0.port__w_data ),
    .A2(net839),
    .B1(net2165),
    .Y(_18084_));
 sky130_fd_sc_hd__a21oi_2 _40021_ (.A1(net900),
    .A2(net839),
    .B1(_18084_),
    .Y(_05130_));
 sky130_fd_sc_hd__o21ai_0 _40022_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__1.port__w_data ),
    .A2(net839),
    .B1(net2164),
    .Y(_18085_));
 sky130_fd_sc_hd__a21oi_2 _40023_ (.A1(net868),
    .A2(net839),
    .B1(_18085_),
    .Y(_05131_));
 sky130_fd_sc_hd__o21ai_0 _40024_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__2.port__w_data ),
    .A2(net839),
    .B1(net2166),
    .Y(_18086_));
 sky130_fd_sc_hd__a21oi_2 _40025_ (.A1(_17954_),
    .A2(net839),
    .B1(_18086_),
    .Y(_05132_));
 sky130_fd_sc_hd__o21ai_0 _40026_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__3.port__w_data ),
    .A2(net839),
    .B1(net2164),
    .Y(_18087_));
 sky130_fd_sc_hd__a21oi_2 _40027_ (.A1(_17960_),
    .A2(net839),
    .B1(_18087_),
    .Y(_05133_));
 sky130_fd_sc_hd__o21ai_0 _40028_ (.A1(\inst$top.soc.gpio_open_drain._gpio.w_data$38 ),
    .A2(net839),
    .B1(net2164),
    .Y(_18088_));
 sky130_fd_sc_hd__a21oi_1 _40029_ (.A1(net867),
    .A2(net840),
    .B1(_18088_),
    .Y(_05134_));
 sky130_fd_sc_hd__inv_1 _40030_ (.A(net839),
    .Y(_18089_));
 sky130_fd_sc_hd__inv_1 _40031_ (.A(_17972_),
    .Y(_18090_));
 sky130_fd_sc_hd__o21ai_0 _40032_ (.A1(_18090_),
    .A2(_18089_),
    .B1(net2164),
    .Y(_18091_));
 sky130_fd_sc_hd__a21oi_2 _40033_ (.A1(_18009_),
    .A2(_18089_),
    .B1(_18091_),
    .Y(_05135_));
 sky130_fd_sc_hd__o21ai_0 _40034_ (.A1(\inst$top.soc.gpio_open_drain._gpio.w_data$50 ),
    .A2(net840),
    .B1(net2164),
    .Y(_18092_));
 sky130_fd_sc_hd__a21oi_1 _40035_ (.A1(_17977_),
    .A2(net840),
    .B1(_18092_),
    .Y(_05136_));
 sky130_fd_sc_hd__inv_1 _40036_ (.A(_17982_),
    .Y(_18093_));
 sky130_fd_sc_hd__o21ai_0 _40037_ (.A1(_18093_),
    .A2(_18089_),
    .B1(net2164),
    .Y(_18094_));
 sky130_fd_sc_hd__a21oi_2 _40038_ (.A1(_18013_),
    .A2(_18089_),
    .B1(_18094_),
    .Y(_05137_));
 sky130_fd_sc_hd__nor2_1 _40039_ (.A(_17885_),
    .B(_17870_),
    .Y(_18095_));
 sky130_fd_sc_hd__clkinv_1 _40040_ (.A(_18095_),
    .Y(_18096_));
 sky130_fd_sc_hd__nor2_1 _40041_ (.A(_09270_),
    .B(_17844_),
    .Y(_18097_));
 sky130_fd_sc_hd__nand2_1 _40042_ (.A(_18097_),
    .B(_09301_),
    .Y(_18098_));
 sky130_fd_sc_hd__inv_1 _40043_ (.A(_18098_),
    .Y(_18099_));
 sky130_fd_sc_hd__inv_1 _40044_ (.A(_09273_),
    .Y(_18100_));
 sky130_fd_sc_hd__nor2_1 _40045_ (.A(_09276_),
    .B(_18100_),
    .Y(_18101_));
 sky130_fd_sc_hd__nand3_1 _40046_ (.A(_18099_),
    .B(_17882_),
    .C(_18101_),
    .Y(_18102_));
 sky130_fd_sc_hd__nand4_1 _40047_ (.A(_18099_),
    .B(_17882_),
    .C(_17931_),
    .D(_18101_),
    .Y(_18103_));
 sky130_fd_sc_hd__nand3_1 _40048_ (.A(_18103_),
    .B(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[6] ),
    .C(net2140),
    .Y(_18104_));
 sky130_fd_sc_hd__o31ai_2 _40049_ (.A1(net2984),
    .A2(_18096_),
    .A3(_18102_),
    .B1(_18104_),
    .Y(_05138_));
 sky130_fd_sc_hd__nor2_1 _40050_ (.A(net2984),
    .B(_18103_),
    .Y(_05139_));
 sky130_fd_sc_hd__a21oi_1 _40051_ (.A1(_17872_),
    .A2(_17873_),
    .B1(_18102_),
    .Y(_05140_));
 sky130_fd_sc_hd__nand3_1 _40052_ (.A(_18103_),
    .B(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[1] ),
    .C(net2137),
    .Y(_18105_));
 sky130_fd_sc_hd__o21ai_1 _40053_ (.A1(_18044_),
    .A2(_18102_),
    .B1(_18105_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand2_1 _40054_ (.A(net2132),
    .B(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[0] ),
    .Y(_18106_));
 sky130_fd_sc_hd__o21ai_1 _40055_ (.A1(net2984),
    .A2(_18103_),
    .B1(_18106_),
    .Y(_05142_));
 sky130_fd_sc_hd__nor4_2 _40056_ (.A(net2979),
    .B(\inst$top.soc.bus__addr[3] ),
    .C(_17856_),
    .D(_18102_),
    .Y(_05143_));
 sky130_fd_sc_hd__nor4_2 _40057_ (.A(net2979),
    .B(\inst$top.soc.bus__addr[3] ),
    .C(_17831_),
    .D(_18102_),
    .Y(_05144_));
 sky130_fd_sc_hd__inv_1 _40058_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[3] ),
    .Y(_18107_));
 sky130_fd_sc_hd__o21ai_0 _40059_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[0] ),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb ),
    .B1(net2126),
    .Y(_18108_));
 sky130_fd_sc_hd__a21oi_1 _40060_ (.A1(_18107_),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb ),
    .B1(_18108_),
    .Y(_05145_));
 sky130_fd_sc_hd__inv_1 _40061_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[4] ),
    .Y(_18109_));
 sky130_fd_sc_hd__o21ai_0 _40063_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[1] ),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb ),
    .B1(net2128),
    .Y(_18111_));
 sky130_fd_sc_hd__a21oi_1 _40064_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb ),
    .A2(_18109_),
    .B1(_18111_),
    .Y(_05146_));
 sky130_fd_sc_hd__inv_1 _40065_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.port__w_data ),
    .Y(_18112_));
 sky130_fd_sc_hd__o21ai_0 _40066_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.raw_enable._storage ),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb ),
    .B1(net2129),
    .Y(_18113_));
 sky130_fd_sc_hd__a21oi_1 _40067_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb ),
    .A2(_18112_),
    .B1(_18113_),
    .Y(_05147_));
 sky130_fd_sc_hd__inv_1 _40068_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.RawControl.port__w_data ),
    .Y(_18114_));
 sky130_fd_sc_hd__o21ai_0 _40069_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[0] ),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb ),
    .B1(net2063),
    .Y(_18115_));
 sky130_fd_sc_hd__a21oi_1 _40070_ (.A1(_18114_),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb ),
    .B1(_18115_),
    .Y(_05148_));
 sky130_fd_sc_hd__inv_1 _40071_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[2] ),
    .Y(_18116_));
 sky130_fd_sc_hd__o21ai_0 _40072_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[1] ),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb ),
    .B1(net2063),
    .Y(_18117_));
 sky130_fd_sc_hd__a21oi_1 _40073_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb ),
    .A2(_18116_),
    .B1(_18117_),
    .Y(_05149_));
 sky130_fd_sc_hd__o21ai_0 _40075_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[0] ),
    .A2(net2581),
    .B1(net2129),
    .Y(_18119_));
 sky130_fd_sc_hd__a21oi_1 _40076_ (.A1(_18112_),
    .A2(net2581),
    .B1(_18119_),
    .Y(_05150_));
 sky130_fd_sc_hd__o21ai_0 _40077_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[1] ),
    .A2(net2580),
    .B1(net2061),
    .Y(_18120_));
 sky130_fd_sc_hd__a21oi_1 _40078_ (.A1(_18114_),
    .A2(net2580),
    .B1(_18120_),
    .Y(_05151_));
 sky130_fd_sc_hd__o21ai_0 _40079_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[2] ),
    .A2(net2580),
    .B1(net2061),
    .Y(_18121_));
 sky130_fd_sc_hd__a21oi_1 _40080_ (.A1(_18116_),
    .A2(net2580),
    .B1(_18121_),
    .Y(_05152_));
 sky130_fd_sc_hd__o21ai_0 _40081_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[3] ),
    .A2(net2580),
    .B1(net2126),
    .Y(_18122_));
 sky130_fd_sc_hd__a21oi_1 _40082_ (.A1(_18107_),
    .A2(net2580),
    .B1(_18122_),
    .Y(_05153_));
 sky130_fd_sc_hd__o21ai_0 _40083_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[4] ),
    .A2(net2580),
    .B1(net2126),
    .Y(_18123_));
 sky130_fd_sc_hd__a21oi_1 _40084_ (.A1(_18109_),
    .A2(net2581),
    .B1(_18123_),
    .Y(_05154_));
 sky130_fd_sc_hd__inv_1 _40085_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[5] ),
    .Y(_18124_));
 sky130_fd_sc_hd__o21ai_0 _40086_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[5] ),
    .A2(net2580),
    .B1(net2129),
    .Y(_18125_));
 sky130_fd_sc_hd__a21oi_1 _40087_ (.A1(net2581),
    .A2(_18124_),
    .B1(_18125_),
    .Y(_05155_));
 sky130_fd_sc_hd__inv_1 _40088_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[6] ),
    .Y(_18126_));
 sky130_fd_sc_hd__o21ai_0 _40090_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[6] ),
    .A2(net2580),
    .B1(net2128),
    .Y(_18128_));
 sky130_fd_sc_hd__a21oi_1 _40091_ (.A1(net2581),
    .A2(_18126_),
    .B1(_18128_),
    .Y(_05156_));
 sky130_fd_sc_hd__inv_1 _40092_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[7] ),
    .Y(_18129_));
 sky130_fd_sc_hd__o21ai_0 _40093_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[7] ),
    .A2(net2581),
    .B1(net2131),
    .Y(_18130_));
 sky130_fd_sc_hd__a21oi_1 _40094_ (.A1(net2581),
    .A2(_18129_),
    .B1(_18130_),
    .Y(_05157_));
 sky130_fd_sc_hd__inv_1 _40096_ (.A(net2580),
    .Y(_18132_));
 sky130_fd_sc_hd__nor2_1 _40097_ (.A(net2948),
    .B(_18132_),
    .Y(_05158_));
 sky130_fd_sc_hd__nor2_2 _40098_ (.A(_09277_),
    .B(_18098_),
    .Y(_18133_));
 sky130_fd_sc_hd__nand2_1 _40099_ (.A(_18133_),
    .B(_17866_),
    .Y(_18134_));
 sky130_fd_sc_hd__nor3_2 _40100_ (.A(net2983),
    .B(_18096_),
    .C(_18134_),
    .Y(_05159_));
 sky130_fd_sc_hd__nor2_1 _40101_ (.A(\inst$top.soc.bus__addr[2] ),
    .B(_19850_),
    .Y(_18135_));
 sky130_fd_sc_hd__inv_1 _40102_ (.A(_18135_),
    .Y(_18136_));
 sky130_fd_sc_hd__nor2_1 _40103_ (.A(_17885_),
    .B(_18136_),
    .Y(_18137_));
 sky130_fd_sc_hd__inv_1 _40104_ (.A(_18137_),
    .Y(_18138_));
 sky130_fd_sc_hd__nor3_2 _40105_ (.A(net2983),
    .B(_18138_),
    .C(_18134_),
    .Y(_05160_));
 sky130_fd_sc_hd__nor2_1 _40106_ (.A(_18044_),
    .B(_18134_),
    .Y(_05161_));
 sky130_fd_sc_hd__nor2_1 _40107_ (.A(\inst$top.soc.spiflash.ctrl.fsm_state[3] ),
    .B(\inst$top.soc.spiflash.ctrl.fsm_state[2] ),
    .Y(_18139_));
 sky130_fd_sc_hd__inv_1 _40108_ (.A(_18139_),
    .Y(_18140_));
 sky130_fd_sc_hd__inv_1 _40109_ (.A(\inst$top.soc.spiflash.ctrl.fsm_state[0] ),
    .Y(_18141_));
 sky130_fd_sc_hd__nor2_1 _40110_ (.A(\inst$top.soc.spiflash.ctrl.fsm_state[1] ),
    .B(_18141_),
    .Y(_18142_));
 sky130_fd_sc_hd__inv_1 _40111_ (.A(_18142_),
    .Y(_18143_));
 sky130_fd_sc_hd__nor2_1 _40112_ (.A(_18140_),
    .B(_18143_),
    .Y(_18144_));
 sky130_fd_sc_hd__nand4_1 _40113_ (.A(_18133_),
    .B(_17882_),
    .C(_18095_),
    .D(_18144_),
    .Y(_18145_));
 sky130_fd_sc_hd__nand2_1 _40114_ (.A(_18133_),
    .B(_17882_),
    .Y(_18146_));
 sky130_fd_sc_hd__nor2_1 _40115_ (.A(_17885_),
    .B(_18146_),
    .Y(_18147_));
 sky130_fd_sc_hd__nor2_1 _40117_ (.A(_17868_),
    .B(_19850_),
    .Y(_18149_));
 sky130_fd_sc_hd__inv_1 _40118_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.raw_enable._storage ),
    .Y(_18150_));
 sky130_fd_sc_hd__nor2_1 _40119_ (.A(_18150_),
    .B(_17874_),
    .Y(_18151_));
 sky130_fd_sc_hd__a221oi_1 _40120_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[0] ),
    .A2(_18135_),
    .B1(\inst$top.soc.spiflash.ctrl.r_data[0] ),
    .B2(_18149_),
    .C1(_18151_),
    .Y(_18152_));
 sky130_fd_sc_hd__o21ai_0 _40121_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[0] ),
    .A2(net808),
    .B1(net2129),
    .Y(_18153_));
 sky130_fd_sc_hd__a31oi_1 _40122_ (.A1(_18145_),
    .A2(net809),
    .A3(_18152_),
    .B1(_18153_),
    .Y(_05162_));
 sky130_fd_sc_hd__nand2_1 _40123_ (.A(_17830_),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[0] ),
    .Y(_18154_));
 sky130_fd_sc_hd__nand2_1 _40124_ (.A(_18135_),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[1] ),
    .Y(_18155_));
 sky130_fd_sc_hd__nand2_1 _40125_ (.A(_18149_),
    .B(\inst$top.soc.spiflash.ctrl.r_data[1] ),
    .Y(_18156_));
 sky130_fd_sc_hd__o21ai_0 _40126_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[1] ),
    .A2(net808),
    .B1(net2126),
    .Y(_18157_));
 sky130_fd_sc_hd__a41oi_1 _40127_ (.A1(net808),
    .A2(_18154_),
    .A3(_18155_),
    .A4(_18156_),
    .B1(_18157_),
    .Y(_05163_));
 sky130_fd_sc_hd__nand2_1 _40128_ (.A(_17830_),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[1] ),
    .Y(_18158_));
 sky130_fd_sc_hd__nand2_1 _40129_ (.A(_18135_),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[2] ),
    .Y(_18159_));
 sky130_fd_sc_hd__nand2_1 _40130_ (.A(_18149_),
    .B(\inst$top.soc.spiflash.ctrl.r_data[2] ),
    .Y(_18160_));
 sky130_fd_sc_hd__o21ai_0 _40131_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[2] ),
    .A2(net808),
    .B1(net2119),
    .Y(_18161_));
 sky130_fd_sc_hd__a41oi_2 _40132_ (.A1(net808),
    .A2(_18158_),
    .A3(_18159_),
    .A4(_18160_),
    .B1(_18161_),
    .Y(_05164_));
 sky130_fd_sc_hd__nand2_1 _40133_ (.A(_17830_),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[0] ),
    .Y(_18162_));
 sky130_fd_sc_hd__nand2_1 _40134_ (.A(_18135_),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[3] ),
    .Y(_18163_));
 sky130_fd_sc_hd__nand2_1 _40135_ (.A(_18149_),
    .B(\inst$top.soc.spiflash.ctrl.r_data[3] ),
    .Y(_18164_));
 sky130_fd_sc_hd__o21ai_0 _40136_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[3] ),
    .A2(net808),
    .B1(net2126),
    .Y(_18165_));
 sky130_fd_sc_hd__a41oi_2 _40137_ (.A1(net808),
    .A2(_18162_),
    .A3(_18163_),
    .A4(_18164_),
    .B1(_18165_),
    .Y(_05165_));
 sky130_fd_sc_hd__inv_1 _40138_ (.A(net808),
    .Y(_18166_));
 sky130_fd_sc_hd__a221oi_1 _40139_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[4] ),
    .A2(_18135_),
    .B1(\inst$top.soc.spiflash.ctrl.r_data[4] ),
    .B2(_18149_),
    .C1(_18166_),
    .Y(_18167_));
 sky130_fd_sc_hd__nand4_1 _40140_ (.A(_18133_),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[1] ),
    .C(_17882_),
    .D(_17886_),
    .Y(_18168_));
 sky130_fd_sc_hd__o21ai_0 _40141_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[4] ),
    .A2(net809),
    .B1(net2131),
    .Y(_18169_));
 sky130_fd_sc_hd__a21oi_2 _40142_ (.A1(_18167_),
    .A2(_18168_),
    .B1(_18169_),
    .Y(_05166_));
 sky130_fd_sc_hd__a21oi_1 _40143_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[5] ),
    .A2(_18135_),
    .B1(_18166_),
    .Y(_18170_));
 sky130_fd_sc_hd__nand3_1 _40144_ (.A(net809),
    .B(\inst$top.soc.spiflash.ctrl.r_data[5] ),
    .C(_18149_),
    .Y(_18171_));
 sky130_fd_sc_hd__o21ai_0 _40145_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[5] ),
    .A2(net809),
    .B1(net2123),
    .Y(_18172_));
 sky130_fd_sc_hd__a21oi_2 _40146_ (.A1(_18170_),
    .A2(_18171_),
    .B1(_18172_),
    .Y(_05167_));
 sky130_fd_sc_hd__a21oi_1 _40147_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[6] ),
    .A2(_18135_),
    .B1(_18166_),
    .Y(_18173_));
 sky130_fd_sc_hd__nand3_1 _40148_ (.A(net808),
    .B(\inst$top.soc.spiflash.ctrl.r_data[6] ),
    .C(_18149_),
    .Y(_18174_));
 sky130_fd_sc_hd__o21ai_0 _40149_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[6] ),
    .A2(net808),
    .B1(net2119),
    .Y(_18175_));
 sky130_fd_sc_hd__a21oi_2 _40150_ (.A1(_18173_),
    .A2(_18174_),
    .B1(_18175_),
    .Y(_05168_));
 sky130_fd_sc_hd__a21oi_1 _40151_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[7] ),
    .A2(_18135_),
    .B1(_18166_),
    .Y(_18176_));
 sky130_fd_sc_hd__nand3_1 _40152_ (.A(net809),
    .B(\inst$top.soc.spiflash.ctrl.r_data[7] ),
    .C(_18149_),
    .Y(_18177_));
 sky130_fd_sc_hd__o21ai_0 _40153_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[7] ),
    .A2(net809),
    .B1(net2129),
    .Y(_18178_));
 sky130_fd_sc_hd__a21oi_2 _40154_ (.A1(_18176_),
    .A2(_18177_),
    .B1(_18178_),
    .Y(_05169_));
 sky130_fd_sc_hd__nor2_1 _40155_ (.A(net2981),
    .B(_18166_),
    .Y(_05170_));
 sky130_fd_sc_hd__nor2_1 _40156_ (.A(_17885_),
    .B(_18134_),
    .Y(_18179_));
 sky130_fd_sc_hd__o21ai_0 _40158_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.port__w_data ),
    .A2(_18179_),
    .B1(net2129),
    .Y(_18181_));
 sky130_fd_sc_hd__a21oi_2 _40159_ (.A1(_17941_),
    .A2(_18179_),
    .B1(_18181_),
    .Y(_05171_));
 sky130_fd_sc_hd__o21ai_0 _40160_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawControl.port__w_data ),
    .A2(net807),
    .B1(net2063),
    .Y(_18182_));
 sky130_fd_sc_hd__a21oi_2 _40161_ (.A1(_17948_),
    .A2(net807),
    .B1(_18182_),
    .Y(_05172_));
 sky130_fd_sc_hd__o21ai_0 _40162_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[2] ),
    .A2(net807),
    .B1(net2063),
    .Y(_18183_));
 sky130_fd_sc_hd__a21oi_2 _40163_ (.A1(_17954_),
    .A2(net807),
    .B1(_18183_),
    .Y(_05173_));
 sky130_fd_sc_hd__o21ai_0 _40164_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[3] ),
    .A2(net807),
    .B1(net2126),
    .Y(_18184_));
 sky130_fd_sc_hd__a21oi_2 _40165_ (.A1(_17960_),
    .A2(net807),
    .B1(_18184_),
    .Y(_05174_));
 sky130_fd_sc_hd__o21ai_0 _40167_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[4] ),
    .A2(net807),
    .B1(net2128),
    .Y(_18186_));
 sky130_fd_sc_hd__a21oi_1 _40168_ (.A1(_17967_),
    .A2(net807),
    .B1(_18186_),
    .Y(_05175_));
 sky130_fd_sc_hd__nor3_1 _40169_ (.A(_09256_),
    .B(_17862_),
    .C(_17865_),
    .Y(_18187_));
 sky130_fd_sc_hd__nand3_1 _40170_ (.A(_18133_),
    .B(_17859_),
    .C(_18187_),
    .Y(_18188_));
 sky130_fd_sc_hd__o21ai_0 _40171_ (.A1(_18090_),
    .A2(_18188_),
    .B1(net2123),
    .Y(_18189_));
 sky130_fd_sc_hd__a21oi_1 _40172_ (.A1(_18124_),
    .A2(_18188_),
    .B1(_18189_),
    .Y(_05176_));
 sky130_fd_sc_hd__o21ai_0 _40173_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[6] ),
    .A2(net807),
    .B1(net2119),
    .Y(_18190_));
 sky130_fd_sc_hd__a21oi_1 _40174_ (.A1(_17977_),
    .A2(net807),
    .B1(_18190_),
    .Y(_05177_));
 sky130_fd_sc_hd__o21ai_0 _40175_ (.A1(_18093_),
    .A2(_18188_),
    .B1(net2123),
    .Y(_18191_));
 sky130_fd_sc_hd__a21oi_1 _40176_ (.A1(_18129_),
    .A2(_18188_),
    .B1(_18191_),
    .Y(_05178_));
 sky130_fd_sc_hd__nor2_1 _40177_ (.A(\inst$top.soc.spiflash.ctrl.fsm_state[1] ),
    .B(\inst$top.soc.spiflash.ctrl.fsm_state[0] ),
    .Y(_18192_));
 sky130_fd_sc_hd__inv_1 _40178_ (.A(_18192_),
    .Y(_18193_));
 sky130_fd_sc_hd__nor2_1 _40179_ (.A(_18140_),
    .B(_18193_),
    .Y(_18194_));
 sky130_fd_sc_hd__inv_1 _40180_ (.A(_18194_),
    .Y(_18195_));
 sky130_fd_sc_hd__nor2_1 _40181_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.raw_enable._storage ),
    .B(_18195_),
    .Y(_18196_));
 sky130_fd_sc_hd__inv_2 _40182_ (.A(\inst$top.soc.spiflash.ctrl.fsm_state[2] ),
    .Y(_18197_));
 sky130_fd_sc_hd__nor2_1 _40183_ (.A(\inst$top.soc.spiflash.ctrl.fsm_state[3] ),
    .B(_18197_),
    .Y(_18198_));
 sky130_fd_sc_hd__inv_1 _40184_ (.A(_18198_),
    .Y(_18199_));
 sky130_fd_sc_hd__inv_1 _40185_ (.A(\inst$top.soc.spiflash.ctrl.fsm_state[1] ),
    .Y(_18200_));
 sky130_fd_sc_hd__nor2_1 _40186_ (.A(_18200_),
    .B(_18140_),
    .Y(_18201_));
 sky130_fd_sc_hd__inv_1 _40187_ (.A(_18201_),
    .Y(_18202_));
 sky130_fd_sc_hd__o21ai_0 _40188_ (.A1(_18199_),
    .A2(_18192_),
    .B1(_18202_),
    .Y(_18203_));
 sky130_fd_sc_hd__inv_1 _40189_ (.A(\inst$top.soc.spiflash.phy.enframer.cycle[2] ),
    .Y(_18204_));
 sky130_fd_sc_hd__nor2_1 _40190_ (.A(_18193_),
    .B(_18199_),
    .Y(_18205_));
 sky130_fd_sc_hd__nor2_1 _40191_ (.A(_18201_),
    .B(_18194_),
    .Y(_18206_));
 sky130_fd_sc_hd__nand2_1 _40192_ (.A(\inst$top.soc.spiflash.ctrl.fsm_state[1] ),
    .B(\inst$top.soc.spiflash.ctrl.fsm_state[0] ),
    .Y(_18207_));
 sky130_fd_sc_hd__nor2_1 _40193_ (.A(_18207_),
    .B(_18199_),
    .Y(_18208_));
 sky130_fd_sc_hd__inv_1 _40194_ (.A(_18208_),
    .Y(_18209_));
 sky130_fd_sc_hd__nand2_1 _40195_ (.A(_18206_),
    .B(_18209_),
    .Y(_18210_));
 sky130_fd_sc_hd__nor2_1 _40196_ (.A(_18205_),
    .B(_18210_),
    .Y(_18211_));
 sky130_fd_sc_hd__inv_1 _40197_ (.A(_18211_),
    .Y(_18212_));
 sky130_fd_sc_hd__a21oi_1 _40198_ (.A1(_18204_),
    .A2(_02746_),
    .B1(_18212_),
    .Y(_18213_));
 sky130_fd_sc_hd__inv_1 _40199_ (.A(\inst$top.soc.spiflash.phy.deframer.cycle[2] ),
    .Y(_18214_));
 sky130_fd_sc_hd__inv_2 _40200_ (.A(\inst$top.soc.spiflash.phy.io_streamer.skid_at ),
    .Y(_18215_));
 sky130_fd_sc_hd__nand2_1 _40201_ (.A(_18215_),
    .B(\inst$top.soc.spiflash.phy.io_streamer.meta_0[0] ),
    .Y(_18216_));
 sky130_fd_sc_hd__nand2_1 _40202_ (.A(\inst$top.soc.spiflash.phy.io_streamer.skid_at ),
    .B(\inst$top.soc.spiflash.phy.io_streamer.skid_1.meta[0] ),
    .Y(_18217_));
 sky130_fd_sc_hd__nand2_1 _40203_ (.A(_18216_),
    .B(_18217_),
    .Y(_18218_));
 sky130_fd_sc_hd__inv_1 _40204_ (.A(\inst$top.soc.spiflash.phy.io_streamer.skid_1.meta[2] ),
    .Y(_18219_));
 sky130_fd_sc_hd__nand2_1 _40205_ (.A(_18219_),
    .B(\inst$top.soc.spiflash.phy.io_streamer.skid_at ),
    .Y(_18220_));
 sky130_fd_sc_hd__o21ai_1 _40206_ (.A1(\inst$top.soc.spiflash.phy.io_streamer.skid_at ),
    .A2(\inst$top.soc.spiflash.phy.io_streamer.meta_0[2] ),
    .B1(_18220_),
    .Y(_18221_));
 sky130_fd_sc_hd__nor2_2 _40207_ (.A(_18218_),
    .B(_18221_),
    .Y(_18222_));
 sky130_fd_sc_hd__inv_1 _40208_ (.A(_18222_),
    .Y(_18223_));
 sky130_fd_sc_hd__nand2_1 _40209_ (.A(_18221_),
    .B(_18218_),
    .Y(_18224_));
 sky130_fd_sc_hd__inv_1 _40210_ (.A(\inst$top.soc.spiflash.phy.io_streamer.skid_1.meta[1] ),
    .Y(_18225_));
 sky130_fd_sc_hd__nand2_1 _40211_ (.A(_18215_),
    .B(\inst$top.soc.spiflash.phy.io_streamer.meta_0[1] ),
    .Y(_18226_));
 sky130_fd_sc_hd__o21ai_0 _40212_ (.A1(_18215_),
    .A2(_18225_),
    .B1(_18226_),
    .Y(_18227_));
 sky130_fd_sc_hd__nand3_1 _40213_ (.A(_18223_),
    .B(_18224_),
    .C(_18227_),
    .Y(_18228_));
 sky130_fd_sc_hd__inv_1 _40214_ (.A(_18228_),
    .Y(_18229_));
 sky130_fd_sc_hd__nand2_1 _40215_ (.A(_18222_),
    .B(_18227_),
    .Y(_18230_));
 sky130_fd_sc_hd__inv_1 _40216_ (.A(_18230_),
    .Y(_18231_));
 sky130_fd_sc_hd__nand2_1 _40217_ (.A(_18231_),
    .B(\inst$top.soc.spiflash.phy.deframer.cycle[1] ),
    .Y(_18232_));
 sky130_fd_sc_hd__nor2_1 _40218_ (.A(\inst$top.soc.spiflash.phy.io_streamer.skid_at ),
    .B(\inst$top.soc.spiflash.phy.io_streamer.i_en_0 ),
    .Y(_18233_));
 sky130_fd_sc_hd__inv_1 _40219_ (.A(_18233_),
    .Y(_18234_));
 sky130_fd_sc_hd__nand2_1 _40220_ (.A(_18234_),
    .B(\inst$top.soc.spiflash.phy.deframer.cycle[0] ),
    .Y(_18235_));
 sky130_fd_sc_hd__a21oi_1 _40221_ (.A1(_18223_),
    .A2(_18214_),
    .B1(_18235_),
    .Y(_18236_));
 sky130_fd_sc_hd__o21a_1 _40222_ (.A1(\inst$top.soc.spiflash.phy.deframer.cycle[1] ),
    .A2(_18231_),
    .B1(_18236_),
    .X(_18237_));
 sky130_fd_sc_hd__o211ai_2 _40223_ (.A1(_18214_),
    .A2(_18229_),
    .B1(_18232_),
    .C1(_18237_),
    .Y(_18238_));
 sky130_fd_sc_hd__inv_2 _40224_ (.A(_18238_),
    .Y(_18239_));
 sky130_fd_sc_hd__inv_2 _40225_ (.A(_18205_),
    .Y(_18240_));
 sky130_fd_sc_hd__inv_1 _40226_ (.A(\inst$top.soc.spiflash.ctrl.fsm_state[3] ),
    .Y(_18241_));
 sky130_fd_sc_hd__nor3_1 _40227_ (.A(_18241_),
    .B(\inst$top.soc.spiflash.ctrl.fsm_state[2] ),
    .C(_18193_),
    .Y(_18242_));
 sky130_fd_sc_hd__inv_1 _40228_ (.A(_18242_),
    .Y(_18243_));
 sky130_fd_sc_hd__nand3_1 _40229_ (.A(_18239_),
    .B(_18240_),
    .C(_18243_),
    .Y(_18244_));
 sky130_fd_sc_hd__nand2_1 _40230_ (.A(_18244_),
    .B(_18215_),
    .Y(_18245_));
 sky130_fd_sc_hd__inv_2 _40231_ (.A(_18245_),
    .Y(_18246_));
 sky130_fd_sc_hd__nand2_1 _40232_ (.A(\inst$top.soc.spiflash.ctrl.o_data_count[2] ),
    .B(_02729_),
    .Y(_18247_));
 sky130_fd_sc_hd__inv_1 _40233_ (.A(_18247_),
    .Y(_18248_));
 sky130_fd_sc_hd__nand4_1 _40234_ (.A(net1082),
    .B(_09256_),
    .C(_09346_),
    .D(_18196_),
    .Y(_18249_));
 sky130_fd_sc_hd__o211ai_1 _40235_ (.A1(_18199_),
    .A2(_18248_),
    .B1(_18200_),
    .C1(_18249_),
    .Y(_18250_));
 sky130_fd_sc_hd__nand3_1 _40236_ (.A(_18250_),
    .B(_18241_),
    .C(_18143_),
    .Y(_18251_));
 sky130_fd_sc_hd__nor2_1 _40237_ (.A(_18143_),
    .B(_18199_),
    .Y(_18252_));
 sky130_fd_sc_hd__inv_1 _40238_ (.A(_18252_),
    .Y(_18253_));
 sky130_fd_sc_hd__nand2_1 _40239_ (.A(_18251_),
    .B(_18253_),
    .Y(_18254_));
 sky130_fd_sc_hd__nand2_1 _40240_ (.A(_18246_),
    .B(_18254_),
    .Y(_18255_));
 sky130_fd_sc_hd__inv_1 _40241_ (.A(_18255_),
    .Y(_18256_));
 sky130_fd_sc_hd__nor2_1 _40242_ (.A(\inst$top.soc.spiflash.phy.io_clocker.fsm_state ),
    .B(_18211_),
    .Y(_18257_));
 sky130_fd_sc_hd__inv_1 _40243_ (.A(_18257_),
    .Y(_18258_));
 sky130_fd_sc_hd__nor2_1 _40244_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[7] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[6] ),
    .Y(_18259_));
 sky130_fd_sc_hd__nor2_1 _40245_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[5] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[4] ),
    .Y(_18260_));
 sky130_fd_sc_hd__nand2_1 _40246_ (.A(_18259_),
    .B(_18260_),
    .Y(_18261_));
 sky130_fd_sc_hd__nor2_1 _40247_ (.A(_02741_),
    .B(_02743_),
    .Y(_18262_));
 sky130_fd_sc_hd__nor2_1 _40248_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[13] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[12] ),
    .Y(_18263_));
 sky130_fd_sc_hd__inv_1 _40249_ (.A(_18263_),
    .Y(_18264_));
 sky130_fd_sc_hd__nor2_1 _40250_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[14] ),
    .B(_18264_),
    .Y(_18265_));
 sky130_fd_sc_hd__nor2_1 _40251_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[11] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[10] ),
    .Y(_18266_));
 sky130_fd_sc_hd__nor2_1 _40252_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[9] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[8] ),
    .Y(_18267_));
 sky130_fd_sc_hd__nand2_1 _40253_ (.A(_18266_),
    .B(_18267_),
    .Y(_18268_));
 sky130_fd_sc_hd__inv_1 _40254_ (.A(_18268_),
    .Y(_18269_));
 sky130_fd_sc_hd__inv_1 _40255_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[15] ),
    .Y(_18270_));
 sky130_fd_sc_hd__nor2_1 _40256_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[3] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[2] ),
    .Y(_18271_));
 sky130_fd_sc_hd__nand4_1 _40257_ (.A(_18265_),
    .B(_18269_),
    .C(_18270_),
    .D(_18271_),
    .Y(_18272_));
 sky130_fd_sc_hd__nor3_1 _40258_ (.A(_18261_),
    .B(_18262_),
    .C(_18272_),
    .Y(_18273_));
 sky130_fd_sc_hd__nand3_1 _40259_ (.A(_18256_),
    .B(_18258_),
    .C(_18273_),
    .Y(_18274_));
 sky130_fd_sc_hd__nor2_1 _40260_ (.A(_18213_),
    .B(_18274_),
    .Y(_18275_));
 sky130_fd_sc_hd__inv_1 _40261_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[1] ),
    .Y(_18276_));
 sky130_fd_sc_hd__nor2_1 _40262_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[0] ),
    .B(_18276_),
    .Y(_18277_));
 sky130_fd_sc_hd__nor2_1 _40263_ (.A(_18277_),
    .B(_18240_),
    .Y(_18278_));
 sky130_fd_sc_hd__inv_1 _40264_ (.A(_18278_),
    .Y(_18279_));
 sky130_fd_sc_hd__inv_1 _40265_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[0] ),
    .Y(_18280_));
 sky130_fd_sc_hd__nor3_1 _40266_ (.A(_18276_),
    .B(_18280_),
    .C(_18202_),
    .Y(_18281_));
 sky130_fd_sc_hd__o21ai_0 _40267_ (.A1(_18276_),
    .A2(_18240_),
    .B1(_18209_),
    .Y(_18282_));
 sky130_fd_sc_hd__nor2_1 _40268_ (.A(_18281_),
    .B(_18282_),
    .Y(_18283_));
 sky130_fd_sc_hd__inv_1 _40269_ (.A(_18281_),
    .Y(_18284_));
 sky130_fd_sc_hd__o21ai_1 _40270_ (.A1(_18279_),
    .A2(_18283_),
    .B1(_18284_),
    .Y(_18285_));
 sky130_fd_sc_hd__inv_1 _40271_ (.A(_18277_),
    .Y(_18286_));
 sky130_fd_sc_hd__nor2_1 _40272_ (.A(_18286_),
    .B(_18202_),
    .Y(_18287_));
 sky130_fd_sc_hd__nor2_1 _40273_ (.A(_18208_),
    .B(_18287_),
    .Y(_18288_));
 sky130_fd_sc_hd__nand2_1 _40274_ (.A(_18288_),
    .B(_18279_),
    .Y(_18289_));
 sky130_fd_sc_hd__nor2_1 _40275_ (.A(_18289_),
    .B(_18283_),
    .Y(_18290_));
 sky130_fd_sc_hd__inv_1 _40276_ (.A(_18210_),
    .Y(_18291_));
 sky130_fd_sc_hd__a21oi_1 _40277_ (.A1(_18290_),
    .A2(_18291_),
    .B1(_18287_),
    .Y(_18292_));
 sky130_fd_sc_hd__inv_1 _40278_ (.A(_18285_),
    .Y(_18293_));
 sky130_fd_sc_hd__nand3_1 _40279_ (.A(_18292_),
    .B(_18204_),
    .C(_18293_),
    .Y(_18294_));
 sky130_fd_sc_hd__nand2_1 _40280_ (.A(_18292_),
    .B(_18293_),
    .Y(_18295_));
 sky130_fd_sc_hd__nand2_1 _40281_ (.A(_18295_),
    .B(\inst$top.soc.spiflash.phy.enframer.cycle[2] ),
    .Y(_18296_));
 sky130_fd_sc_hd__a21oi_1 _40282_ (.A1(_18285_),
    .A2(net2578),
    .B1(_02744_),
    .Y(_18297_));
 sky130_fd_sc_hd__o2111ai_1 _40283_ (.A1(net2578),
    .A2(_18285_),
    .B1(_18294_),
    .C1(_18296_),
    .D1(_18297_),
    .Y(_18298_));
 sky130_fd_sc_hd__nand2_1 _40284_ (.A(_18298_),
    .B(_18212_),
    .Y(_18299_));
 sky130_fd_sc_hd__nand2_1 _40285_ (.A(_18275_),
    .B(_18299_),
    .Y(_18300_));
 sky130_fd_sc_hd__o21ai_0 _40286_ (.A1(_18196_),
    .A2(_18203_),
    .B1(_18300_),
    .Y(_18301_));
 sky130_fd_sc_hd__nand2_1 _40287_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.RawControl.port__w_data ),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb$16 ),
    .Y(_18302_));
 sky130_fd_sc_hd__inv_1 _40288_ (.A(_18144_),
    .Y(_18303_));
 sky130_fd_sc_hd__nor2_1 _40289_ (.A(_18150_),
    .B(_18303_),
    .Y(_18304_));
 sky130_fd_sc_hd__inv_1 _40290_ (.A(_18304_),
    .Y(_18305_));
 sky130_fd_sc_hd__nor2_1 _40291_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12.w_stb ),
    .B(_18305_),
    .Y(_18306_));
 sky130_fd_sc_hd__nor2_1 _40292_ (.A(_18243_),
    .B(_18239_),
    .Y(_18307_));
 sky130_fd_sc_hd__nand3_1 _40293_ (.A(net1082),
    .B(_09256_),
    .C(_09346_),
    .Y(_18308_));
 sky130_fd_sc_hd__nand2_1 _40294_ (.A(_18308_),
    .B(_18194_),
    .Y(_18309_));
 sky130_fd_sc_hd__a21oi_1 _40295_ (.A1(_18192_),
    .A2(_18197_),
    .B1(_18241_),
    .Y(_18310_));
 sky130_fd_sc_hd__nor2_1 _40296_ (.A(\inst$top.soc.spiflash.ctrl.fsm_state[0] ),
    .B(_18200_),
    .Y(_18311_));
 sky130_fd_sc_hd__nand2_1 _40297_ (.A(_18311_),
    .B(_18139_),
    .Y(_18312_));
 sky130_fd_sc_hd__nor2_1 _40298_ (.A(_02725_),
    .B(_18312_),
    .Y(_18313_));
 sky130_fd_sc_hd__inv_1 _40299_ (.A(\inst$top.soc.spiflash.ctrl.o_dummy_count[0] ),
    .Y(_18314_));
 sky130_fd_sc_hd__inv_1 _40300_ (.A(\inst$top.soc.spiflash.ctrl.o_dummy_count[1] ),
    .Y(_18315_));
 sky130_fd_sc_hd__nor2_1 _40301_ (.A(_18207_),
    .B(_18140_),
    .Y(_18316_));
 sky130_fd_sc_hd__inv_1 _40302_ (.A(_18316_),
    .Y(_18317_));
 sky130_fd_sc_hd__a21oi_1 _40303_ (.A1(_18314_),
    .A2(_18315_),
    .B1(_18317_),
    .Y(_18318_));
 sky130_fd_sc_hd__nor3_1 _40304_ (.A(_18310_),
    .B(_18313_),
    .C(_18318_),
    .Y(_18319_));
 sky130_fd_sc_hd__o21ai_0 _40305_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.raw_enable._storage ),
    .A2(_18309_),
    .B1(_18319_),
    .Y(_18320_));
 sky130_fd_sc_hd__inv_1 _40306_ (.A(\inst$top.soc.spiflash.ctrl.i_data_count[2] ),
    .Y(_18321_));
 sky130_fd_sc_hd__a31oi_1 _40307_ (.A1(_18239_),
    .A2(_02738_),
    .A3(_18321_),
    .B1(_18240_),
    .Y(_18322_));
 sky130_fd_sc_hd__a2111oi_0 _40308_ (.A1(_18302_),
    .A2(_18306_),
    .B1(_18307_),
    .C1(_18320_),
    .D1(_18322_),
    .Y(_18323_));
 sky130_fd_sc_hd__nand2_1 _40309_ (.A(_18301_),
    .B(_18323_),
    .Y(_18324_));
 sky130_fd_sc_hd__nand2_1 _40310_ (.A(_18198_),
    .B(_18311_),
    .Y(_18325_));
 sky130_fd_sc_hd__o21ai_0 _40311_ (.A1(_18150_),
    .A2(_18302_),
    .B1(_18144_),
    .Y(_18326_));
 sky130_fd_sc_hd__inv_1 _40312_ (.A(_18312_),
    .Y(_18327_));
 sky130_fd_sc_hd__o21ai_0 _40314_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[0] ),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[1] ),
    .B1(_18327_),
    .Y(_18329_));
 sky130_fd_sc_hd__nor2_1 _40315_ (.A(\inst$top.soc.spiflash.ctrl.fsm_state[3] ),
    .B(_18192_),
    .Y(_18330_));
 sky130_fd_sc_hd__or2_2 _40316_ (.A(_18194_),
    .B(_18310_),
    .X(_18331_));
 sky130_fd_sc_hd__nand2_1 _40317_ (.A(_18331_),
    .B(_18150_),
    .Y(_18332_));
 sky130_fd_sc_hd__inv_1 _40318_ (.A(_18332_),
    .Y(_18333_));
 sky130_fd_sc_hd__a41oi_1 _40319_ (.A1(_18325_),
    .A2(_18326_),
    .A3(_18329_),
    .A4(_18330_),
    .B1(_18333_),
    .Y(_18334_));
 sky130_fd_sc_hd__o21ai_0 _40320_ (.A1(_18334_),
    .A2(_18324_),
    .B1(net2059),
    .Y(_18335_));
 sky130_fd_sc_hd__a21oi_2 _40321_ (.A1(_18141_),
    .A2(_18324_),
    .B1(_18335_),
    .Y(_05179_));
 sky130_fd_sc_hd__nand3_1 _40322_ (.A(_18332_),
    .B(_18305_),
    .C(_18329_),
    .Y(_18336_));
 sky130_fd_sc_hd__o21ai_0 _40323_ (.A1(_18336_),
    .A2(_18324_),
    .B1(net2059),
    .Y(_18337_));
 sky130_fd_sc_hd__a21oi_2 _40324_ (.A1(_18200_),
    .A2(_18324_),
    .B1(_18337_),
    .Y(_05180_));
 sky130_fd_sc_hd__nor3_1 _40325_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[0] ),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[1] ),
    .C(_18312_),
    .Y(_18338_));
 sky130_fd_sc_hd__nor3_1 _40326_ (.A(_18205_),
    .B(_18316_),
    .C(_18338_),
    .Y(_18339_));
 sky130_fd_sc_hd__nand2_1 _40327_ (.A(_18339_),
    .B(_18303_),
    .Y(_18340_));
 sky130_fd_sc_hd__o21ai_0 _40328_ (.A1(_18340_),
    .A2(_18324_),
    .B1(net2059),
    .Y(_18341_));
 sky130_fd_sc_hd__a21oi_2 _40329_ (.A1(_18197_),
    .A2(_18324_),
    .B1(_18341_),
    .Y(_05181_));
 sky130_fd_sc_hd__nor2_1 _40330_ (.A(_18208_),
    .B(_18324_),
    .Y(_18342_));
 sky130_fd_sc_hd__a211oi_2 _40331_ (.A1(_18324_),
    .A2(_18241_),
    .B1(net2947),
    .C1(_18342_),
    .Y(_05182_));
 sky130_fd_sc_hd__nor2_1 _40332_ (.A(_18240_),
    .B(_18238_),
    .Y(_18343_));
 sky130_fd_sc_hd__inv_1 _40333_ (.A(_18343_),
    .Y(_18344_));
 sky130_fd_sc_hd__nand2_1 _40334_ (.A(_18344_),
    .B(\inst$top.soc.spiflash.ctrl.i_data_count[0] ),
    .Y(_18345_));
 sky130_fd_sc_hd__nand2_1 _40335_ (.A(_18343_),
    .B(_02732_),
    .Y(_18346_));
 sky130_fd_sc_hd__nand4_1 _40336_ (.A(_18239_),
    .B(_02738_),
    .C(_18321_),
    .D(_18205_),
    .Y(_18347_));
 sky130_fd_sc_hd__nand2_1 _40337_ (.A(_18347_),
    .B(net2052),
    .Y(_18348_));
 sky130_fd_sc_hd__a21oi_1 _40338_ (.A1(_18345_),
    .A2(_18346_),
    .B1(_18348_),
    .Y(_05183_));
 sky130_fd_sc_hd__o21ai_0 _40339_ (.A1(_02735_),
    .A2(_18344_),
    .B1(net2048),
    .Y(_18349_));
 sky130_fd_sc_hd__a21oi_1 _40340_ (.A1(_02733_),
    .A2(_18344_),
    .B1(_18349_),
    .Y(_05184_));
 sky130_fd_sc_hd__nand2_1 _40341_ (.A(_18343_),
    .B(_02738_),
    .Y(_18350_));
 sky130_fd_sc_hd__nand3_1 _40342_ (.A(_18350_),
    .B(net2053),
    .C(\inst$top.soc.spiflash.ctrl.i_data_count[2] ),
    .Y(_18351_));
 sky130_fd_sc_hd__inv_2 _40343_ (.A(_18351_),
    .Y(_05185_));
 sky130_fd_sc_hd__inv_1 _40344_ (.A(_02741_),
    .Y(_18352_));
 sky130_fd_sc_hd__inv_1 _40345_ (.A(_18271_),
    .Y(_18353_));
 sky130_fd_sc_hd__nor2_1 _40346_ (.A(_18352_),
    .B(_18353_),
    .Y(_18354_));
 sky130_fd_sc_hd__inv_1 _40347_ (.A(_18354_),
    .Y(_18355_));
 sky130_fd_sc_hd__nand2_1 _40348_ (.A(_18271_),
    .B(_02743_),
    .Y(_18356_));
 sky130_fd_sc_hd__nor2_1 _40349_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[15] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[14] ),
    .Y(_18357_));
 sky130_fd_sc_hd__nand3_1 _40350_ (.A(_18269_),
    .B(_18263_),
    .C(_18357_),
    .Y(_18358_));
 sky130_fd_sc_hd__a211oi_1 _40351_ (.A1(_18355_),
    .A2(_18356_),
    .B1(_18261_),
    .C1(_18358_),
    .Y(_18359_));
 sky130_fd_sc_hd__o211a_1 _40352_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.fsm_state ),
    .A2(_18211_),
    .B1(_18359_),
    .C1(_18246_),
    .X(_18360_));
 sky130_fd_sc_hd__inv_1 _40353_ (.A(_18213_),
    .Y(_18361_));
 sky130_fd_sc_hd__nand4_1 _40354_ (.A(_18360_),
    .B(_18299_),
    .C(_18361_),
    .D(_18254_),
    .Y(_18362_));
 sky130_fd_sc_hd__o21ai_0 _40355_ (.A1(_18327_),
    .A2(_18194_),
    .B1(_18309_),
    .Y(_18363_));
 sky130_fd_sc_hd__a21oi_1 _40356_ (.A1(_18362_),
    .A2(_18194_),
    .B1(_18363_),
    .Y(_18364_));
 sky130_fd_sc_hd__o21ai_0 _40357_ (.A1(_02725_),
    .A2(_18300_),
    .B1(net1638),
    .Y(_18365_));
 sky130_fd_sc_hd__and2_1 _40358_ (.A(_18364_),
    .B(_18365_),
    .X(_18366_));
 sky130_fd_sc_hd__nor2_1 _40359_ (.A(\inst$top.soc.spiflash.ctrl.o_addr_count[0] ),
    .B(_18366_),
    .Y(_18367_));
 sky130_fd_sc_hd__nand2_1 _40360_ (.A(net1638),
    .B(_02723_),
    .Y(_18368_));
 sky130_fd_sc_hd__nand2_1 _40361_ (.A(_18366_),
    .B(_18368_),
    .Y(_18369_));
 sky130_fd_sc_hd__nand2_1 _40362_ (.A(_18369_),
    .B(net2027),
    .Y(_18370_));
 sky130_fd_sc_hd__nor2_2 _40363_ (.A(_18367_),
    .B(_18370_),
    .Y(_05186_));
 sky130_fd_sc_hd__nor2_1 _40364_ (.A(\inst$top.soc.spiflash.ctrl.o_addr_count[1] ),
    .B(_18366_),
    .Y(_18371_));
 sky130_fd_sc_hd__nand4_1 _40365_ (.A(_18364_),
    .B(_18365_),
    .C(_02726_),
    .D(net1638),
    .Y(_18372_));
 sky130_fd_sc_hd__nand2_1 _40366_ (.A(_18372_),
    .B(net2049),
    .Y(_18373_));
 sky130_fd_sc_hd__nor2_2 _40367_ (.A(_18371_),
    .B(_18373_),
    .Y(_05187_));
 sky130_fd_sc_hd__nor3_1 _40368_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[14] ),
    .B(_18264_),
    .C(_18261_),
    .Y(_18374_));
 sky130_fd_sc_hd__nand3_1 _40369_ (.A(_18374_),
    .B(_18270_),
    .C(_18269_),
    .Y(_18375_));
 sky130_fd_sc_hd__a21oi_1 _40370_ (.A1(_18356_),
    .A2(_18355_),
    .B1(_18375_),
    .Y(_18376_));
 sky130_fd_sc_hd__nand2_1 _40371_ (.A(_18256_),
    .B(_18376_),
    .Y(_18377_));
 sky130_fd_sc_hd__nor3b_1 _40372_ (.A(_18257_),
    .B(_18377_),
    .C_N(_18299_),
    .Y(_18378_));
 sky130_fd_sc_hd__nand4_1 _40373_ (.A(_18378_),
    .B(_18205_),
    .C(_18361_),
    .D(_18247_),
    .Y(_18379_));
 sky130_fd_sc_hd__xor2_1 _40374_ (.A(\inst$top.soc.spiflash.ctrl.o_data_count[0] ),
    .B(_18379_),
    .X(_18380_));
 sky130_fd_sc_hd__nor2_2 _40375_ (.A(_18348_),
    .B(_18380_),
    .Y(_05188_));
 sky130_fd_sc_hd__inv_1 _40376_ (.A(_18300_),
    .Y(_18381_));
 sky130_fd_sc_hd__nand3b_1 _40377_ (.A_N(_02730_),
    .B(_18381_),
    .C(_18247_),
    .Y(_18382_));
 sky130_fd_sc_hd__o21ai_0 _40378_ (.A1(_18248_),
    .A2(_18300_),
    .B1(_02728_),
    .Y(_18383_));
 sky130_fd_sc_hd__nand3_1 _40379_ (.A(_18382_),
    .B(_18383_),
    .C(_18322_),
    .Y(_18384_));
 sky130_fd_sc_hd__nand2_1 _40380_ (.A(_18240_),
    .B(\inst$top.soc.spiflash.ctrl.o_data_count[1] ),
    .Y(_18385_));
 sky130_fd_sc_hd__a21oi_1 _40381_ (.A1(_18384_),
    .A2(_18385_),
    .B1(net2947),
    .Y(_05189_));
 sky130_fd_sc_hd__nand3_1 _40382_ (.A(_18378_),
    .B(_02731_),
    .C(_18361_),
    .Y(_18386_));
 sky130_fd_sc_hd__inv_1 _40383_ (.A(\inst$top.soc.spiflash.ctrl.o_data_count[2] ),
    .Y(_18387_));
 sky130_fd_sc_hd__nand2_1 _40384_ (.A(_18386_),
    .B(_18387_),
    .Y(_18388_));
 sky130_fd_sc_hd__nor2_1 _40385_ (.A(_02729_),
    .B(_18387_),
    .Y(_18389_));
 sky130_fd_sc_hd__nand4_1 _40386_ (.A(_18378_),
    .B(_02731_),
    .C(_18361_),
    .D(_18389_),
    .Y(_18390_));
 sky130_fd_sc_hd__nand3_1 _40387_ (.A(_18388_),
    .B(_18390_),
    .C(_18322_),
    .Y(_18391_));
 sky130_fd_sc_hd__nand2_1 _40388_ (.A(_18240_),
    .B(\inst$top.soc.spiflash.ctrl.o_data_count[2] ),
    .Y(_18392_));
 sky130_fd_sc_hd__a21oi_2 _40389_ (.A1(_18391_),
    .A2(_18392_),
    .B1(net2947),
    .Y(_05190_));
 sky130_fd_sc_hd__nor3_1 _40390_ (.A(\inst$top.soc.spiflash.ctrl.o_dummy_count[0] ),
    .B(\inst$top.soc.spiflash.ctrl.o_dummy_count[1] ),
    .C(_18317_),
    .Y(_18393_));
 sky130_fd_sc_hd__nor4_1 _40391_ (.A(_18202_),
    .B(_18313_),
    .C(_18338_),
    .D(_18393_),
    .Y(_18394_));
 sky130_fd_sc_hd__nand2_1 _40392_ (.A(_18381_),
    .B(_18394_),
    .Y(_18395_));
 sky130_fd_sc_hd__nand2_1 _40393_ (.A(_18316_),
    .B(_18314_),
    .Y(_18396_));
 sky130_fd_sc_hd__o21ai_0 _40394_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[0] ),
    .A2(_18316_),
    .B1(_18396_),
    .Y(_18397_));
 sky130_fd_sc_hd__o21ai_0 _40395_ (.A1(_18397_),
    .A2(_18395_),
    .B1(net2059),
    .Y(_18398_));
 sky130_fd_sc_hd__a21oi_2 _40396_ (.A1(_18314_),
    .A2(_18395_),
    .B1(_18398_),
    .Y(_05191_));
 sky130_fd_sc_hd__nand2_1 _40397_ (.A(_18317_),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[1] ),
    .Y(_18399_));
 sky130_fd_sc_hd__o21ai_0 _40398_ (.A1(_18315_),
    .A2(_18317_),
    .B1(_18399_),
    .Y(_18400_));
 sky130_fd_sc_hd__xor2_1 _40399_ (.A(_18397_),
    .B(_18400_),
    .X(_18401_));
 sky130_fd_sc_hd__o21ai_0 _40400_ (.A1(_18401_),
    .A2(_18395_),
    .B1(net2059),
    .Y(_18402_));
 sky130_fd_sc_hd__a21oi_2 _40401_ (.A1(_18315_),
    .A2(_18395_),
    .B1(_18402_),
    .Y(_05192_));
 sky130_fd_sc_hd__nor2_1 _40402_ (.A(_18243_),
    .B(_18238_),
    .Y(_18403_));
 sky130_fd_sc_hd__inv_1 _40404_ (.A(\inst$top.soc.spiflash.phy.io_streamer.buffer_io1.i_ff ),
    .Y(_18405_));
 sky130_fd_sc_hd__nand2_1 _40405_ (.A(\inst$top.soc.spiflash.phy.io_streamer.skid_at ),
    .B(\inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io1 ),
    .Y(_18406_));
 sky130_fd_sc_hd__o21ai_0 _40406_ (.A1(\inst$top.soc.spiflash.phy.io_streamer.skid_at ),
    .A2(_18405_),
    .B1(_18406_),
    .Y(_18407_));
 sky130_fd_sc_hd__inv_1 _40407_ (.A(_18407_),
    .Y(_18408_));
 sky130_fd_sc_hd__inv_1 _40408_ (.A(\inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io0 ),
    .Y(_18409_));
 sky130_fd_sc_hd__nand2_1 _40409_ (.A(_18409_),
    .B(\inst$top.soc.spiflash.phy.io_streamer.skid_at ),
    .Y(_18410_));
 sky130_fd_sc_hd__o211ai_1 _40410_ (.A1(\inst$top.soc.spiflash.phy.io_streamer.skid_at ),
    .A2(\inst$top.soc.spiflash.phy.io_streamer.buffer_io0.i_ff ),
    .B1(_18410_),
    .C1(_18222_),
    .Y(_18411_));
 sky130_fd_sc_hd__o21a_1 _40411_ (.A1(_18408_),
    .A2(_18228_),
    .B1(_18411_),
    .X(_18412_));
 sky130_fd_sc_hd__o21ai_0 _40414_ (.A1(\inst$top.soc.spiflash.ctrl.r_data[0] ),
    .A2(_18403_),
    .B1(net2125),
    .Y(_18415_));
 sky130_fd_sc_hd__a21oi_1 _40415_ (.A1(net882),
    .A2(_18412_),
    .B1(_18415_),
    .Y(_05193_));
 sky130_fd_sc_hd__a22oi_1 _40416_ (.A1(_18222_),
    .A2(_18407_),
    .B1(_18229_),
    .B2(\inst$top.soc.spiflash.phy.deframer.data_reg[0] ),
    .Y(_18416_));
 sky130_fd_sc_hd__o21ai_0 _40417_ (.A1(\inst$top.soc.spiflash.ctrl.r_data[1] ),
    .A2(net882),
    .B1(net2057),
    .Y(_18417_));
 sky130_fd_sc_hd__a21oi_1 _40418_ (.A1(net882),
    .A2(_18416_),
    .B1(_18417_),
    .Y(_05194_));
 sky130_fd_sc_hd__nand2_1 _40419_ (.A(_18229_),
    .B(\inst$top.soc.spiflash.phy.deframer.data_reg[1] ),
    .Y(_18418_));
 sky130_fd_sc_hd__nor2_1 _40420_ (.A(_18227_),
    .B(_18223_),
    .Y(_18419_));
 sky130_fd_sc_hd__nand2_1 _40421_ (.A(_18419_),
    .B(\inst$top.soc.spiflash.phy.deframer.data_reg[0] ),
    .Y(_18420_));
 sky130_fd_sc_hd__inv_1 _40422_ (.A(\inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io2 ),
    .Y(_18421_));
 sky130_fd_sc_hd__nand2_1 _40423_ (.A(_18215_),
    .B(\inst$top.soc.spiflash.phy.io_streamer.buffer_io2.i_ff ),
    .Y(_18422_));
 sky130_fd_sc_hd__o21ai_0 _40424_ (.A1(_18215_),
    .A2(_18421_),
    .B1(_18422_),
    .Y(_18423_));
 sky130_fd_sc_hd__nand2_1 _40425_ (.A(_18231_),
    .B(_18423_),
    .Y(_18424_));
 sky130_fd_sc_hd__nand3_1 _40426_ (.A(_18418_),
    .B(_18420_),
    .C(_18424_),
    .Y(_18425_));
 sky130_fd_sc_hd__inv_1 _40427_ (.A(_18403_),
    .Y(_18426_));
 sky130_fd_sc_hd__nor2_1 _40428_ (.A(_18425_),
    .B(_18426_),
    .Y(_18427_));
 sky130_fd_sc_hd__o21ai_0 _40429_ (.A1(\inst$top.soc.spiflash.ctrl.r_data[2] ),
    .A2(net882),
    .B1(net2057),
    .Y(_18428_));
 sky130_fd_sc_hd__nor2_1 _40430_ (.A(_18427_),
    .B(_18428_),
    .Y(_05195_));
 sky130_fd_sc_hd__inv_1 _40431_ (.A(\inst$top.soc.spiflash.phy.deframer.data_reg[2] ),
    .Y(_18429_));
 sky130_fd_sc_hd__nand2_1 _40432_ (.A(_18419_),
    .B(\inst$top.soc.spiflash.phy.deframer.data_reg[1] ),
    .Y(_18430_));
 sky130_fd_sc_hd__inv_1 _40433_ (.A(\inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io3 ),
    .Y(_18431_));
 sky130_fd_sc_hd__nand2_1 _40434_ (.A(_18215_),
    .B(\inst$top.soc.spiflash.phy.io_streamer.buffer_io3.i_ff ),
    .Y(_18432_));
 sky130_fd_sc_hd__o21ai_0 _40435_ (.A1(_18215_),
    .A2(_18431_),
    .B1(_18432_),
    .Y(_18433_));
 sky130_fd_sc_hd__nand2_1 _40436_ (.A(_18231_),
    .B(_18433_),
    .Y(_18434_));
 sky130_fd_sc_hd__o211ai_1 _40437_ (.A1(_18429_),
    .A2(_18228_),
    .B1(_18430_),
    .C1(_18434_),
    .Y(_18435_));
 sky130_fd_sc_hd__nor2_1 _40438_ (.A(_18435_),
    .B(_18426_),
    .Y(_18436_));
 sky130_fd_sc_hd__o21ai_0 _40439_ (.A1(\inst$top.soc.spiflash.ctrl.r_data[3] ),
    .A2(net882),
    .B1(net2119),
    .Y(_18437_));
 sky130_fd_sc_hd__nor2_1 _40440_ (.A(_18436_),
    .B(_18437_),
    .Y(_05196_));
 sky130_fd_sc_hd__inv_1 _40441_ (.A(\inst$top.soc.spiflash.phy.deframer.data_reg[3] ),
    .Y(_18438_));
 sky130_fd_sc_hd__nand2_1 _40442_ (.A(_18419_),
    .B(\inst$top.soc.spiflash.phy.deframer.data_reg[2] ),
    .Y(_18439_));
 sky130_fd_sc_hd__nand2_1 _40443_ (.A(_18231_),
    .B(\inst$top.soc.spiflash.phy.deframer.data_reg[0] ),
    .Y(_18440_));
 sky130_fd_sc_hd__o211ai_1 _40444_ (.A1(_18438_),
    .A2(_18228_),
    .B1(_18439_),
    .C1(_18440_),
    .Y(_18441_));
 sky130_fd_sc_hd__nor2_1 _40445_ (.A(_18441_),
    .B(_18426_),
    .Y(_18442_));
 sky130_fd_sc_hd__o21ai_0 _40446_ (.A1(\inst$top.soc.spiflash.ctrl.r_data[4] ),
    .A2(net882),
    .B1(net2119),
    .Y(_18443_));
 sky130_fd_sc_hd__nor2_1 _40447_ (.A(_18442_),
    .B(_18443_),
    .Y(_05197_));
 sky130_fd_sc_hd__nand2_1 _40448_ (.A(_18426_),
    .B(\inst$top.soc.spiflash.ctrl.r_data[5] ),
    .Y(_18444_));
 sky130_fd_sc_hd__nand2_1 _40449_ (.A(_18229_),
    .B(\inst$top.soc.spiflash.phy.deframer.data_reg[4] ),
    .Y(_18445_));
 sky130_fd_sc_hd__nand2_1 _40450_ (.A(_18419_),
    .B(\inst$top.soc.spiflash.phy.deframer.data_reg[3] ),
    .Y(_18446_));
 sky130_fd_sc_hd__nand2_1 _40451_ (.A(_18231_),
    .B(\inst$top.soc.spiflash.phy.deframer.data_reg[1] ),
    .Y(_18447_));
 sky130_fd_sc_hd__nand3_1 _40452_ (.A(_18445_),
    .B(_18446_),
    .C(_18447_),
    .Y(_18448_));
 sky130_fd_sc_hd__nand2_1 _40453_ (.A(net882),
    .B(_18448_),
    .Y(_18449_));
 sky130_fd_sc_hd__a21oi_1 _40454_ (.A1(_18444_),
    .A2(_18449_),
    .B1(net2979),
    .Y(_05198_));
 sky130_fd_sc_hd__nand2_1 _40455_ (.A(_18419_),
    .B(\inst$top.soc.spiflash.phy.deframer.data_reg[4] ),
    .Y(_18450_));
 sky130_fd_sc_hd__nand2_1 _40456_ (.A(_18229_),
    .B(\inst$top.soc.spiflash.phy.deframer.data_reg[5] ),
    .Y(_18451_));
 sky130_fd_sc_hd__o211ai_1 _40457_ (.A1(_18429_),
    .A2(_18230_),
    .B1(_18450_),
    .C1(_18451_),
    .Y(_18452_));
 sky130_fd_sc_hd__nor2_1 _40458_ (.A(_18452_),
    .B(_18426_),
    .Y(_18453_));
 sky130_fd_sc_hd__o21ai_0 _40459_ (.A1(\inst$top.soc.spiflash.ctrl.r_data[6] ),
    .A2(net882),
    .B1(net2119),
    .Y(_18454_));
 sky130_fd_sc_hd__nor2_1 _40460_ (.A(_18453_),
    .B(_18454_),
    .Y(_05199_));
 sky130_fd_sc_hd__nand2_1 _40461_ (.A(_18419_),
    .B(\inst$top.soc.spiflash.phy.deframer.data_reg[5] ),
    .Y(_18455_));
 sky130_fd_sc_hd__o21ai_0 _40462_ (.A1(_18438_),
    .A2(_18230_),
    .B1(_18455_),
    .Y(_18456_));
 sky130_fd_sc_hd__a21oi_1 _40463_ (.A1(\inst$top.soc.spiflash.phy.deframer.data_reg[6] ),
    .A2(_18229_),
    .B1(_18456_),
    .Y(_18457_));
 sky130_fd_sc_hd__o21ai_0 _40464_ (.A1(\inst$top.soc.spiflash.ctrl.r_data[7] ),
    .A2(net882),
    .B1(net2119),
    .Y(_18458_));
 sky130_fd_sc_hd__a21oi_1 _40465_ (.A1(net882),
    .A2(_18457_),
    .B1(_18458_),
    .Y(_05200_));
 sky130_fd_sc_hd__inv_1 _40466_ (.A(\inst$top.soc.spiflash.ctrl.raw_tx_data[0] ),
    .Y(_18459_));
 sky130_fd_sc_hd__nand3_1 _40467_ (.A(_18304_),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12.w_stb ),
    .C(_18302_),
    .Y(_18460_));
 sky130_fd_sc_hd__o21ai_0 _40469_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[0] ),
    .A2(net1023),
    .B1(net2061),
    .Y(_18462_));
 sky130_fd_sc_hd__a21oi_1 _40470_ (.A1(_18459_),
    .A2(net1023),
    .B1(_18462_),
    .Y(_05201_));
 sky130_fd_sc_hd__inv_1 _40471_ (.A(\inst$top.soc.spiflash.ctrl.raw_tx_data[1] ),
    .Y(_18463_));
 sky130_fd_sc_hd__o21ai_0 _40472_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[1] ),
    .A2(net1023),
    .B1(net2061),
    .Y(_18464_));
 sky130_fd_sc_hd__a21oi_1 _40473_ (.A1(_18463_),
    .A2(net1023),
    .B1(_18464_),
    .Y(_05202_));
 sky130_fd_sc_hd__inv_1 _40474_ (.A(\inst$top.soc.spiflash.ctrl.raw_tx_data[2] ),
    .Y(_18465_));
 sky130_fd_sc_hd__o21ai_0 _40475_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[2] ),
    .A2(net1022),
    .B1(net2059),
    .Y(_18466_));
 sky130_fd_sc_hd__a21oi_1 _40476_ (.A1(_18465_),
    .A2(net1022),
    .B1(_18466_),
    .Y(_05203_));
 sky130_fd_sc_hd__inv_1 _40477_ (.A(\inst$top.soc.spiflash.ctrl.raw_tx_data[3] ),
    .Y(_18467_));
 sky130_fd_sc_hd__o21ai_0 _40478_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[3] ),
    .A2(net1022),
    .B1(net2061),
    .Y(_18468_));
 sky130_fd_sc_hd__a21oi_1 _40479_ (.A1(_18467_),
    .A2(net1023),
    .B1(_18468_),
    .Y(_05204_));
 sky130_fd_sc_hd__inv_1 _40480_ (.A(\inst$top.soc.spiflash.ctrl.raw_tx_data[4] ),
    .Y(_18469_));
 sky130_fd_sc_hd__o21ai_0 _40481_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[4] ),
    .A2(net1022),
    .B1(net2059),
    .Y(_18470_));
 sky130_fd_sc_hd__a21oi_1 _40482_ (.A1(_18469_),
    .A2(net1022),
    .B1(_18470_),
    .Y(_05205_));
 sky130_fd_sc_hd__inv_1 _40483_ (.A(\inst$top.soc.spiflash.ctrl.raw_tx_data[5] ),
    .Y(_18471_));
 sky130_fd_sc_hd__o21ai_0 _40484_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[5] ),
    .A2(net1022),
    .B1(net2059),
    .Y(_18472_));
 sky130_fd_sc_hd__a21oi_1 _40485_ (.A1(_18471_),
    .A2(net1022),
    .B1(_18472_),
    .Y(_05206_));
 sky130_fd_sc_hd__inv_1 _40486_ (.A(\inst$top.soc.spiflash.ctrl.raw_tx_data[6] ),
    .Y(_18473_));
 sky130_fd_sc_hd__o21ai_0 _40487_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[6] ),
    .A2(net1022),
    .B1(net2061),
    .Y(_18474_));
 sky130_fd_sc_hd__a21oi_1 _40488_ (.A1(_18473_),
    .A2(net1023),
    .B1(_18474_),
    .Y(_05207_));
 sky130_fd_sc_hd__inv_1 _40489_ (.A(\inst$top.soc.spiflash.ctrl.raw_tx_data[7] ),
    .Y(_18475_));
 sky130_fd_sc_hd__o21ai_0 _40492_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[7] ),
    .A2(net1022),
    .B1(net2059),
    .Y(_18478_));
 sky130_fd_sc_hd__a21oi_1 _40493_ (.A1(_18475_),
    .A2(net1022),
    .B1(_18478_),
    .Y(_05208_));
 sky130_fd_sc_hd__nand3_1 _40494_ (.A(_18253_),
    .B(net2052),
    .C(_18325_),
    .Y(_18479_));
 sky130_fd_sc_hd__a21oi_1 _40495_ (.A1(_18347_),
    .A2(_12692_),
    .B1(_18479_),
    .Y(_05209_));
 sky130_fd_sc_hd__nand3_1 _40496_ (.A(_18343_),
    .B(_18321_),
    .C(_02734_),
    .Y(_18480_));
 sky130_fd_sc_hd__inv_1 _40497_ (.A(net866),
    .Y(_18481_));
 sky130_fd_sc_hd__o21ai_0 _40498_ (.A1(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[0] ),
    .A2(_18481_),
    .B1(net2052),
    .Y(_18482_));
 sky130_fd_sc_hd__a21oi_1 _40499_ (.A1(_18412_),
    .A2(_18481_),
    .B1(_18482_),
    .Y(_05210_));
 sky130_fd_sc_hd__nand3_1 _40500_ (.A(_18343_),
    .B(_18321_),
    .C(_02737_),
    .Y(_18483_));
 sky130_fd_sc_hd__o21ai_0 _40502_ (.A1(_18425_),
    .A2(_18483_),
    .B1(net2055),
    .Y(_18485_));
 sky130_fd_sc_hd__a21oi_1 _40503_ (.A1(_12720_),
    .A2(net865),
    .B1(_18485_),
    .Y(_05211_));
 sky130_fd_sc_hd__o21ai_0 _40504_ (.A1(_18435_),
    .A2(net865),
    .B1(net2054),
    .Y(_18486_));
 sky130_fd_sc_hd__a21oi_1 _40505_ (.A1(_12730_),
    .A2(net865),
    .B1(_18486_),
    .Y(_05212_));
 sky130_fd_sc_hd__inv_1 _40506_ (.A(net865),
    .Y(_18487_));
 sky130_fd_sc_hd__nor2_1 _40507_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[12] ),
    .B(_18487_),
    .Y(_18488_));
 sky130_fd_sc_hd__o21ai_0 _40508_ (.A1(_18441_),
    .A2(net865),
    .B1(net2056),
    .Y(_18489_));
 sky130_fd_sc_hd__nor2_1 _40509_ (.A(_18488_),
    .B(_18489_),
    .Y(_05213_));
 sky130_fd_sc_hd__nor2_1 _40510_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[13] ),
    .B(_18487_),
    .Y(_18490_));
 sky130_fd_sc_hd__o21ai_0 _40511_ (.A1(_18448_),
    .A2(net865),
    .B1(net2056),
    .Y(_18491_));
 sky130_fd_sc_hd__nor2_1 _40512_ (.A(_18490_),
    .B(_18491_),
    .Y(_05214_));
 sky130_fd_sc_hd__o21ai_0 _40513_ (.A1(_18452_),
    .A2(net865),
    .B1(net2054),
    .Y(_18492_));
 sky130_fd_sc_hd__a21oi_1 _40514_ (.A1(_12751_),
    .A2(net865),
    .B1(_18492_),
    .Y(_05215_));
 sky130_fd_sc_hd__inv_1 _40515_ (.A(_18457_),
    .Y(_18493_));
 sky130_fd_sc_hd__o21ai_0 _40516_ (.A1(_18493_),
    .A2(net865),
    .B1(net2054),
    .Y(_18494_));
 sky130_fd_sc_hd__a21oi_1 _40517_ (.A1(_12759_),
    .A2(net865),
    .B1(_18494_),
    .Y(_05216_));
 sky130_fd_sc_hd__nand3_1 _40518_ (.A(_18343_),
    .B(_18321_),
    .C(_02736_),
    .Y(_18495_));
 sky130_fd_sc_hd__inv_1 _40520_ (.A(_18412_),
    .Y(_18497_));
 sky130_fd_sc_hd__nand3_1 _40521_ (.A(_18343_),
    .B(_18321_),
    .C(_02736_),
    .Y(_18498_));
 sky130_fd_sc_hd__o21ai_0 _40522_ (.A1(_18497_),
    .A2(_18498_),
    .B1(net2125),
    .Y(_18499_));
 sky130_fd_sc_hd__a21oi_1 _40523_ (.A1(_12766_),
    .A2(_18495_),
    .B1(_18499_),
    .Y(_05217_));
 sky130_fd_sc_hd__inv_1 _40524_ (.A(_18416_),
    .Y(_18500_));
 sky130_fd_sc_hd__o21ai_0 _40525_ (.A1(_18500_),
    .A2(_18498_),
    .B1(net2057),
    .Y(_18501_));
 sky130_fd_sc_hd__a21oi_1 _40526_ (.A1(_12773_),
    .A2(_18495_),
    .B1(_18501_),
    .Y(_05218_));
 sky130_fd_sc_hd__o21ai_0 _40527_ (.A1(_18425_),
    .A2(_18498_),
    .B1(net2055),
    .Y(_18502_));
 sky130_fd_sc_hd__a21oi_1 _40528_ (.A1(_12781_),
    .A2(_18495_),
    .B1(_18502_),
    .Y(_05219_));
 sky130_fd_sc_hd__o21ai_0 _40529_ (.A1(_18435_),
    .A2(_18498_),
    .B1(net2120),
    .Y(_18503_));
 sky130_fd_sc_hd__a21oi_1 _40530_ (.A1(_12790_),
    .A2(_18495_),
    .B1(_18503_),
    .Y(_05220_));
 sky130_fd_sc_hd__o21ai_0 _40532_ (.A1(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[1] ),
    .A2(_18481_),
    .B1(net2052),
    .Y(_18505_));
 sky130_fd_sc_hd__a21oi_1 _40533_ (.A1(_18416_),
    .A2(_18481_),
    .B1(_18505_),
    .Y(_05221_));
 sky130_fd_sc_hd__o21ai_0 _40534_ (.A1(_18441_),
    .A2(_18498_),
    .B1(net2125),
    .Y(_18506_));
 sky130_fd_sc_hd__a21oi_1 _40535_ (.A1(_12805_),
    .A2(_18495_),
    .B1(_18506_),
    .Y(_05222_));
 sky130_fd_sc_hd__o21ai_0 _40536_ (.A1(_18448_),
    .A2(_18498_),
    .B1(net2119),
    .Y(_18507_));
 sky130_fd_sc_hd__a21oi_1 _40537_ (.A1(_12812_),
    .A2(_18495_),
    .B1(_18507_),
    .Y(_05223_));
 sky130_fd_sc_hd__o21ai_0 _40538_ (.A1(_18452_),
    .A2(_18498_),
    .B1(net2120),
    .Y(_18508_));
 sky130_fd_sc_hd__a21oi_1 _40539_ (.A1(_12819_),
    .A2(_18495_),
    .B1(_18508_),
    .Y(_05224_));
 sky130_fd_sc_hd__o21ai_0 _40540_ (.A1(_18493_),
    .A2(_18495_),
    .B1(net2057),
    .Y(_18509_));
 sky130_fd_sc_hd__a21oi_1 _40541_ (.A1(_12826_),
    .A2(_18495_),
    .B1(_18509_),
    .Y(_05225_));
 sky130_fd_sc_hd__clkinv_1 _40542_ (.A(_18347_),
    .Y(_18510_));
 sky130_fd_sc_hd__o21ai_0 _40543_ (.A1(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[24] ),
    .A2(_18510_),
    .B1(net2052),
    .Y(_18511_));
 sky130_fd_sc_hd__a21oi_1 _40544_ (.A1(_18510_),
    .A2(_18412_),
    .B1(_18511_),
    .Y(_05226_));
 sky130_fd_sc_hd__o21ai_0 _40545_ (.A1(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[25] ),
    .A2(_18510_),
    .B1(net2051),
    .Y(_18512_));
 sky130_fd_sc_hd__a21oi_1 _40546_ (.A1(_18510_),
    .A2(_18416_),
    .B1(_18512_),
    .Y(_05227_));
 sky130_fd_sc_hd__nor2_1 _40547_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[26] ),
    .B(_18510_),
    .Y(_18513_));
 sky130_fd_sc_hd__o21ai_0 _40548_ (.A1(_18425_),
    .A2(_18347_),
    .B1(net2052),
    .Y(_18514_));
 sky130_fd_sc_hd__nor2_1 _40549_ (.A(_18513_),
    .B(_18514_),
    .Y(_05228_));
 sky130_fd_sc_hd__nor2_1 _40550_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[27] ),
    .B(_18510_),
    .Y(_18515_));
 sky130_fd_sc_hd__o21ai_0 _40551_ (.A1(_18435_),
    .A2(_18347_),
    .B1(net2051),
    .Y(_18516_));
 sky130_fd_sc_hd__nor2_1 _40552_ (.A(_18515_),
    .B(_18516_),
    .Y(_05229_));
 sky130_fd_sc_hd__nor2_1 _40553_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[28] ),
    .B(_18510_),
    .Y(_18517_));
 sky130_fd_sc_hd__o21ai_0 _40554_ (.A1(_18441_),
    .A2(_18347_),
    .B1(net2051),
    .Y(_18518_));
 sky130_fd_sc_hd__nor2_1 _40555_ (.A(_18517_),
    .B(_18518_),
    .Y(_05230_));
 sky130_fd_sc_hd__nor2_1 _40556_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[29] ),
    .B(_18510_),
    .Y(_18519_));
 sky130_fd_sc_hd__o21ai_0 _40557_ (.A1(_18448_),
    .A2(_18347_),
    .B1(net2051),
    .Y(_18520_));
 sky130_fd_sc_hd__nor2_1 _40558_ (.A(_18519_),
    .B(_18520_),
    .Y(_05231_));
 sky130_fd_sc_hd__o21ai_0 _40560_ (.A1(_18425_),
    .A2(net866),
    .B1(net2053),
    .Y(_18522_));
 sky130_fd_sc_hd__a21oi_1 _40561_ (.A1(_12878_),
    .A2(net866),
    .B1(_18522_),
    .Y(_05232_));
 sky130_fd_sc_hd__nor2_1 _40562_ (.A(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[30] ),
    .B(_18510_),
    .Y(_18523_));
 sky130_fd_sc_hd__o21ai_0 _40563_ (.A1(_18452_),
    .A2(_18347_),
    .B1(net2051),
    .Y(_18524_));
 sky130_fd_sc_hd__nor2_1 _40564_ (.A(_18523_),
    .B(_18524_),
    .Y(_05233_));
 sky130_fd_sc_hd__o21ai_0 _40565_ (.A1(_18493_),
    .A2(_18347_),
    .B1(net2054),
    .Y(_18525_));
 sky130_fd_sc_hd__a21oi_1 _40566_ (.A1(_12892_),
    .A2(_18347_),
    .B1(_18525_),
    .Y(_05234_));
 sky130_fd_sc_hd__o21ai_0 _40567_ (.A1(_18435_),
    .A2(net866),
    .B1(net2053),
    .Y(_18526_));
 sky130_fd_sc_hd__a21oi_1 _40568_ (.A1(_12899_),
    .A2(net866),
    .B1(_18526_),
    .Y(_05235_));
 sky130_fd_sc_hd__o21ai_0 _40570_ (.A1(_18441_),
    .A2(net866),
    .B1(net2053),
    .Y(_18528_));
 sky130_fd_sc_hd__a21oi_1 _40571_ (.A1(_12907_),
    .A2(net866),
    .B1(_18528_),
    .Y(_05236_));
 sky130_fd_sc_hd__o21ai_0 _40572_ (.A1(_18448_),
    .A2(_18480_),
    .B1(net2056),
    .Y(_18529_));
 sky130_fd_sc_hd__a21oi_1 _40573_ (.A1(_12914_),
    .A2(_18480_),
    .B1(_18529_),
    .Y(_05237_));
 sky130_fd_sc_hd__o21ai_0 _40574_ (.A1(_18452_),
    .A2(net866),
    .B1(net2053),
    .Y(_18530_));
 sky130_fd_sc_hd__a21oi_1 _40575_ (.A1(_12921_),
    .A2(_18480_),
    .B1(_18530_),
    .Y(_05238_));
 sky130_fd_sc_hd__o21ai_0 _40576_ (.A1(_18493_),
    .A2(net866),
    .B1(net2054),
    .Y(_18531_));
 sky130_fd_sc_hd__a21oi_1 _40577_ (.A1(_12928_),
    .A2(net866),
    .B1(_18531_),
    .Y(_05239_));
 sky130_fd_sc_hd__o21ai_0 _40578_ (.A1(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[8] ),
    .A2(_18487_),
    .B1(net2056),
    .Y(_18532_));
 sky130_fd_sc_hd__a21oi_1 _40579_ (.A1(_18412_),
    .A2(_18487_),
    .B1(_18532_),
    .Y(_05240_));
 sky130_fd_sc_hd__o21ai_0 _40580_ (.A1(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[9] ),
    .A2(_18487_),
    .B1(net2057),
    .Y(_18533_));
 sky130_fd_sc_hd__a21oi_1 _40581_ (.A1(_18416_),
    .A2(_18487_),
    .B1(_18533_),
    .Y(_05241_));
 sky130_fd_sc_hd__inv_1 _40582_ (.A(_18244_),
    .Y(_18534_));
 sky130_fd_sc_hd__nor2_1 _40583_ (.A(_18233_),
    .B(_18534_),
    .Y(_18535_));
 sky130_fd_sc_hd__nand2_1 _40585_ (.A(net828),
    .B(\inst$top.soc.spiflash.phy.deframer.cycle[0] ),
    .Y(_18537_));
 sky130_fd_sc_hd__o211ai_1 _40586_ (.A1(\inst$top.soc.spiflash.phy.deframer.cycle[0] ),
    .A2(_18234_),
    .B1(net2047),
    .C1(_18537_),
    .Y(_18538_));
 sky130_fd_sc_hd__inv_2 _40587_ (.A(_18538_),
    .Y(_05242_));
 sky130_fd_sc_hd__clkinv_1 _40588_ (.A(net828),
    .Y(_18539_));
 sky130_fd_sc_hd__nand2_1 _40589_ (.A(_18539_),
    .B(\inst$top.soc.spiflash.phy.deframer.cycle[1] ),
    .Y(_18540_));
 sky130_fd_sc_hd__nand3_1 _40590_ (.A(_18238_),
    .B(_02750_),
    .C(_18234_),
    .Y(_18541_));
 sky130_fd_sc_hd__a21oi_1 _40591_ (.A1(_18540_),
    .A2(_18541_),
    .B1(net2947),
    .Y(_05243_));
 sky130_fd_sc_hd__nand2_1 _40592_ (.A(net828),
    .B(_02749_),
    .Y(_18542_));
 sky130_fd_sc_hd__nand2_1 _40593_ (.A(_18542_),
    .B(_18214_),
    .Y(_18543_));
 sky130_fd_sc_hd__nand4_1 _40594_ (.A(_18543_),
    .B(net2048),
    .C(_18344_),
    .D(_18426_),
    .Y(_18544_));
 sky130_fd_sc_hd__a31oi_1 _40595_ (.A1(\inst$top.soc.spiflash.phy.deframer.cycle[2] ),
    .A2(_02749_),
    .A3(net828),
    .B1(_18544_),
    .Y(_05244_));
 sky130_fd_sc_hd__o21ai_0 _40596_ (.A1(\inst$top.soc.spiflash.phy.deframer.data_reg[0] ),
    .A2(_18535_),
    .B1(net2047),
    .Y(_18545_));
 sky130_fd_sc_hd__a21oi_1 _40597_ (.A1(_18412_),
    .A2(net828),
    .B1(_18545_),
    .Y(_05245_));
 sky130_fd_sc_hd__o21ai_0 _40598_ (.A1(\inst$top.soc.spiflash.phy.deframer.data_reg[1] ),
    .A2(net828),
    .B1(net2048),
    .Y(_18546_));
 sky130_fd_sc_hd__a21oi_1 _40599_ (.A1(_18416_),
    .A2(net828),
    .B1(_18546_),
    .Y(_05246_));
 sky130_fd_sc_hd__o21ai_0 _40600_ (.A1(_18425_),
    .A2(_18539_),
    .B1(net2047),
    .Y(_18547_));
 sky130_fd_sc_hd__a21oi_1 _40601_ (.A1(_18429_),
    .A2(_18539_),
    .B1(_18547_),
    .Y(_05247_));
 sky130_fd_sc_hd__o21ai_0 _40602_ (.A1(_18435_),
    .A2(_18539_),
    .B1(net2047),
    .Y(_18548_));
 sky130_fd_sc_hd__a21oi_1 _40603_ (.A1(_18438_),
    .A2(_18539_),
    .B1(_18548_),
    .Y(_05248_));
 sky130_fd_sc_hd__nor2_1 _40604_ (.A(_18441_),
    .B(_18539_),
    .Y(_18549_));
 sky130_fd_sc_hd__o21ai_0 _40605_ (.A1(\inst$top.soc.spiflash.phy.deframer.data_reg[4] ),
    .A2(net828),
    .B1(net2047),
    .Y(_18550_));
 sky130_fd_sc_hd__nor2_1 _40606_ (.A(_18549_),
    .B(_18550_),
    .Y(_05249_));
 sky130_fd_sc_hd__nor2_1 _40607_ (.A(_18448_),
    .B(_18539_),
    .Y(_18551_));
 sky130_fd_sc_hd__o21ai_0 _40608_ (.A1(\inst$top.soc.spiflash.phy.deframer.data_reg[5] ),
    .A2(net828),
    .B1(net2047),
    .Y(_18552_));
 sky130_fd_sc_hd__nor2_1 _40609_ (.A(_18551_),
    .B(_18552_),
    .Y(_05250_));
 sky130_fd_sc_hd__nor2_1 _40610_ (.A(_18452_),
    .B(_18539_),
    .Y(_18553_));
 sky130_fd_sc_hd__o21ai_0 _40611_ (.A1(\inst$top.soc.spiflash.phy.deframer.data_reg[6] ),
    .A2(net828),
    .B1(net2048),
    .Y(_18554_));
 sky130_fd_sc_hd__nor2_1 _40612_ (.A(_18553_),
    .B(_18554_),
    .Y(_05251_));
 sky130_fd_sc_hd__inv_1 _40613_ (.A(_18274_),
    .Y(_18555_));
 sky130_fd_sc_hd__a21oi_1 _40615_ (.A1(_18300_),
    .A2(_18555_),
    .B1(net2579),
    .Y(_18557_));
 sky130_fd_sc_hd__a211oi_2 _40616_ (.A1(net2579),
    .A2(_18555_),
    .B1(net2944),
    .C1(_18557_),
    .Y(_05252_));
 sky130_fd_sc_hd__nand3_1 _40617_ (.A(_18300_),
    .B(_02747_),
    .C(_18555_),
    .Y(_18558_));
 sky130_fd_sc_hd__nand2_1 _40618_ (.A(_18274_),
    .B(net2578),
    .Y(_18559_));
 sky130_fd_sc_hd__a21oi_1 _40619_ (.A1(_18558_),
    .A2(_18559_),
    .B1(net2944),
    .Y(_05253_));
 sky130_fd_sc_hd__nand2_1 _40620_ (.A(_18555_),
    .B(_02748_),
    .Y(_18560_));
 sky130_fd_sc_hd__nand2_1 _40621_ (.A(_18560_),
    .B(\inst$top.soc.spiflash.phy.enframer.cycle[2] ),
    .Y(_18561_));
 sky130_fd_sc_hd__nand3_1 _40622_ (.A(_18555_),
    .B(_18204_),
    .C(_02748_),
    .Y(_18562_));
 sky130_fd_sc_hd__a211oi_2 _40623_ (.A1(_18561_),
    .A2(_18562_),
    .B1(net2944),
    .C1(_18381_),
    .Y(_05254_));
 sky130_fd_sc_hd__nor2_1 _40624_ (.A(_18258_),
    .B(_18255_),
    .Y(_18563_));
 sky130_fd_sc_hd__nand2_1 _40625_ (.A(_18563_),
    .B(_18376_),
    .Y(_18564_));
 sky130_fd_sc_hd__inv_1 _40626_ (.A(_18376_),
    .Y(_18565_));
 sky130_fd_sc_hd__o21ai_0 _40627_ (.A1(_18565_),
    .A2(_18245_),
    .B1(\inst$top.soc.spiflash.phy.io_clocker.fsm_state ),
    .Y(_18566_));
 sky130_fd_sc_hd__a21oi_1 _40628_ (.A1(_18564_),
    .A2(_18566_),
    .B1(net2947),
    .Y(_05255_));
 sky130_fd_sc_hd__inv_1 _40629_ (.A(_18563_),
    .Y(_18567_));
 sky130_fd_sc_hd__nand2_1 _40630_ (.A(_18246_),
    .B(\inst$top.soc.spiflash.phy.io_clocker.fsm_state ),
    .Y(_18568_));
 sky130_fd_sc_hd__nand2_1 _40631_ (.A(_18568_),
    .B(_18273_),
    .Y(_18569_));
 sky130_fd_sc_hd__inv_1 _40632_ (.A(_18569_),
    .Y(_18570_));
 sky130_fd_sc_hd__nand2_2 _40633_ (.A(_18567_),
    .B(_18570_),
    .Y(_18571_));
 sky130_fd_sc_hd__nand2_1 _40634_ (.A(_18571_),
    .B(_02739_),
    .Y(_18572_));
 sky130_fd_sc_hd__nand3_1 _40635_ (.A(_18567_),
    .B(_18570_),
    .C(\inst$top.soc.spiflash.phy.io_clocker.timer[0] ),
    .Y(_18573_));
 sky130_fd_sc_hd__a21oi_2 _40636_ (.A1(_18571_),
    .A2(_18273_),
    .B1(net2932),
    .Y(_18574_));
 sky130_fd_sc_hd__inv_1 _40637_ (.A(_18574_),
    .Y(_18575_));
 sky130_fd_sc_hd__a21oi_2 _40638_ (.A1(_18572_),
    .A2(_18573_),
    .B1(_18575_),
    .Y(_05256_));
 sky130_fd_sc_hd__nand3_1 _40639_ (.A(_18568_),
    .B(_18258_),
    .C(_18376_),
    .Y(_18576_));
 sky130_fd_sc_hd__nor2_1 _40640_ (.A(_18261_),
    .B(_18355_),
    .Y(_18577_));
 sky130_fd_sc_hd__nor2_1 _40641_ (.A(\inst$top.soc.spiflash.phy.io_clocker.fsm_state ),
    .B(_18565_),
    .Y(_18578_));
 sky130_fd_sc_hd__nand2_1 _40642_ (.A(_18255_),
    .B(_18578_),
    .Y(_18579_));
 sky130_fd_sc_hd__nand3_1 _40643_ (.A(_18576_),
    .B(_18577_),
    .C(_18579_),
    .Y(_18580_));
 sky130_fd_sc_hd__nor3_1 _40644_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[9] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[8] ),
    .C(_18580_),
    .Y(_18581_));
 sky130_fd_sc_hd__o21ai_0 _40645_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[10] ),
    .A2(_18581_),
    .B1(_18574_),
    .Y(_18582_));
 sky130_fd_sc_hd__a21oi_1 _40646_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[10] ),
    .A2(_18581_),
    .B1(_18582_),
    .Y(_05257_));
 sky130_fd_sc_hd__nor2_1 _40647_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[7] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[8] ),
    .Y(_18583_));
 sky130_fd_sc_hd__inv_1 _40648_ (.A(_18583_),
    .Y(_18584_));
 sky130_fd_sc_hd__nor2_1 _40649_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[2] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[1] ),
    .Y(_18585_));
 sky130_fd_sc_hd__inv_1 _40650_ (.A(_18585_),
    .Y(_18586_));
 sky130_fd_sc_hd__nor3_1 _40651_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[3] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[4] ),
    .C(_18586_),
    .Y(_18587_));
 sky130_fd_sc_hd__inv_1 _40652_ (.A(_18587_),
    .Y(_18588_));
 sky130_fd_sc_hd__nor4_1 _40653_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[5] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[6] ),
    .C(_18584_),
    .D(_18588_),
    .Y(_18589_));
 sky130_fd_sc_hd__nand3_1 _40654_ (.A(_18571_),
    .B(_02739_),
    .C(_18589_),
    .Y(_18590_));
 sky130_fd_sc_hd__nor3_1 _40655_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[9] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[10] ),
    .C(_18590_),
    .Y(_18591_));
 sky130_fd_sc_hd__o21ai_0 _40656_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[11] ),
    .A2(_18591_),
    .B1(_18574_),
    .Y(_18592_));
 sky130_fd_sc_hd__a21oi_1 _40657_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[11] ),
    .A2(_18591_),
    .B1(_18592_),
    .Y(_05258_));
 sky130_fd_sc_hd__nor2_1 _40658_ (.A(_18268_),
    .B(_18580_),
    .Y(_18593_));
 sky130_fd_sc_hd__o21ai_0 _40659_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[12] ),
    .A2(_18593_),
    .B1(_18574_),
    .Y(_18594_));
 sky130_fd_sc_hd__a21oi_1 _40660_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[12] ),
    .A2(_18593_),
    .B1(_18594_),
    .Y(_05259_));
 sky130_fd_sc_hd__inv_1 _40661_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[13] ),
    .Y(_18595_));
 sky130_fd_sc_hd__nor2_1 _40662_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[11] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[12] ),
    .Y(_18596_));
 sky130_fd_sc_hd__nand2_1 _40663_ (.A(_18591_),
    .B(_18596_),
    .Y(_18597_));
 sky130_fd_sc_hd__o21bai_1 _40664_ (.A1(_18595_),
    .A2(_18597_),
    .B1_N(_18575_),
    .Y(_18598_));
 sky130_fd_sc_hd__a21oi_2 _40665_ (.A1(_18595_),
    .A2(_18597_),
    .B1(_18598_),
    .Y(_05260_));
 sky130_fd_sc_hd__nand3_1 _40666_ (.A(_18266_),
    .B(_18267_),
    .C(_18263_),
    .Y(_18599_));
 sky130_fd_sc_hd__nor2_1 _40667_ (.A(_18599_),
    .B(_18580_),
    .Y(_18600_));
 sky130_fd_sc_hd__o21ai_0 _40668_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[14] ),
    .A2(_18600_),
    .B1(_18574_),
    .Y(_18601_));
 sky130_fd_sc_hd__a21oi_1 _40669_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[14] ),
    .A2(_18600_),
    .B1(_18601_),
    .Y(_05261_));
 sky130_fd_sc_hd__inv_1 _40670_ (.A(_18590_),
    .Y(_18602_));
 sky130_fd_sc_hd__nor2_1 _40671_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[9] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[10] ),
    .Y(_18603_));
 sky130_fd_sc_hd__nor3_1 _40672_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[11] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[14] ),
    .C(_18264_),
    .Y(_18604_));
 sky130_fd_sc_hd__nand3_1 _40673_ (.A(_18602_),
    .B(_18603_),
    .C(_18604_),
    .Y(_18605_));
 sky130_fd_sc_hd__o21ai_0 _40674_ (.A1(_18270_),
    .A2(_18605_),
    .B1(_18574_),
    .Y(_18606_));
 sky130_fd_sc_hd__a21oi_1 _40675_ (.A1(_18270_),
    .A2(_18605_),
    .B1(_18606_),
    .Y(_05262_));
 sky130_fd_sc_hd__nor2_1 _40676_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[1] ),
    .B(_18571_),
    .Y(_18607_));
 sky130_fd_sc_hd__a211oi_2 _40677_ (.A1(_02742_),
    .A2(_18571_),
    .B1(_18607_),
    .C1(_18575_),
    .Y(_05263_));
 sky130_fd_sc_hd__a21oi_1 _40678_ (.A1(_18571_),
    .A2(_02741_),
    .B1(\inst$top.soc.spiflash.phy.io_clocker.timer[2] ),
    .Y(_18608_));
 sky130_fd_sc_hd__a211oi_2 _40679_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[2] ),
    .A2(_02741_),
    .B1(_18608_),
    .C1(_18575_),
    .Y(_05264_));
 sky130_fd_sc_hd__nor2_1 _40680_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[0] ),
    .B(_18586_),
    .Y(_18609_));
 sky130_fd_sc_hd__xnor2_1 _40681_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[3] ),
    .B(_18609_),
    .Y(_18610_));
 sky130_fd_sc_hd__nor3_1 _40682_ (.A(net2932),
    .B(_18610_),
    .C(_18359_),
    .Y(_05265_));
 sky130_fd_sc_hd__xnor2_1 _40683_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[4] ),
    .B(_18354_),
    .Y(_18611_));
 sky130_fd_sc_hd__nor3_1 _40684_ (.A(net2932),
    .B(_18611_),
    .C(_18359_),
    .Y(_05266_));
 sky130_fd_sc_hd__nor2_1 _40685_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[0] ),
    .B(_18588_),
    .Y(_18612_));
 sky130_fd_sc_hd__nor4_1 _40686_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[3] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[4] ),
    .C(_18586_),
    .D(_18572_),
    .Y(_18613_));
 sky130_fd_sc_hd__o21ai_0 _40687_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[5] ),
    .A2(_18613_),
    .B1(_18574_),
    .Y(_18614_));
 sky130_fd_sc_hd__a21oi_2 _40688_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[5] ),
    .A2(_18612_),
    .B1(_18614_),
    .Y(_05267_));
 sky130_fd_sc_hd__nand3_1 _40689_ (.A(_18260_),
    .B(_18271_),
    .C(_02741_),
    .Y(_18615_));
 sky130_fd_sc_hd__xor2_1 _40690_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[6] ),
    .B(_18615_),
    .X(_18616_));
 sky130_fd_sc_hd__nor3_1 _40691_ (.A(net2932),
    .B(_18616_),
    .C(_18359_),
    .Y(_05268_));
 sky130_fd_sc_hd__inv_1 _40692_ (.A(_18612_),
    .Y(_18617_));
 sky130_fd_sc_hd__nor3_1 _40693_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[5] ),
    .B(\inst$top.soc.spiflash.phy.io_clocker.timer[6] ),
    .C(_18617_),
    .Y(_18618_));
 sky130_fd_sc_hd__a21oi_1 _40694_ (.A1(_18571_),
    .A2(_18618_),
    .B1(\inst$top.soc.spiflash.phy.io_clocker.timer[7] ),
    .Y(_18619_));
 sky130_fd_sc_hd__a211oi_2 _40695_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[7] ),
    .A2(_18618_),
    .B1(_18619_),
    .C1(_18575_),
    .Y(_05269_));
 sky130_fd_sc_hd__inv_1 _40696_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[8] ),
    .Y(_18620_));
 sky130_fd_sc_hd__nand2_1 _40697_ (.A(_18580_),
    .B(_18620_),
    .Y(_18621_));
 sky130_fd_sc_hd__nand2_1 _40698_ (.A(_18574_),
    .B(_18621_),
    .Y(_18622_));
 sky130_fd_sc_hd__a21oi_1 _40699_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[8] ),
    .A2(_18577_),
    .B1(_18622_),
    .Y(_05270_));
 sky130_fd_sc_hd__o21ai_0 _40700_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[9] ),
    .A2(_18602_),
    .B1(_18574_),
    .Y(_18623_));
 sky130_fd_sc_hd__a21oi_1 _40701_ (.A1(\inst$top.soc.spiflash.phy.io_clocker.timer[9] ),
    .A2(_18602_),
    .B1(_18623_),
    .Y(_05271_));
 sky130_fd_sc_hd__a211oi_1 _40702_ (.A1(_18240_),
    .A2(_18209_),
    .B1(net2944),
    .C1(_18274_),
    .Y(_05272_));
 sky130_fd_sc_hd__nor2_1 _40703_ (.A(net2947),
    .B(_18291_),
    .Y(_05273_));
 sky130_fd_sc_hd__nand2_1 _40704_ (.A(_18289_),
    .B(net2047),
    .Y(_18624_));
 sky130_fd_sc_hd__inv_2 _40705_ (.A(_18624_),
    .Y(_05274_));
 sky130_fd_sc_hd__o21ai_0 _40706_ (.A1(_18281_),
    .A2(_18282_),
    .B1(net2049),
    .Y(_18625_));
 sky130_fd_sc_hd__inv_2 _40707_ (.A(_18625_),
    .Y(_05275_));
 sky130_fd_sc_hd__inv_1 _40708_ (.A(_18377_),
    .Y(_18626_));
 sky130_fd_sc_hd__o21ai_0 _40709_ (.A1(\inst$top.soc.spiflash.phy.io_streamer.o_latch.sck.o ),
    .A2(_18626_),
    .B1(_18564_),
    .Y(_18627_));
 sky130_fd_sc_hd__inv_2 _40710_ (.A(_18627_),
    .Y(\inst$top.soc.spiflash.phy.io_streamer.buffer_sck.o ));
 sky130_fd_sc_hd__nand2_1 _40711_ (.A(_18627_),
    .B(net2027),
    .Y(_05276_));
 sky130_fd_sc_hd__nand3_1 _40712_ (.A(_18246_),
    .B(_18254_),
    .C(_18359_),
    .Y(_18628_));
 sky130_fd_sc_hd__nand2_1 _40714_ (.A(net806),
    .B(\inst$top.soc.spiflash.phy.io_streamer.o_latch.cs.o ),
    .Y(_18630_));
 sky130_fd_sc_hd__o21ai_2 _40715_ (.A1(_18211_),
    .A2(net806),
    .B1(_18630_),
    .Y(\inst$top.soc.spiflash.phy.io_streamer.buffer_cs.o ));
 sky130_fd_sc_hd__inv_1 _40716_ (.A(\inst$top.soc.spiflash.phy.io_streamer.buffer_cs.o ),
    .Y(_18631_));
 sky130_fd_sc_hd__nor2_1 _40717_ (.A(net2932),
    .B(_18631_),
    .Y(_05277_));
 sky130_fd_sc_hd__nor2_1 _40718_ (.A(\inst$top.soc.spiflash.ctrl.o_addr_count[0] ),
    .B(\inst$top.soc.spiflash.ctrl.o_addr_count[1] ),
    .Y(_18632_));
 sky130_fd_sc_hd__inv_1 _40719_ (.A(_18632_),
    .Y(_18633_));
 sky130_fd_sc_hd__nor2_1 _40720_ (.A(\inst$top.soc.spiflash.ctrl.o_addr_count[0] ),
    .B(_02724_),
    .Y(_18634_));
 sky130_fd_sc_hd__nand2_1 _40721_ (.A(_09329_),
    .B(_18634_),
    .Y(_18635_));
 sky130_fd_sc_hd__nand2_1 _40722_ (.A(_02724_),
    .B(\inst$top.soc.spiflash.ctrl.o_addr_count[0] ),
    .Y(_18636_));
 sky130_fd_sc_hd__inv_1 _40723_ (.A(_18636_),
    .Y(_18637_));
 sky130_fd_sc_hd__nand2_1 _40724_ (.A(_09283_),
    .B(_18637_),
    .Y(_18638_));
 sky130_fd_sc_hd__o211ai_1 _40725_ (.A1(_18633_),
    .A2(_17868_),
    .B1(_18635_),
    .C1(_18638_),
    .Y(_18639_));
 sky130_fd_sc_hd__o21ai_0 _40726_ (.A1(_18465_),
    .A2(_18209_),
    .B1(_18317_),
    .Y(_18640_));
 sky130_fd_sc_hd__a21oi_1 _40727_ (.A1(_18639_),
    .A2(net1638),
    .B1(_18640_),
    .Y(_18641_));
 sky130_fd_sc_hd__inv_1 _40728_ (.A(_18641_),
    .Y(_18642_));
 sky130_fd_sc_hd__nor2_1 _40729_ (.A(_02744_),
    .B(_18642_),
    .Y(_18643_));
 sky130_fd_sc_hd__nor3_1 _40730_ (.A(\inst$top.soc.spiflash.ctrl.o_addr_count[0] ),
    .B(_02724_),
    .C(_09330_),
    .Y(_18644_));
 sky130_fd_sc_hd__o22ai_1 _40731_ (.A1(_18636_),
    .A2(_09285_),
    .B1(_19850_),
    .B2(_18633_),
    .Y(_18645_));
 sky130_fd_sc_hd__o21ai_0 _40732_ (.A1(_18644_),
    .A2(_18645_),
    .B1(net1638),
    .Y(_18646_));
 sky130_fd_sc_hd__a21oi_1 _40733_ (.A1(_18276_),
    .A2(_18280_),
    .B1(_18195_),
    .Y(_18647_));
 sky130_fd_sc_hd__a211oi_1 _40734_ (.A1(\inst$top.soc.spiflash.ctrl.raw_tx_data[3] ),
    .A2(_18208_),
    .B1(_18316_),
    .C1(_18647_),
    .Y(_18648_));
 sky130_fd_sc_hd__nand2_1 _40735_ (.A(_18646_),
    .B(_18648_),
    .Y(_18649_));
 sky130_fd_sc_hd__inv_1 _40736_ (.A(_18649_),
    .Y(_18650_));
 sky130_fd_sc_hd__nand2_1 _40737_ (.A(_18650_),
    .B(_02744_),
    .Y(_18651_));
 sky130_fd_sc_hd__nand2_1 _40738_ (.A(_18651_),
    .B(_02745_),
    .Y(_18652_));
 sky130_fd_sc_hd__nand2_1 _40739_ (.A(_09290_),
    .B(_18634_),
    .Y(_18653_));
 sky130_fd_sc_hd__nand2_1 _40740_ (.A(\inst$top.soc.bus__adr[7] ),
    .B(_18637_),
    .Y(_18654_));
 sky130_fd_sc_hd__nand3_1 _40741_ (.A(_09298_),
    .B(\inst$top.soc.spiflash.ctrl.o_addr_count[0] ),
    .C(\inst$top.soc.spiflash.ctrl.o_addr_count[1] ),
    .Y(_18655_));
 sky130_fd_sc_hd__nand3_1 _40742_ (.A(_18653_),
    .B(_18654_),
    .C(_18655_),
    .Y(_18656_));
 sky130_fd_sc_hd__nand2_1 _40743_ (.A(_18195_),
    .B(_18317_),
    .Y(_18657_));
 sky130_fd_sc_hd__a221oi_1 _40744_ (.A1(\inst$top.soc.spiflash.ctrl.raw_tx_data[1] ),
    .A2(_18208_),
    .B1(_18656_),
    .B2(_18327_),
    .C1(_18657_),
    .Y(_18658_));
 sky130_fd_sc_hd__nand2_1 _40745_ (.A(_18658_),
    .B(_02744_),
    .Y(_18659_));
 sky130_fd_sc_hd__nand2_1 _40746_ (.A(_09292_),
    .B(_18634_),
    .Y(_18660_));
 sky130_fd_sc_hd__o21ai_0 _40747_ (.A1(_19859_),
    .A2(_18636_),
    .B1(_18660_),
    .Y(_18661_));
 sky130_fd_sc_hd__nor3_1 _40748_ (.A(_02723_),
    .B(_02724_),
    .C(_17834_),
    .Y(_18662_));
 sky130_fd_sc_hd__o21ai_0 _40749_ (.A1(_18661_),
    .A2(_18662_),
    .B1(net1638),
    .Y(_18663_));
 sky130_fd_sc_hd__a21oi_1 _40750_ (.A1(\inst$top.soc.spiflash.ctrl.raw_tx_data[0] ),
    .A2(_18208_),
    .B1(_18657_),
    .Y(_18664_));
 sky130_fd_sc_hd__nand3_1 _40751_ (.A(_18663_),
    .B(net2579),
    .C(_18664_),
    .Y(_18665_));
 sky130_fd_sc_hd__nand3_1 _40752_ (.A(_18659_),
    .B(net2578),
    .C(_18665_),
    .Y(_18666_));
 sky130_fd_sc_hd__o211ai_1 _40753_ (.A1(_18643_),
    .A2(_18652_),
    .B1(\inst$top.soc.spiflash.phy.enframer.cycle[2] ),
    .C1(_18666_),
    .Y(_18667_));
 sky130_fd_sc_hd__nand2_1 _40754_ (.A(_09261_),
    .B(_18634_),
    .Y(_18668_));
 sky130_fd_sc_hd__nand2_1 _40755_ (.A(_09321_),
    .B(_18637_),
    .Y(_18669_));
 sky130_fd_sc_hd__nand2_1 _40756_ (.A(\inst$top.soc.bus__adr[3] ),
    .B(_18632_),
    .Y(_18670_));
 sky130_fd_sc_hd__nand3_1 _40757_ (.A(_18668_),
    .B(_18669_),
    .C(_18670_),
    .Y(_18671_));
 sky130_fd_sc_hd__o21ai_0 _40758_ (.A1(_18276_),
    .A2(_18195_),
    .B1(_18317_),
    .Y(_18672_));
 sky130_fd_sc_hd__nor2_1 _40759_ (.A(_18471_),
    .B(_18209_),
    .Y(_18673_));
 sky130_fd_sc_hd__a211oi_1 _40760_ (.A1(_18671_),
    .A2(net1638),
    .B1(_18672_),
    .C1(_18673_),
    .Y(_18674_));
 sky130_fd_sc_hd__nand2_1 _40761_ (.A(_18674_),
    .B(_02744_),
    .Y(_18675_));
 sky130_fd_sc_hd__nand2_1 _40762_ (.A(_09259_),
    .B(_18634_),
    .Y(_18676_));
 sky130_fd_sc_hd__o221ai_1 _40763_ (.A1(_18636_),
    .A2(_09316_),
    .B1(_18633_),
    .B2(_19868_),
    .C1(_18676_),
    .Y(_18677_));
 sky130_fd_sc_hd__nand2_1 _40764_ (.A(_18677_),
    .B(net1638),
    .Y(_18678_));
 sky130_fd_sc_hd__a221oi_1 _40765_ (.A1(_18194_),
    .A2(_18277_),
    .B1(_18208_),
    .B2(\inst$top.soc.spiflash.ctrl.raw_tx_data[4] ),
    .C1(_18316_),
    .Y(_18679_));
 sky130_fd_sc_hd__nand3_1 _40766_ (.A(_18678_),
    .B(net2579),
    .C(_18679_),
    .Y(_18680_));
 sky130_fd_sc_hd__nand3_1 _40767_ (.A(_18675_),
    .B(net2578),
    .C(_18680_),
    .Y(_18681_));
 sky130_fd_sc_hd__nand3_1 _40768_ (.A(_18194_),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[1] ),
    .C(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[0] ),
    .Y(_18682_));
 sky130_fd_sc_hd__nand2_1 _40769_ (.A(_09268_),
    .B(_18634_),
    .Y(_18683_));
 sky130_fd_sc_hd__nand2_1 _40770_ (.A(_09324_),
    .B(_18637_),
    .Y(_18684_));
 sky130_fd_sc_hd__nand2_1 _40771_ (.A(\inst$top.soc.bus__adr[4] ),
    .B(_18632_),
    .Y(_18685_));
 sky130_fd_sc_hd__nand3_1 _40772_ (.A(_18683_),
    .B(_18684_),
    .C(_18685_),
    .Y(_18686_));
 sky130_fd_sc_hd__nand2_1 _40773_ (.A(_18686_),
    .B(net1638),
    .Y(_18687_));
 sky130_fd_sc_hd__o2111ai_1 _40774_ (.A1(_18473_),
    .A2(_18209_),
    .B1(_18317_),
    .C1(_18682_),
    .D1(_18687_),
    .Y(_18688_));
 sky130_fd_sc_hd__a21oi_1 _40775_ (.A1(\inst$top.soc.spiflash.ctrl.raw_tx_data[7] ),
    .A2(_18208_),
    .B1(_18672_),
    .Y(_18689_));
 sky130_fd_sc_hd__nand2_1 _40776_ (.A(_09265_),
    .B(_18634_),
    .Y(_18690_));
 sky130_fd_sc_hd__nand2_1 _40777_ (.A(_09314_),
    .B(_18637_),
    .Y(_18691_));
 sky130_fd_sc_hd__nand2_1 _40778_ (.A(\inst$top.soc.bus__adr[5] ),
    .B(_18632_),
    .Y(_18692_));
 sky130_fd_sc_hd__nand3_1 _40779_ (.A(_18690_),
    .B(_18691_),
    .C(_18692_),
    .Y(_18693_));
 sky130_fd_sc_hd__nand2_1 _40780_ (.A(_18693_),
    .B(net1638),
    .Y(_18694_));
 sky130_fd_sc_hd__nand3_1 _40781_ (.A(_18689_),
    .B(_02744_),
    .C(_18694_),
    .Y(_18695_));
 sky130_fd_sc_hd__o211ai_1 _40782_ (.A1(_02744_),
    .A2(_18688_),
    .B1(_02745_),
    .C1(_18695_),
    .Y(_18696_));
 sky130_fd_sc_hd__nand3_1 _40783_ (.A(_18681_),
    .B(_18204_),
    .C(_18696_),
    .Y(_18697_));
 sky130_fd_sc_hd__nand2_1 _40784_ (.A(_18283_),
    .B(_18289_),
    .Y(_18698_));
 sky130_fd_sc_hd__inv_1 _40785_ (.A(_18698_),
    .Y(_18699_));
 sky130_fd_sc_hd__nor2_1 _40786_ (.A(_18290_),
    .B(_18699_),
    .Y(_18700_));
 sky130_fd_sc_hd__nor2_1 _40787_ (.A(net2579),
    .B(_18688_),
    .Y(_18701_));
 sky130_fd_sc_hd__nand2_1 _40788_ (.A(_18287_),
    .B(_02745_),
    .Y(_18702_));
 sky130_fd_sc_hd__inv_1 _40789_ (.A(_18702_),
    .Y(_18703_));
 sky130_fd_sc_hd__nand2_1 _40790_ (.A(_18680_),
    .B(_18703_),
    .Y(_18704_));
 sky130_fd_sc_hd__o211ai_1 _40791_ (.A1(net2579),
    .A2(_18642_),
    .B1(net2578),
    .C1(_18287_),
    .Y(_18705_));
 sky130_fd_sc_hd__nand3_1 _40792_ (.A(_18678_),
    .B(_02744_),
    .C(_18679_),
    .Y(_18706_));
 sky130_fd_sc_hd__nor2_1 _40793_ (.A(net2578),
    .B(_18284_),
    .Y(_18707_));
 sky130_fd_sc_hd__nand2_1 _40794_ (.A(_18706_),
    .B(_18707_),
    .Y(_18708_));
 sky130_fd_sc_hd__nand2_1 _40795_ (.A(_18705_),
    .B(_18708_),
    .Y(_18709_));
 sky130_fd_sc_hd__nand2_1 _40796_ (.A(_18709_),
    .B(_18665_),
    .Y(_18710_));
 sky130_fd_sc_hd__o21ai_0 _40797_ (.A1(_18701_),
    .A2(_18704_),
    .B1(_18710_),
    .Y(_18711_));
 sky130_fd_sc_hd__a32o_1 _40798_ (.A1(_18667_),
    .A2(_18697_),
    .A3(_18700_),
    .B1(_18711_),
    .B2(_18204_),
    .X(_18712_));
 sky130_fd_sc_hd__inv_1 _40799_ (.A(net806),
    .Y(_18713_));
 sky130_fd_sc_hd__nand2_1 _40800_ (.A(_18712_),
    .B(_18713_),
    .Y(_18714_));
 sky130_fd_sc_hd__nand2_1 _40801_ (.A(net806),
    .B(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io0.o ),
    .Y(_18715_));
 sky130_fd_sc_hd__nand2_1 _40802_ (.A(_18714_),
    .B(_18715_),
    .Y(\inst$top.soc.spiflash.phy.io_streamer.buffer_io0.o ));
 sky130_fd_sc_hd__a21oi_1 _40803_ (.A1(_18714_),
    .A2(_18715_),
    .B1(net2954),
    .Y(_05278_));
 sky130_fd_sc_hd__nor2_1 _40804_ (.A(_18210_),
    .B(_18699_),
    .Y(_18716_));
 sky130_fd_sc_hd__nand2_1 _40805_ (.A(net806),
    .B(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io0.oe ),
    .Y(_18717_));
 sky130_fd_sc_hd__o21ai_1 _40806_ (.A1(_18716_),
    .A2(net806),
    .B1(_18717_),
    .Y(\inst$top.soc.spiflash.phy.io_streamer.buffer_io0.oe ));
 sky130_fd_sc_hd__inv_1 _40807_ (.A(\inst$top.soc.spiflash.phy.io_streamer.buffer_io0.oe ),
    .Y(_18718_));
 sky130_fd_sc_hd__nor2_1 _40808_ (.A(net2933),
    .B(_18718_),
    .Y(_05279_));
 sky130_fd_sc_hd__inv_1 _40809_ (.A(_18695_),
    .Y(_18719_));
 sky130_fd_sc_hd__a211oi_1 _40810_ (.A1(_18674_),
    .A2(net2579),
    .B1(_18702_),
    .C1(_18719_),
    .Y(_18720_));
 sky130_fd_sc_hd__nand3_1 _40811_ (.A(_18651_),
    .B(net2578),
    .C(_18287_),
    .Y(_18721_));
 sky130_fd_sc_hd__nand2_1 _40812_ (.A(_18675_),
    .B(_18707_),
    .Y(_18722_));
 sky130_fd_sc_hd__a22oi_1 _40813_ (.A1(_18658_),
    .A2(net2579),
    .B1(_18721_),
    .B2(_18722_),
    .Y(_18723_));
 sky130_fd_sc_hd__o21ai_0 _40814_ (.A1(_18720_),
    .A2(_18723_),
    .B1(_18204_),
    .Y(_18724_));
 sky130_fd_sc_hd__or2_2 _40815_ (.A(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io1.o ),
    .B(_18626_),
    .X(_18725_));
 sky130_fd_sc_hd__inv_1 _40816_ (.A(_18725_),
    .Y(_18726_));
 sky130_fd_sc_hd__a21oi_1 _40817_ (.A1(_18626_),
    .A2(_18724_),
    .B1(_18726_),
    .Y(\inst$top.soc.spiflash.phy.io_streamer.buffer_io1.o ));
 sky130_fd_sc_hd__a211oi_2 _40818_ (.A1(_18626_),
    .A2(_18724_),
    .B1(net2944),
    .C1(_18726_),
    .Y(_05280_));
 sky130_fd_sc_hd__o21ai_0 _40819_ (.A1(_18281_),
    .A2(_18287_),
    .B1(_18713_),
    .Y(_18727_));
 sky130_fd_sc_hd__nand2_1 _40820_ (.A(net806),
    .B(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io1.oe ),
    .Y(_18728_));
 sky130_fd_sc_hd__nand2_1 _40821_ (.A(_18727_),
    .B(_18728_),
    .Y(\inst$top.soc.spiflash.phy.io_streamer.buffer_io1.oe ));
 sky130_fd_sc_hd__a21oi_1 _40822_ (.A1(_18727_),
    .A2(_18728_),
    .B1(net2932),
    .Y(_05281_));
 sky130_fd_sc_hd__nor2_1 _40823_ (.A(\inst$top.soc.spiflash.phy.enframer.cycle[2] ),
    .B(\inst$top.soc.spiflash.phy.enframer.cycle[1] ),
    .Y(_18729_));
 sky130_fd_sc_hd__inv_1 _40824_ (.A(_18729_),
    .Y(_18730_));
 sky130_fd_sc_hd__nor3_1 _40825_ (.A(_18730_),
    .B(_18701_),
    .C(_18643_),
    .Y(_18731_));
 sky130_fd_sc_hd__nand3_1 _40826_ (.A(_18713_),
    .B(_18281_),
    .C(_18731_),
    .Y(_18732_));
 sky130_fd_sc_hd__nand2_1 _40827_ (.A(net806),
    .B(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io2.o ),
    .Y(_18733_));
 sky130_fd_sc_hd__nand2_1 _40828_ (.A(_18732_),
    .B(_18733_),
    .Y(\inst$top.soc.spiflash.phy.io_streamer.buffer_io2.o ));
 sky130_fd_sc_hd__a21oi_1 _40830_ (.A1(_18732_),
    .A2(_18733_),
    .B1(net2946),
    .Y(_05282_));
 sky130_fd_sc_hd__nand2_1 _40831_ (.A(_18713_),
    .B(_18281_),
    .Y(_18735_));
 sky130_fd_sc_hd__nand2_1 _40832_ (.A(_18628_),
    .B(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io2.oe ),
    .Y(_18736_));
 sky130_fd_sc_hd__nand2_1 _40833_ (.A(_18735_),
    .B(_18736_),
    .Y(\inst$top.soc.spiflash.phy.io_streamer.buffer_io2.oe ));
 sky130_fd_sc_hd__a21oi_1 _40834_ (.A1(_18735_),
    .A2(_18736_),
    .B1(net2965),
    .Y(_05283_));
 sky130_fd_sc_hd__a211oi_1 _40835_ (.A1(_18650_),
    .A2(\inst$top.soc.spiflash.phy.enframer.cycle[0] ),
    .B1(_18719_),
    .C1(_18730_),
    .Y(_18737_));
 sky130_fd_sc_hd__nand3_1 _40836_ (.A(_18713_),
    .B(_18281_),
    .C(_18737_),
    .Y(_18738_));
 sky130_fd_sc_hd__nand2_1 _40837_ (.A(net806),
    .B(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io3.o ),
    .Y(_18739_));
 sky130_fd_sc_hd__nand2_1 _40838_ (.A(_18738_),
    .B(_18739_),
    .Y(\inst$top.soc.spiflash.phy.io_streamer.buffer_io3.o ));
 sky130_fd_sc_hd__a21oi_1 _40839_ (.A1(_18738_),
    .A2(_18739_),
    .B1(net2946),
    .Y(_05284_));
 sky130_fd_sc_hd__nand2_1 _40840_ (.A(net806),
    .B(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io3.oe ),
    .Y(_18740_));
 sky130_fd_sc_hd__nand2_1 _40841_ (.A(_18735_),
    .B(_18740_),
    .Y(\inst$top.soc.spiflash.phy.io_streamer.buffer_io3.oe ));
 sky130_fd_sc_hd__a21oi_1 _40842_ (.A1(_18735_),
    .A2(_18740_),
    .B1(net2965),
    .Y(_05285_));
 sky130_fd_sc_hd__nand2_1 _40843_ (.A(_18534_),
    .B(\inst$top.soc.spiflash.phy.io_streamer.i_en_0 ),
    .Y(_18741_));
 sky130_fd_sc_hd__o21ai_0 _40846_ (.A1(\inst$top.soc.spiflash.phy.io_streamer.buffer_io0.i_ff ),
    .A2(net827),
    .B1(net2047),
    .Y(_18744_));
 sky130_fd_sc_hd__a21oi_1 _40847_ (.A1(_18409_),
    .A2(net827),
    .B1(_18744_),
    .Y(_05286_));
 sky130_fd_sc_hd__nand2_1 _40848_ (.A(net827),
    .B(\inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io1 ),
    .Y(_18745_));
 sky130_fd_sc_hd__nand3_1 _40849_ (.A(_18534_),
    .B(\inst$top.soc.spiflash.phy.io_streamer.i_en_0 ),
    .C(\inst$top.soc.spiflash.phy.io_streamer.buffer_io1.i_ff ),
    .Y(_18746_));
 sky130_fd_sc_hd__a21oi_1 _40850_ (.A1(_18745_),
    .A2(_18746_),
    .B1(net2947),
    .Y(_05287_));
 sky130_fd_sc_hd__o21ai_0 _40851_ (.A1(\inst$top.soc.spiflash.phy.io_streamer.buffer_io2.i_ff ),
    .A2(_18741_),
    .B1(net2048),
    .Y(_18747_));
 sky130_fd_sc_hd__a21oi_1 _40852_ (.A1(_18421_),
    .A2(_18741_),
    .B1(_18747_),
    .Y(_05288_));
 sky130_fd_sc_hd__o21ai_0 _40853_ (.A1(\inst$top.soc.spiflash.phy.io_streamer.buffer_io3.i_ff ),
    .A2(net827),
    .B1(net2048),
    .Y(_18748_));
 sky130_fd_sc_hd__a21oi_1 _40854_ (.A1(_18431_),
    .A2(net827),
    .B1(_18748_),
    .Y(_05289_));
 sky130_fd_sc_hd__nand2_1 _40855_ (.A(net827),
    .B(\inst$top.soc.spiflash.phy.io_streamer.skid_1.meta[0] ),
    .Y(_18749_));
 sky130_fd_sc_hd__nand3_1 _40856_ (.A(_18534_),
    .B(\inst$top.soc.spiflash.phy.io_streamer.i_en_0 ),
    .C(\inst$top.soc.spiflash.phy.io_streamer.meta_0[0] ),
    .Y(_18750_));
 sky130_fd_sc_hd__a21oi_1 _40857_ (.A1(_18749_),
    .A2(_18750_),
    .B1(net2947),
    .Y(_05290_));
 sky130_fd_sc_hd__o21ai_0 _40858_ (.A1(\inst$top.soc.spiflash.phy.io_streamer.meta_0[1] ),
    .A2(net827),
    .B1(net2047),
    .Y(_18751_));
 sky130_fd_sc_hd__a21oi_1 _40859_ (.A1(_18225_),
    .A2(net827),
    .B1(_18751_),
    .Y(_05291_));
 sky130_fd_sc_hd__o21ai_0 _40860_ (.A1(\inst$top.soc.spiflash.phy.io_streamer.meta_0[2] ),
    .A2(net827),
    .B1(net2047),
    .Y(_18752_));
 sky130_fd_sc_hd__a21oi_1 _40861_ (.A1(_18219_),
    .A2(net827),
    .B1(_18752_),
    .Y(_05292_));
 sky130_fd_sc_hd__a211oi_1 _40862_ (.A1(\inst$top.soc.spiflash.phy.io_streamer.skid_at ),
    .A2(\inst$top.soc.spiflash.phy.io_streamer.i_en_0 ),
    .B1(net2947),
    .C1(_18244_),
    .Y(_05293_));
 sky130_fd_sc_hd__nor2_1 _40863_ (.A(net2951),
    .B(_09347_),
    .Y(_05294_));
 sky130_fd_sc_hd__nand2_1 _40865_ (.A(net547),
    .B(_02879_),
    .Y(_18754_));
 sky130_fd_sc_hd__o21ai_1 _40866_ (.A1(net1835),
    .A2(_02879_),
    .B1(_18754_),
    .Y(_18755_));
 sky130_fd_sc_hd__inv_1 _40867_ (.A(_02882_),
    .Y(_18756_));
 sky130_fd_sc_hd__nor2_1 _40868_ (.A(net1766),
    .B(_09353_),
    .Y(_18757_));
 sky130_fd_sc_hd__nor2_1 _40869_ (.A(net1637),
    .B(_18757_),
    .Y(_18758_));
 sky130_fd_sc_hd__inv_1 _40870_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.Config.enable._storage ),
    .Y(_18759_));
 sky130_fd_sc_hd__nor2_1 _40871_ (.A(net2995),
    .B(_18759_),
    .Y(_18760_));
 sky130_fd_sc_hd__o21ai_0 _40873_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.bitno[0] ),
    .A2(_18758_),
    .B1(net1856),
    .Y(_18762_));
 sky130_fd_sc_hd__a31oi_1 _40874_ (.A1(net1835),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.bitno[0] ),
    .A3(_18758_),
    .B1(_18762_),
    .Y(_05295_));
 sky130_fd_sc_hd__inv_1 _40875_ (.A(_18758_),
    .Y(_18763_));
 sky130_fd_sc_hd__nand2_1 _40876_ (.A(_18763_),
    .B(\inst$top.soc.uart_0._phy.rx.lower.bitno[1] ),
    .Y(_18764_));
 sky130_fd_sc_hd__nor2_1 _40878_ (.A(_02717_),
    .B(_18756_),
    .Y(_18766_));
 sky130_fd_sc_hd__nand2_1 _40879_ (.A(_18758_),
    .B(_18766_),
    .Y(_18767_));
 sky130_fd_sc_hd__inv_1 _40880_ (.A(net1856),
    .Y(_18768_));
 sky130_fd_sc_hd__a21oi_1 _40882_ (.A1(_18764_),
    .A2(_18767_),
    .B1(net1765),
    .Y(_05296_));
 sky130_fd_sc_hd__inv_1 _40883_ (.A(_02716_),
    .Y(_18770_));
 sky130_fd_sc_hd__nor2_1 _40884_ (.A(_18770_),
    .B(_18763_),
    .Y(_18771_));
 sky130_fd_sc_hd__nor2_1 _40886_ (.A(net1835),
    .B(net1637),
    .Y(_18773_));
 sky130_fd_sc_hd__clkinv_1 _40887_ (.A(_18773_),
    .Y(_18774_));
 sky130_fd_sc_hd__o21ai_0 _40888_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.bitno[2] ),
    .A2(_18771_),
    .B1(_18774_),
    .Y(_18775_));
 sky130_fd_sc_hd__a211oi_1 _40889_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.bitno[2] ),
    .A2(_18771_),
    .B1(net1765),
    .C1(_18775_),
    .Y(_05297_));
 sky130_fd_sc_hd__nor2_1 _40890_ (.A(\inst$top.soc.uart_0._phy.rx.lower.bitno[2] ),
    .B(\inst$top.soc.uart_0._phy.rx.lower.bitno[1] ),
    .Y(_18776_));
 sky130_fd_sc_hd__nand2_1 _40891_ (.A(_18776_),
    .B(_02714_),
    .Y(_18777_));
 sky130_fd_sc_hd__or3_1 _40892_ (.A(\inst$top.soc.uart_0._phy.rx.lower.bitno[3] ),
    .B(_18777_),
    .C(_18763_),
    .X(_18778_));
 sky130_fd_sc_hd__o21ai_0 _40893_ (.A1(_18777_),
    .A2(_18763_),
    .B1(\inst$top.soc.uart_0._phy.rx.lower.bitno[3] ),
    .Y(_18779_));
 sky130_fd_sc_hd__a31oi_1 _40895_ (.A1(_18778_),
    .A2(_18774_),
    .A3(_18779_),
    .B1(net1765),
    .Y(_05298_));
 sky130_fd_sc_hd__inv_1 _40896_ (.A(\inst$top.soc.uart_0._phy.rx.lower.shreg[1] ),
    .Y(_18781_));
 sky130_fd_sc_hd__o21ai_0 _40899_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.data[0] ),
    .A2(net1837),
    .B1(net1855),
    .Y(_18784_));
 sky130_fd_sc_hd__a21oi_1 _40900_ (.A1(_18781_),
    .A2(net1837),
    .B1(_18784_),
    .Y(_05299_));
 sky130_fd_sc_hd__inv_1 _40901_ (.A(net1836),
    .Y(_18785_));
 sky130_fd_sc_hd__nand2_1 _40902_ (.A(_18785_),
    .B(\inst$top.soc.uart_0._phy.rx.lower.data[1] ),
    .Y(_18786_));
 sky130_fd_sc_hd__nand2_1 _40903_ (.A(net1837),
    .B(\inst$top.soc.uart_0._phy.rx.lower.shreg[2] ),
    .Y(_18787_));
 sky130_fd_sc_hd__a21oi_1 _40904_ (.A1(_18786_),
    .A2(_18787_),
    .B1(net1764),
    .Y(_05300_));
 sky130_fd_sc_hd__inv_1 _40905_ (.A(\inst$top.soc.uart_0._phy.rx.lower.shreg[3] ),
    .Y(_18788_));
 sky130_fd_sc_hd__o21ai_0 _40906_ (.A1(net1836),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.data[2] ),
    .B1(net1854),
    .Y(_18789_));
 sky130_fd_sc_hd__a21oi_1 _40907_ (.A1(net1836),
    .A2(_18788_),
    .B1(_18789_),
    .Y(_05301_));
 sky130_fd_sc_hd__inv_1 _40908_ (.A(\inst$top.soc.uart_0._phy.rx.lower.shreg[4] ),
    .Y(_18790_));
 sky130_fd_sc_hd__o21ai_0 _40909_ (.A1(net1836),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.data[3] ),
    .B1(net1856),
    .Y(_18791_));
 sky130_fd_sc_hd__a21oi_1 _40910_ (.A1(net1836),
    .A2(_18790_),
    .B1(_18791_),
    .Y(_05302_));
 sky130_fd_sc_hd__inv_1 _40911_ (.A(\inst$top.soc.uart_0._phy.rx.lower.shreg[5] ),
    .Y(_18792_));
 sky130_fd_sc_hd__o21ai_0 _40912_ (.A1(net1836),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.data[4] ),
    .B1(net1854),
    .Y(_18793_));
 sky130_fd_sc_hd__a21oi_1 _40913_ (.A1(net1836),
    .A2(_18792_),
    .B1(_18793_),
    .Y(_05303_));
 sky130_fd_sc_hd__inv_1 _40914_ (.A(\inst$top.soc.uart_0._phy.rx.lower.shreg[6] ),
    .Y(_18794_));
 sky130_fd_sc_hd__o21ai_0 _40915_ (.A1(net1837),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.data[5] ),
    .B1(net1855),
    .Y(_18795_));
 sky130_fd_sc_hd__a21oi_1 _40916_ (.A1(net1837),
    .A2(_18794_),
    .B1(_18795_),
    .Y(_05304_));
 sky130_fd_sc_hd__nand2_1 _40917_ (.A(_18785_),
    .B(\inst$top.soc.uart_0._phy.rx.lower.data[6] ),
    .Y(_18796_));
 sky130_fd_sc_hd__nand2_1 _40918_ (.A(net1836),
    .B(\inst$top.soc.uart_0._phy.rx.lower.shreg[7] ),
    .Y(_18797_));
 sky130_fd_sc_hd__a21oi_1 _40919_ (.A1(_18796_),
    .A2(_18797_),
    .B1(net1764),
    .Y(_05305_));
 sky130_fd_sc_hd__inv_1 _40920_ (.A(\inst$top.soc.uart_0._phy.rx.lower.shreg[8] ),
    .Y(_18798_));
 sky130_fd_sc_hd__o21ai_0 _40921_ (.A1(net1836),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.data[7] ),
    .B1(net1854),
    .Y(_18799_));
 sky130_fd_sc_hd__a21oi_1 _40922_ (.A1(net1836),
    .A2(_18798_),
    .B1(_18799_),
    .Y(_05306_));
 sky130_fd_sc_hd__inv_1 _40923_ (.A(\inst$top.soc.uart_0._phy.rx.lower.shreg.start ),
    .Y(_18800_));
 sky130_fd_sc_hd__o21ai_0 _40924_ (.A1(\inst$top.soc.uart_0._phy.rx.err.frame ),
    .A2(net1837),
    .B1(net1855),
    .Y(_18801_));
 sky130_fd_sc_hd__a31oi_1 _40925_ (.A1(_18800_),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.shreg.stop ),
    .A3(net1837),
    .B1(_18801_),
    .Y(_05307_));
 sky130_fd_sc_hd__nor2_1 _40926_ (.A(\inst$top.soc.uart_0._phy.rx.lower.bitno[3] ),
    .B(\inst$top.soc.uart_0._phy.rx.lower.bitno[2] ),
    .Y(_18802_));
 sky130_fd_sc_hd__a21oi_1 _40927_ (.A1(_18802_),
    .A2(_02718_),
    .B1(net1766),
    .Y(_18803_));
 sky130_fd_sc_hd__nor3b_1 _40928_ (.A(_02883_),
    .B(_18803_),
    .C_N(_18754_),
    .Y(_18804_));
 sky130_fd_sc_hd__o21ai_0 _40929_ (.A1(_18756_),
    .A2(_09353_),
    .B1(_18804_),
    .Y(_18805_));
 sky130_fd_sc_hd__or2_2 _40930_ (.A(_02880_),
    .B(_18805_),
    .X(_18806_));
 sky130_fd_sc_hd__nand2_1 _40931_ (.A(_18805_),
    .B(\inst$top.soc.uart_0._phy.rx.lower.fsm_state[0] ),
    .Y(_18807_));
 sky130_fd_sc_hd__a21oi_1 _40932_ (.A1(_18806_),
    .A2(_18807_),
    .B1(net1765),
    .Y(_05308_));
 sky130_fd_sc_hd__nor2_1 _40934_ (.A(_18756_),
    .B(_07483_),
    .Y(_18809_));
 sky130_fd_sc_hd__a22oi_1 _40936_ (.A1(net1226),
    .A2(_18804_),
    .B1(_18805_),
    .B2(\inst$top.soc.uart_0._phy.rx.lower.fsm_state[1] ),
    .Y(_18811_));
 sky130_fd_sc_hd__nor2_1 _40937_ (.A(net1764),
    .B(_18811_),
    .Y(_05309_));
 sky130_fd_sc_hd__nor2_1 _40938_ (.A(_18785_),
    .B(net1763),
    .Y(_05310_));
 sky130_fd_sc_hd__o21ai_0 _40939_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.shreg.start ),
    .A2(_18809_),
    .B1(net1855),
    .Y(_18812_));
 sky130_fd_sc_hd__a21oi_1 _40940_ (.A1(_18781_),
    .A2(_18809_),
    .B1(_18812_),
    .Y(_05311_));
 sky130_fd_sc_hd__inv_2 _40941_ (.A(net1226),
    .Y(_18813_));
 sky130_fd_sc_hd__o21ai_0 _40942_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.shreg[2] ),
    .A2(_18813_),
    .B1(net1855),
    .Y(_18814_));
 sky130_fd_sc_hd__a21oi_1 _40943_ (.A1(_18781_),
    .A2(_18813_),
    .B1(_18814_),
    .Y(_05312_));
 sky130_fd_sc_hd__o21ai_0 _40944_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.shreg[2] ),
    .A2(_18809_),
    .B1(net1854),
    .Y(_18815_));
 sky130_fd_sc_hd__a21oi_1 _40945_ (.A1(_18788_),
    .A2(net1226),
    .B1(_18815_),
    .Y(_05313_));
 sky130_fd_sc_hd__o21ai_0 _40946_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.shreg[3] ),
    .A2(net1226),
    .B1(net1854),
    .Y(_18816_));
 sky130_fd_sc_hd__a21oi_1 _40947_ (.A1(_18790_),
    .A2(net1226),
    .B1(_18816_),
    .Y(_05314_));
 sky130_fd_sc_hd__o21ai_0 _40948_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.shreg[4] ),
    .A2(net1226),
    .B1(net1854),
    .Y(_18817_));
 sky130_fd_sc_hd__a21oi_1 _40949_ (.A1(_18792_),
    .A2(net1226),
    .B1(_18817_),
    .Y(_05315_));
 sky130_fd_sc_hd__o21ai_0 _40950_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.shreg[6] ),
    .A2(_18813_),
    .B1(net1854),
    .Y(_18818_));
 sky130_fd_sc_hd__a21oi_1 _40951_ (.A1(_18792_),
    .A2(_18813_),
    .B1(_18818_),
    .Y(_05316_));
 sky130_fd_sc_hd__o21ai_0 _40952_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.shreg[7] ),
    .A2(_18813_),
    .B1(net1854),
    .Y(_18819_));
 sky130_fd_sc_hd__a21oi_1 _40953_ (.A1(_18794_),
    .A2(_18813_),
    .B1(_18819_),
    .Y(_05317_));
 sky130_fd_sc_hd__o21ai_0 _40954_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.shreg[7] ),
    .A2(net1226),
    .B1(net1854),
    .Y(_18820_));
 sky130_fd_sc_hd__a21oi_1 _40955_ (.A1(_18798_),
    .A2(net1226),
    .B1(_18820_),
    .Y(_05318_));
 sky130_fd_sc_hd__o21ai_0 _40956_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.shreg.stop ),
    .A2(_18813_),
    .B1(net1854),
    .Y(_18821_));
 sky130_fd_sc_hd__a21oi_1 _40957_ (.A1(_18798_),
    .A2(_18813_),
    .B1(_18821_),
    .Y(_05319_));
 sky130_fd_sc_hd__nor2_1 _40958_ (.A(net547),
    .B(_18813_),
    .Y(_18822_));
 sky130_fd_sc_hd__o21ai_0 _40959_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.shreg.stop ),
    .A2(net1226),
    .B1(net1855),
    .Y(_18823_));
 sky130_fd_sc_hd__nor2_1 _40960_ (.A(_18822_),
    .B(_18823_),
    .Y(_05320_));
 sky130_fd_sc_hd__inv_1 _40961_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[1] ),
    .Y(_18824_));
 sky130_fd_sc_hd__nand2_1 _40962_ (.A(_18754_),
    .B(net1835),
    .Y(_18825_));
 sky130_fd_sc_hd__a21oi_1 _40964_ (.A1(net1636),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.timer[0] ),
    .B1(net1762),
    .Y(_18827_));
 sky130_fd_sc_hd__o221ai_1 _40965_ (.A1(_18824_),
    .A2(_18774_),
    .B1(_18825_),
    .B2(_07485_),
    .C1(_18827_),
    .Y(_05321_));
 sky130_fd_sc_hd__inv_1 _40966_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[2] ),
    .Y(_18828_));
 sky130_fd_sc_hd__o21bai_1 _40967_ (.A1(_18828_),
    .A2(net1667),
    .B1_N(\inst$top.soc.uart_0._phy.rx.lower.timer[2] ),
    .Y(_18829_));
 sky130_fd_sc_hd__inv_1 _40968_ (.A(_18829_),
    .Y(_18830_));
 sky130_fd_sc_hd__nand2_1 _40969_ (.A(_18830_),
    .B(_02721_),
    .Y(_18831_));
 sky130_fd_sc_hd__inv_1 _40970_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[4] ),
    .Y(_18832_));
 sky130_fd_sc_hd__o21bai_1 _40971_ (.A1(_18832_),
    .A2(net1667),
    .B1_N(\inst$top.soc.uart_0._phy.rx.lower.timer[4] ),
    .Y(_18833_));
 sky130_fd_sc_hd__inv_1 _40972_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[3] ),
    .Y(_18834_));
 sky130_fd_sc_hd__o21bai_1 _40973_ (.A1(_18834_),
    .A2(net1667),
    .B1_N(\inst$top.soc.uart_0._phy.rx.lower.timer[3] ),
    .Y(_18835_));
 sky130_fd_sc_hd__nor2_1 _40974_ (.A(_18833_),
    .B(_18835_),
    .Y(_18836_));
 sky130_fd_sc_hd__inv_1 _40975_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[5] ),
    .Y(_18837_));
 sky130_fd_sc_hd__o21bai_1 _40976_ (.A1(_18837_),
    .A2(net1667),
    .B1_N(\inst$top.soc.uart_0._phy.rx.lower.timer[5] ),
    .Y(_18838_));
 sky130_fd_sc_hd__inv_1 _40977_ (.A(_18838_),
    .Y(_18839_));
 sky130_fd_sc_hd__nand2_1 _40978_ (.A(_18836_),
    .B(_18839_),
    .Y(_18840_));
 sky130_fd_sc_hd__nor2_1 _40979_ (.A(_18831_),
    .B(_18840_),
    .Y(_18841_));
 sky130_fd_sc_hd__a21oi_1 _40980_ (.A1(_09353_),
    .A2(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[6] ),
    .B1(\inst$top.soc.uart_0._phy.rx.lower.timer[6] ),
    .Y(_18842_));
 sky130_fd_sc_hd__inv_1 _40981_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[7] ),
    .Y(_18843_));
 sky130_fd_sc_hd__o21bai_1 _40982_ (.A1(_18843_),
    .A2(net1667),
    .B1_N(\inst$top.soc.uart_0._phy.rx.lower.timer[7] ),
    .Y(_18844_));
 sky130_fd_sc_hd__inv_1 _40983_ (.A(_18844_),
    .Y(_18845_));
 sky130_fd_sc_hd__nand2_1 _40984_ (.A(_18842_),
    .B(_18845_),
    .Y(_18846_));
 sky130_fd_sc_hd__a21oi_1 _40985_ (.A1(_09353_),
    .A2(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[9] ),
    .B1(\inst$top.soc.uart_0._phy.rx.lower.timer[9] ),
    .Y(_18847_));
 sky130_fd_sc_hd__a21oi_1 _40986_ (.A1(_09353_),
    .A2(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[8] ),
    .B1(\inst$top.soc.uart_0._phy.rx.lower.timer[8] ),
    .Y(_18848_));
 sky130_fd_sc_hd__nand2_1 _40987_ (.A(_18847_),
    .B(_18848_),
    .Y(_18849_));
 sky130_fd_sc_hd__nor2_1 _40988_ (.A(_18846_),
    .B(_18849_),
    .Y(_18850_));
 sky130_fd_sc_hd__nand2_1 _40989_ (.A(_18841_),
    .B(_18850_),
    .Y(_18851_));
 sky130_fd_sc_hd__inv_1 _40990_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[10] ),
    .Y(_18852_));
 sky130_fd_sc_hd__o21ai_0 _40991_ (.A1(_18852_),
    .A2(_07483_),
    .B1(_07471_),
    .Y(_18853_));
 sky130_fd_sc_hd__inv_1 _40992_ (.A(_18853_),
    .Y(_18854_));
 sky130_fd_sc_hd__nand2_1 _40993_ (.A(_18851_),
    .B(_18854_),
    .Y(_18855_));
 sky130_fd_sc_hd__inv_1 _40994_ (.A(_18825_),
    .Y(_18856_));
 sky130_fd_sc_hd__nand3_1 _40995_ (.A(_18841_),
    .B(_18850_),
    .C(_18853_),
    .Y(_18857_));
 sky130_fd_sc_hd__nand3_1 _40996_ (.A(_18855_),
    .B(net1224),
    .C(_18857_),
    .Y(_18858_));
 sky130_fd_sc_hd__nand2_1 _40998_ (.A(net1637),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[10] ),
    .Y(_18860_));
 sky130_fd_sc_hd__nand2_1 _40999_ (.A(_18773_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[11] ),
    .Y(_18861_));
 sky130_fd_sc_hd__a31oi_1 _41000_ (.A1(_18858_),
    .A2(_18860_),
    .A3(_18861_),
    .B1(net1764),
    .Y(_05322_));
 sky130_fd_sc_hd__nand4_1 _41001_ (.A(_18842_),
    .B(_18848_),
    .C(_18845_),
    .D(_18839_),
    .Y(_18862_));
 sky130_fd_sc_hd__inv_1 _41002_ (.A(_18836_),
    .Y(_18863_));
 sky130_fd_sc_hd__nand3_1 _41003_ (.A(_02719_),
    .B(_18830_),
    .C(_02720_),
    .Y(_18864_));
 sky130_fd_sc_hd__nor2_1 _41004_ (.A(_18863_),
    .B(_18864_),
    .Y(_18865_));
 sky130_fd_sc_hd__inv_1 _41005_ (.A(_18865_),
    .Y(_18866_));
 sky130_fd_sc_hd__nor2_1 _41006_ (.A(_18862_),
    .B(_18866_),
    .Y(_18867_));
 sky130_fd_sc_hd__nand3_1 _41007_ (.A(_18867_),
    .B(_18847_),
    .C(_18854_),
    .Y(_18868_));
 sky130_fd_sc_hd__inv_1 _41008_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[11] ),
    .Y(_18869_));
 sky130_fd_sc_hd__o21ai_0 _41009_ (.A1(_18869_),
    .A2(net1668),
    .B1(_07475_),
    .Y(_18870_));
 sky130_fd_sc_hd__nand2_1 _41010_ (.A(_18868_),
    .B(_18870_),
    .Y(_18871_));
 sky130_fd_sc_hd__nor2_1 _41011_ (.A(_18853_),
    .B(_18870_),
    .Y(_18872_));
 sky130_fd_sc_hd__nand3_1 _41012_ (.A(_18867_),
    .B(_18847_),
    .C(_18872_),
    .Y(_18873_));
 sky130_fd_sc_hd__nand2_1 _41013_ (.A(_18871_),
    .B(_18873_),
    .Y(_18874_));
 sky130_fd_sc_hd__nand2_1 _41015_ (.A(_18874_),
    .B(net1225),
    .Y(_18876_));
 sky130_fd_sc_hd__nand2_1 _41016_ (.A(net1637),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[11] ),
    .Y(_18877_));
 sky130_fd_sc_hd__nand2_1 _41017_ (.A(_18773_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[12] ),
    .Y(_18878_));
 sky130_fd_sc_hd__a31oi_1 _41018_ (.A1(_18876_),
    .A2(_18877_),
    .A3(_18878_),
    .B1(net1764),
    .Y(_05323_));
 sky130_fd_sc_hd__inv_1 _41019_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[12] ),
    .Y(_18879_));
 sky130_fd_sc_hd__inv_1 _41020_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[12] ),
    .Y(_18880_));
 sky130_fd_sc_hd__o21ai_0 _41021_ (.A1(_18879_),
    .A2(net1668),
    .B1(_18880_),
    .Y(_18881_));
 sky130_fd_sc_hd__nor2_1 _41022_ (.A(_18838_),
    .B(_18833_),
    .Y(_18882_));
 sky130_fd_sc_hd__nand3_1 _41023_ (.A(_18882_),
    .B(_18842_),
    .C(_18845_),
    .Y(_18883_));
 sky130_fd_sc_hd__nand3_1 _41024_ (.A(_18872_),
    .B(_18847_),
    .C(_18848_),
    .Y(_18884_));
 sky130_fd_sc_hd__nor2_1 _41025_ (.A(_18883_),
    .B(_18884_),
    .Y(_18885_));
 sky130_fd_sc_hd__nor2_1 _41026_ (.A(_18835_),
    .B(_18829_),
    .Y(_18886_));
 sky130_fd_sc_hd__nand2_1 _41027_ (.A(_18886_),
    .B(_02721_),
    .Y(_18887_));
 sky130_fd_sc_hd__inv_1 _41028_ (.A(_18887_),
    .Y(_18888_));
 sky130_fd_sc_hd__nand2_1 _41029_ (.A(_18885_),
    .B(_18888_),
    .Y(_18889_));
 sky130_fd_sc_hd__xnor2_1 _41030_ (.A(_18881_),
    .B(_18889_),
    .Y(_18890_));
 sky130_fd_sc_hd__nand2_1 _41031_ (.A(_18890_),
    .B(net1225),
    .Y(_18891_));
 sky130_fd_sc_hd__nand2_1 _41032_ (.A(_18755_),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[12] ),
    .Y(_18892_));
 sky130_fd_sc_hd__nand2_1 _41033_ (.A(_18773_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[13] ),
    .Y(_18893_));
 sky130_fd_sc_hd__a31oi_1 _41034_ (.A1(_18891_),
    .A2(_18892_),
    .A3(_18893_),
    .B1(net1764),
    .Y(_05324_));
 sky130_fd_sc_hd__inv_1 _41035_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[13] ),
    .Y(_18894_));
 sky130_fd_sc_hd__inv_1 _41036_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[13] ),
    .Y(_18895_));
 sky130_fd_sc_hd__o21ai_0 _41037_ (.A1(_18894_),
    .A2(net1668),
    .B1(_18895_),
    .Y(_18896_));
 sky130_fd_sc_hd__nor2_1 _41038_ (.A(_18870_),
    .B(_18881_),
    .Y(_18897_));
 sky130_fd_sc_hd__nand3_1 _41039_ (.A(_18897_),
    .B(_18847_),
    .C(_18854_),
    .Y(_18898_));
 sky130_fd_sc_hd__inv_1 _41040_ (.A(_18862_),
    .Y(_18899_));
 sky130_fd_sc_hd__nand2_1 _41041_ (.A(_18899_),
    .B(_18865_),
    .Y(_18900_));
 sky130_fd_sc_hd__nor2_1 _41042_ (.A(_18898_),
    .B(_18900_),
    .Y(_18901_));
 sky130_fd_sc_hd__xor2_1 _41043_ (.A(_18896_),
    .B(_18901_),
    .X(_18902_));
 sky130_fd_sc_hd__nand2_1 _41044_ (.A(_18902_),
    .B(net1225),
    .Y(_18903_));
 sky130_fd_sc_hd__nand2_1 _41045_ (.A(net1637),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[13] ),
    .Y(_18904_));
 sky130_fd_sc_hd__nand2_1 _41046_ (.A(_18773_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[14] ),
    .Y(_18905_));
 sky130_fd_sc_hd__a31oi_1 _41047_ (.A1(_18903_),
    .A2(_18904_),
    .A3(_18905_),
    .B1(net1764),
    .Y(_05325_));
 sky130_fd_sc_hd__inv_1 _41048_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[14] ),
    .Y(_18906_));
 sky130_fd_sc_hd__o21bai_1 _41049_ (.A1(_18906_),
    .A2(net1668),
    .B1_N(\inst$top.soc.uart_0._phy.rx.lower.timer[14] ),
    .Y(_18907_));
 sky130_fd_sc_hd__nor2_1 _41050_ (.A(_18881_),
    .B(_18896_),
    .Y(_18908_));
 sky130_fd_sc_hd__nand2_1 _41051_ (.A(_18872_),
    .B(_18908_),
    .Y(_18909_));
 sky130_fd_sc_hd__nor2_1 _41052_ (.A(_18909_),
    .B(_18851_),
    .Y(_18910_));
 sky130_fd_sc_hd__xor2_1 _41053_ (.A(_18907_),
    .B(_18910_),
    .X(_18911_));
 sky130_fd_sc_hd__nand2_1 _41054_ (.A(_18911_),
    .B(net1225),
    .Y(_18912_));
 sky130_fd_sc_hd__nand2_1 _41055_ (.A(net1637),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[14] ),
    .Y(_18913_));
 sky130_fd_sc_hd__nand2_1 _41056_ (.A(_18773_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[15] ),
    .Y(_18914_));
 sky130_fd_sc_hd__a31oi_1 _41057_ (.A1(_18912_),
    .A2(_18913_),
    .A3(_18914_),
    .B1(net1764),
    .Y(_05326_));
 sky130_fd_sc_hd__nor2_1 _41058_ (.A(_18907_),
    .B(_18896_),
    .Y(_18915_));
 sky130_fd_sc_hd__nand2_1 _41059_ (.A(_18897_),
    .B(_18915_),
    .Y(_18916_));
 sky130_fd_sc_hd__nor2_1 _41060_ (.A(_18916_),
    .B(_18868_),
    .Y(_18917_));
 sky130_fd_sc_hd__inv_1 _41061_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[15] ),
    .Y(_18918_));
 sky130_fd_sc_hd__inv_1 _41062_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[15] ),
    .Y(_18919_));
 sky130_fd_sc_hd__o21ai_0 _41063_ (.A1(_18918_),
    .A2(net1668),
    .B1(_18919_),
    .Y(_18920_));
 sky130_fd_sc_hd__nand2_1 _41064_ (.A(_18917_),
    .B(_18920_),
    .Y(_18921_));
 sky130_fd_sc_hd__inv_1 _41065_ (.A(_18896_),
    .Y(_18922_));
 sky130_fd_sc_hd__inv_1 _41066_ (.A(_18907_),
    .Y(_18923_));
 sky130_fd_sc_hd__nand3_1 _41067_ (.A(_18901_),
    .B(_18922_),
    .C(_18923_),
    .Y(_18924_));
 sky130_fd_sc_hd__inv_1 _41068_ (.A(_18920_),
    .Y(_18925_));
 sky130_fd_sc_hd__nand2_1 _41069_ (.A(_18924_),
    .B(_18925_),
    .Y(_18926_));
 sky130_fd_sc_hd__inv_2 _41070_ (.A(net1635),
    .Y(_18927_));
 sky130_fd_sc_hd__inv_1 _41071_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[16] ),
    .Y(_18928_));
 sky130_fd_sc_hd__o22ai_1 _41072_ (.A1(_18919_),
    .A2(_18927_),
    .B1(_18928_),
    .B2(_18774_),
    .Y(_18929_));
 sky130_fd_sc_hd__a31oi_1 _41073_ (.A1(_18921_),
    .A2(_18926_),
    .A3(net1225),
    .B1(_18929_),
    .Y(_18930_));
 sky130_fd_sc_hd__nor2_1 _41074_ (.A(net1763),
    .B(_18930_),
    .Y(_05327_));
 sky130_fd_sc_hd__o21ai_0 _41075_ (.A1(_18928_),
    .A2(net1668),
    .B1(_07476_),
    .Y(_18931_));
 sky130_fd_sc_hd__nand3_1 _41076_ (.A(_18908_),
    .B(_18923_),
    .C(_18925_),
    .Y(_18932_));
 sky130_fd_sc_hd__or2_2 _41077_ (.A(_18887_),
    .B(_18883_),
    .X(_18933_));
 sky130_fd_sc_hd__nor3_1 _41078_ (.A(_18884_),
    .B(_18932_),
    .C(_18933_),
    .Y(_18934_));
 sky130_fd_sc_hd__xor2_1 _41079_ (.A(_18931_),
    .B(_18934_),
    .X(_18935_));
 sky130_fd_sc_hd__inv_1 _41080_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[17] ),
    .Y(_18936_));
 sky130_fd_sc_hd__o22ai_1 _41081_ (.A1(_07476_),
    .A2(_18927_),
    .B1(_18936_),
    .B2(_18774_),
    .Y(_18937_));
 sky130_fd_sc_hd__a21oi_1 _41082_ (.A1(_18935_),
    .A2(net1224),
    .B1(_18937_),
    .Y(_18938_));
 sky130_fd_sc_hd__nor2_1 _41083_ (.A(net1763),
    .B(_18938_),
    .Y(_05328_));
 sky130_fd_sc_hd__inv_1 _41084_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[17] ),
    .Y(_18939_));
 sky130_fd_sc_hd__o21ai_0 _41085_ (.A1(_18936_),
    .A2(net1667),
    .B1(_18939_),
    .Y(_18940_));
 sky130_fd_sc_hd__nor2_1 _41086_ (.A(_18920_),
    .B(_18931_),
    .Y(_18941_));
 sky130_fd_sc_hd__nand2_1 _41087_ (.A(_18941_),
    .B(_18915_),
    .Y(_18942_));
 sky130_fd_sc_hd__nor3_1 _41088_ (.A(_18898_),
    .B(_18942_),
    .C(_18900_),
    .Y(_18943_));
 sky130_fd_sc_hd__xor2_1 _41089_ (.A(_18940_),
    .B(_18943_),
    .X(_18944_));
 sky130_fd_sc_hd__nand2_1 _41090_ (.A(_18944_),
    .B(net1224),
    .Y(_18945_));
 sky130_fd_sc_hd__inv_1 _41091_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[18] ),
    .Y(_18946_));
 sky130_fd_sc_hd__o22ai_1 _41092_ (.A1(_18939_),
    .A2(_18927_),
    .B1(_18946_),
    .B2(_18774_),
    .Y(_18947_));
 sky130_fd_sc_hd__inv_1 _41093_ (.A(_18947_),
    .Y(_18948_));
 sky130_fd_sc_hd__a21oi_1 _41094_ (.A1(_18945_),
    .A2(_18948_),
    .B1(net1763),
    .Y(_05329_));
 sky130_fd_sc_hd__inv_1 _41095_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[18] ),
    .Y(_18949_));
 sky130_fd_sc_hd__o21ai_0 _41096_ (.A1(_18946_),
    .A2(net1667),
    .B1(_18949_),
    .Y(_18950_));
 sky130_fd_sc_hd__nor4_1 _41097_ (.A(_18907_),
    .B(_18920_),
    .C(_18931_),
    .D(_18940_),
    .Y(_18951_));
 sky130_fd_sc_hd__nand2_1 _41098_ (.A(_18910_),
    .B(_18951_),
    .Y(_18952_));
 sky130_fd_sc_hd__xnor2_1 _41099_ (.A(_18950_),
    .B(_18952_),
    .Y(_18953_));
 sky130_fd_sc_hd__nand2_1 _41100_ (.A(_18953_),
    .B(net1224),
    .Y(_18954_));
 sky130_fd_sc_hd__nand2_1 _41101_ (.A(net1636),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[18] ),
    .Y(_18955_));
 sky130_fd_sc_hd__nand2_1 _41102_ (.A(_18773_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[19] ),
    .Y(_18956_));
 sky130_fd_sc_hd__a31oi_1 _41103_ (.A1(_18954_),
    .A2(_18955_),
    .A3(_18956_),
    .B1(net1763),
    .Y(_05330_));
 sky130_fd_sc_hd__nor2_1 _41104_ (.A(_18940_),
    .B(_18950_),
    .Y(_18957_));
 sky130_fd_sc_hd__nand2_1 _41105_ (.A(_18941_),
    .B(_18957_),
    .Y(_18958_));
 sky130_fd_sc_hd__inv_1 _41106_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[19] ),
    .Y(_18959_));
 sky130_fd_sc_hd__o21ai_0 _41107_ (.A1(_18959_),
    .A2(net1668),
    .B1(_07477_),
    .Y(_18960_));
 sky130_fd_sc_hd__o21bai_1 _41108_ (.A1(_18958_),
    .A2(_18924_),
    .B1_N(_18960_),
    .Y(_18961_));
 sky130_fd_sc_hd__nor2_1 _41109_ (.A(_18958_),
    .B(_18924_),
    .Y(_18962_));
 sky130_fd_sc_hd__nand2_1 _41110_ (.A(_18962_),
    .B(_18960_),
    .Y(_18963_));
 sky130_fd_sc_hd__nand3_1 _41111_ (.A(_18961_),
    .B(_18963_),
    .C(net1224),
    .Y(_18964_));
 sky130_fd_sc_hd__inv_1 _41112_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[20] ),
    .Y(_18965_));
 sky130_fd_sc_hd__o22ai_1 _41113_ (.A1(_07477_),
    .A2(_18927_),
    .B1(_18965_),
    .B2(_18774_),
    .Y(_18966_));
 sky130_fd_sc_hd__inv_1 _41114_ (.A(_18966_),
    .Y(_18967_));
 sky130_fd_sc_hd__a21oi_2 _41115_ (.A1(_18964_),
    .A2(_18967_),
    .B1(net1763),
    .Y(_05331_));
 sky130_fd_sc_hd__nand2_1 _41116_ (.A(_18773_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[2] ),
    .Y(_18968_));
 sky130_fd_sc_hd__or2_2 _41117_ (.A(_02722_),
    .B(_18825_),
    .X(_18969_));
 sky130_fd_sc_hd__nand2_1 _41118_ (.A(net1635),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[1] ),
    .Y(_18970_));
 sky130_fd_sc_hd__a31oi_1 _41119_ (.A1(_18968_),
    .A2(_18969_),
    .A3(_18970_),
    .B1(net1762),
    .Y(_05332_));
 sky130_fd_sc_hd__o21ai_0 _41120_ (.A1(_18965_),
    .A2(net1668),
    .B1(_07467_),
    .Y(_18971_));
 sky130_fd_sc_hd__nor2_1 _41121_ (.A(_18931_),
    .B(_18940_),
    .Y(_18972_));
 sky130_fd_sc_hd__nor2_1 _41122_ (.A(_18950_),
    .B(_18960_),
    .Y(_18973_));
 sky130_fd_sc_hd__nand2_1 _41123_ (.A(_18972_),
    .B(_18973_),
    .Y(_18974_));
 sky130_fd_sc_hd__nor2_1 _41124_ (.A(_18974_),
    .B(_18932_),
    .Y(_18975_));
 sky130_fd_sc_hd__nand3_1 _41125_ (.A(_18885_),
    .B(_18975_),
    .C(_18888_),
    .Y(_18976_));
 sky130_fd_sc_hd__xnor2_1 _41126_ (.A(_18971_),
    .B(_18976_),
    .Y(_18977_));
 sky130_fd_sc_hd__nand2_1 _41127_ (.A(_18977_),
    .B(net1224),
    .Y(_18978_));
 sky130_fd_sc_hd__nand2_1 _41128_ (.A(net1635),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[20] ),
    .Y(_18979_));
 sky130_fd_sc_hd__nand2_1 _41129_ (.A(_18773_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[21] ),
    .Y(_18980_));
 sky130_fd_sc_hd__a31oi_1 _41130_ (.A1(_18978_),
    .A2(_18979_),
    .A3(_18980_),
    .B1(net1762),
    .Y(_05333_));
 sky130_fd_sc_hd__inv_1 _41131_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[21] ),
    .Y(_18981_));
 sky130_fd_sc_hd__o21ai_0 _41132_ (.A1(_18981_),
    .A2(net1667),
    .B1(_07466_),
    .Y(_18982_));
 sky130_fd_sc_hd__nor3_1 _41133_ (.A(_18960_),
    .B(_18971_),
    .C(_18958_),
    .Y(_18983_));
 sky130_fd_sc_hd__nand3_1 _41134_ (.A(_18901_),
    .B(_18915_),
    .C(_18983_),
    .Y(_18984_));
 sky130_fd_sc_hd__xnor2_1 _41135_ (.A(_18982_),
    .B(_18984_),
    .Y(_18985_));
 sky130_fd_sc_hd__nand2_1 _41136_ (.A(_18985_),
    .B(net1224),
    .Y(_18986_));
 sky130_fd_sc_hd__inv_1 _41137_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[22] ),
    .Y(_18987_));
 sky130_fd_sc_hd__o22ai_1 _41138_ (.A1(_07466_),
    .A2(_18927_),
    .B1(_18987_),
    .B2(_18774_),
    .Y(_18988_));
 sky130_fd_sc_hd__inv_1 _41139_ (.A(_18988_),
    .Y(_18989_));
 sky130_fd_sc_hd__a21oi_2 _41140_ (.A1(_18986_),
    .A2(_18989_),
    .B1(net1762),
    .Y(_05334_));
 sky130_fd_sc_hd__inv_1 _41141_ (.A(\inst$top.soc.uart_0._phy.rx.lower.timer[22] ),
    .Y(_18990_));
 sky130_fd_sc_hd__o21ai_0 _41142_ (.A1(_18987_),
    .A2(net1667),
    .B1(_18990_),
    .Y(_18991_));
 sky130_fd_sc_hd__nor2_1 _41143_ (.A(_18971_),
    .B(_18982_),
    .Y(_18992_));
 sky130_fd_sc_hd__nand2_1 _41144_ (.A(_18973_),
    .B(_18992_),
    .Y(_18993_));
 sky130_fd_sc_hd__nor2_1 _41145_ (.A(_18993_),
    .B(_18952_),
    .Y(_18994_));
 sky130_fd_sc_hd__a21oi_1 _41146_ (.A1(_18994_),
    .A2(_18991_),
    .B1(_18825_),
    .Y(_18995_));
 sky130_fd_sc_hd__o21ai_0 _41147_ (.A1(_18991_),
    .A2(_18994_),
    .B1(_18995_),
    .Y(_18996_));
 sky130_fd_sc_hd__inv_1 _41148_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[23] ),
    .Y(_18997_));
 sky130_fd_sc_hd__o22ai_1 _41149_ (.A1(_18990_),
    .A2(_18927_),
    .B1(_18997_),
    .B2(_18774_),
    .Y(_18998_));
 sky130_fd_sc_hd__inv_1 _41150_ (.A(_18998_),
    .Y(_18999_));
 sky130_fd_sc_hd__a21oi_1 _41151_ (.A1(_18996_),
    .A2(_18999_),
    .B1(net1762),
    .Y(_05335_));
 sky130_fd_sc_hd__nor3b_1 _41152_ (.A(_18982_),
    .B(_18991_),
    .C_N(_18983_),
    .Y(_19000_));
 sky130_fd_sc_hd__nand2_1 _41153_ (.A(_18917_),
    .B(_19000_),
    .Y(_19001_));
 sky130_fd_sc_hd__a21oi_1 _41154_ (.A1(_09353_),
    .A2(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[23] ),
    .B1(\inst$top.soc.uart_0._phy.rx.lower.timer[23] ),
    .Y(_19002_));
 sky130_fd_sc_hd__nand2_1 _41155_ (.A(_19001_),
    .B(_19002_),
    .Y(_19003_));
 sky130_fd_sc_hd__nand3b_1 _41156_ (.A_N(_19002_),
    .B(_18917_),
    .C(_19000_),
    .Y(_19004_));
 sky130_fd_sc_hd__nand3_1 _41157_ (.A(_19003_),
    .B(_19004_),
    .C(net1224),
    .Y(_19005_));
 sky130_fd_sc_hd__nand2_1 _41158_ (.A(net1636),
    .B(\inst$top.soc.uart_0._phy.rx.lower.timer[23] ),
    .Y(_19006_));
 sky130_fd_sc_hd__a21oi_2 _41159_ (.A1(_19005_),
    .A2(_19006_),
    .B1(net1762),
    .Y(_05336_));
 sky130_fd_sc_hd__nor2_1 _41160_ (.A(_02721_),
    .B(_18830_),
    .Y(_19007_));
 sky130_fd_sc_hd__nand2_1 _41161_ (.A(_18831_),
    .B(net1835),
    .Y(_19008_));
 sky130_fd_sc_hd__o22ai_1 _41162_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[3] ),
    .A2(net1224),
    .B1(_19007_),
    .B2(_19008_),
    .Y(_19009_));
 sky130_fd_sc_hd__o21ai_0 _41163_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.timer[2] ),
    .A2(_18927_),
    .B1(_18760_),
    .Y(_19010_));
 sky130_fd_sc_hd__a21oi_1 _41164_ (.A1(_19009_),
    .A2(_18927_),
    .B1(_19010_),
    .Y(_05337_));
 sky130_fd_sc_hd__xnor2_1 _41165_ (.A(_18835_),
    .B(_18864_),
    .Y(_19011_));
 sky130_fd_sc_hd__a21oi_1 _41166_ (.A1(net1766),
    .A2(_18832_),
    .B1(net1635),
    .Y(_19012_));
 sky130_fd_sc_hd__o21ai_0 _41167_ (.A1(net1766),
    .A2(_19011_),
    .B1(_19012_),
    .Y(_19013_));
 sky130_fd_sc_hd__a21oi_1 _41168_ (.A1(net1635),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.timer[3] ),
    .B1(net1762),
    .Y(_19014_));
 sky130_fd_sc_hd__nand2_1 _41169_ (.A(_19013_),
    .B(_19014_),
    .Y(_05338_));
 sky130_fd_sc_hd__xnor2_1 _41170_ (.A(_18833_),
    .B(_18887_),
    .Y(_19015_));
 sky130_fd_sc_hd__a21oi_1 _41171_ (.A1(net1766),
    .A2(_18837_),
    .B1(net1635),
    .Y(_19016_));
 sky130_fd_sc_hd__o21ai_0 _41172_ (.A1(net1766),
    .A2(_19015_),
    .B1(_19016_),
    .Y(_19017_));
 sky130_fd_sc_hd__a21oi_1 _41173_ (.A1(net1635),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.timer[4] ),
    .B1(net1762),
    .Y(_19018_));
 sky130_fd_sc_hd__nand2_1 _41174_ (.A(_19017_),
    .B(_19018_),
    .Y(_05339_));
 sky130_fd_sc_hd__nor2_1 _41175_ (.A(_18839_),
    .B(_18865_),
    .Y(_19019_));
 sky130_fd_sc_hd__o21ai_0 _41176_ (.A1(_18840_),
    .A2(_18864_),
    .B1(net1835),
    .Y(_19020_));
 sky130_fd_sc_hd__o22ai_1 _41177_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[6] ),
    .A2(net1224),
    .B1(_19019_),
    .B2(_19020_),
    .Y(_19021_));
 sky130_fd_sc_hd__o21ai_0 _41178_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.timer[5] ),
    .A2(_18927_),
    .B1(_18760_),
    .Y(_19022_));
 sky130_fd_sc_hd__a21oi_1 _41179_ (.A1(_19021_),
    .A2(_18927_),
    .B1(_19022_),
    .Y(_05340_));
 sky130_fd_sc_hd__xnor2_1 _41180_ (.A(_18842_),
    .B(_18841_),
    .Y(_19023_));
 sky130_fd_sc_hd__a21oi_1 _41181_ (.A1(net1766),
    .A2(_18843_),
    .B1(net1635),
    .Y(_19024_));
 sky130_fd_sc_hd__o21ai_0 _41182_ (.A1(net1766),
    .A2(_19023_),
    .B1(_19024_),
    .Y(_19025_));
 sky130_fd_sc_hd__a21oi_1 _41183_ (.A1(net1635),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.timer[6] ),
    .B1(net1762),
    .Y(_19026_));
 sky130_fd_sc_hd__nand2_1 _41184_ (.A(_19025_),
    .B(_19026_),
    .Y(_05341_));
 sky130_fd_sc_hd__nand2_1 _41185_ (.A(_18842_),
    .B(_18839_),
    .Y(_19027_));
 sky130_fd_sc_hd__nor2_1 _41186_ (.A(_19027_),
    .B(_18866_),
    .Y(_19028_));
 sky130_fd_sc_hd__xor2_1 _41187_ (.A(_18844_),
    .B(_19028_),
    .X(_19029_));
 sky130_fd_sc_hd__inv_1 _41188_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[8] ),
    .Y(_19030_));
 sky130_fd_sc_hd__a21oi_1 _41189_ (.A1(_19030_),
    .A2(net1766),
    .B1(net1636),
    .Y(_19031_));
 sky130_fd_sc_hd__o21ai_0 _41190_ (.A1(net1766),
    .A2(_19029_),
    .B1(_19031_),
    .Y(_19032_));
 sky130_fd_sc_hd__a21oi_1 _41191_ (.A1(net1635),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.timer[7] ),
    .B1(net1762),
    .Y(_19033_));
 sky130_fd_sc_hd__nand2_1 _41192_ (.A(_19032_),
    .B(_19033_),
    .Y(_05342_));
 sky130_fd_sc_hd__inv_1 _41193_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[9] ),
    .Y(_19034_));
 sky130_fd_sc_hd__xor2_1 _41194_ (.A(_18848_),
    .B(_18933_),
    .X(_19035_));
 sky130_fd_sc_hd__nand2_1 _41195_ (.A(_19035_),
    .B(net1835),
    .Y(_19036_));
 sky130_fd_sc_hd__o21ai_0 _41196_ (.A1(_19034_),
    .A2(net1835),
    .B1(_19036_),
    .Y(_19037_));
 sky130_fd_sc_hd__a21oi_1 _41197_ (.A1(net1637),
    .A2(_07474_),
    .B1(net1764),
    .Y(_19038_));
 sky130_fd_sc_hd__o21ai_0 _41198_ (.A1(net1637),
    .A2(_19037_),
    .B1(_19038_),
    .Y(_19039_));
 sky130_fd_sc_hd__inv_2 _41199_ (.A(_19039_),
    .Y(_05343_));
 sky130_fd_sc_hd__xor2_1 _41200_ (.A(_18847_),
    .B(_18900_),
    .X(_19040_));
 sky130_fd_sc_hd__nand2_1 _41201_ (.A(_19040_),
    .B(net1835),
    .Y(_19041_));
 sky130_fd_sc_hd__o21ai_0 _41202_ (.A1(_18852_),
    .A2(net1835),
    .B1(_19041_),
    .Y(_19042_));
 sky130_fd_sc_hd__a21oi_1 _41203_ (.A1(net1637),
    .A2(_07470_),
    .B1(net1764),
    .Y(_19043_));
 sky130_fd_sc_hd__o21ai_0 _41204_ (.A1(net1637),
    .A2(_19042_),
    .B1(_19043_),
    .Y(_19044_));
 sky130_fd_sc_hd__inv_2 _41205_ (.A(_19044_),
    .Y(_05344_));
 sky130_fd_sc_hd__nand2_1 _41206_ (.A(\inst$top.soc.uart_0._phy.rx.symbols__valid ),
    .B(\inst$top.soc.uart_0._phy.rx.lower.rdy ),
    .Y(_19045_));
 sky130_fd_sc_hd__nor2_1 _41207_ (.A(net2996),
    .B(_19045_),
    .Y(_05345_));
 sky130_fd_sc_hd__inv_1 _41208_ (.A(\inst$top.soc.uart_0._phy.rx.symbols__payload[0] ),
    .Y(_19046_));
 sky130_fd_sc_hd__inv_1 _41209_ (.A(\inst$top.soc.uart_0._phy.rx.lower.rdy ),
    .Y(_19047_));
 sky130_fd_sc_hd__nor2_1 _41210_ (.A(\inst$top.soc.uart_0._phy.rx.symbols__valid ),
    .B(_19047_),
    .Y(_19048_));
 sky130_fd_sc_hd__inv_1 _41211_ (.A(_19048_),
    .Y(_19049_));
 sky130_fd_sc_hd__o21ai_0 _41213_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.data[0] ),
    .A2(net1761),
    .B1(net2161),
    .Y(_19051_));
 sky130_fd_sc_hd__a21oi_1 _41214_ (.A1(_19046_),
    .A2(net1761),
    .B1(_19051_),
    .Y(_05346_));
 sky130_fd_sc_hd__inv_1 _41215_ (.A(\inst$top.soc.uart_0._phy.rx.symbols__payload[1] ),
    .Y(_19052_));
 sky130_fd_sc_hd__o21ai_0 _41216_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.data[1] ),
    .A2(net1761),
    .B1(net2161),
    .Y(_19053_));
 sky130_fd_sc_hd__a21oi_1 _41217_ (.A1(_19052_),
    .A2(net1761),
    .B1(_19053_),
    .Y(_05347_));
 sky130_fd_sc_hd__inv_1 _41218_ (.A(\inst$top.soc.uart_0._phy.rx.symbols__payload[2] ),
    .Y(_19054_));
 sky130_fd_sc_hd__o21ai_0 _41219_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.data[2] ),
    .A2(net1760),
    .B1(net2161),
    .Y(_19055_));
 sky130_fd_sc_hd__a21oi_1 _41220_ (.A1(_19054_),
    .A2(net1761),
    .B1(_19055_),
    .Y(_05348_));
 sky130_fd_sc_hd__inv_1 _41221_ (.A(\inst$top.soc.uart_0._phy.rx.symbols__payload[3] ),
    .Y(_19056_));
 sky130_fd_sc_hd__o21ai_0 _41222_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.data[3] ),
    .A2(net1760),
    .B1(net2161),
    .Y(_19057_));
 sky130_fd_sc_hd__a21oi_1 _41223_ (.A1(_19056_),
    .A2(net1760),
    .B1(_19057_),
    .Y(_05349_));
 sky130_fd_sc_hd__inv_1 _41224_ (.A(\inst$top.soc.uart_0._phy.rx.symbols__payload[4] ),
    .Y(_19058_));
 sky130_fd_sc_hd__o21ai_0 _41225_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.data[4] ),
    .A2(net1760),
    .B1(net2161),
    .Y(_19059_));
 sky130_fd_sc_hd__a21oi_1 _41226_ (.A1(_19058_),
    .A2(net1760),
    .B1(_19059_),
    .Y(_05350_));
 sky130_fd_sc_hd__inv_1 _41227_ (.A(\inst$top.soc.uart_0._phy.rx.symbols__payload[5] ),
    .Y(_19060_));
 sky130_fd_sc_hd__o21ai_0 _41229_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.data[5] ),
    .A2(net1760),
    .B1(net2162),
    .Y(_19062_));
 sky130_fd_sc_hd__a21oi_1 _41230_ (.A1(_19060_),
    .A2(net1760),
    .B1(_19062_),
    .Y(_05351_));
 sky130_fd_sc_hd__inv_1 _41231_ (.A(\inst$top.soc.uart_0._phy.rx.symbols__payload[6] ),
    .Y(_19063_));
 sky130_fd_sc_hd__o21ai_0 _41232_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.data[6] ),
    .A2(net1760),
    .B1(net2162),
    .Y(_19064_));
 sky130_fd_sc_hd__a21oi_1 _41233_ (.A1(_19063_),
    .A2(net1761),
    .B1(_19064_),
    .Y(_05352_));
 sky130_fd_sc_hd__inv_1 _41234_ (.A(\inst$top.soc.uart_0._phy.rx.symbols__payload[7] ),
    .Y(_19065_));
 sky130_fd_sc_hd__o21ai_0 _41235_ (.A1(\inst$top.soc.uart_0._phy.rx.lower.data[7] ),
    .A2(net1760),
    .B1(net2161),
    .Y(_19066_));
 sky130_fd_sc_hd__a21oi_1 _41236_ (.A1(_19065_),
    .A2(net1760),
    .B1(_19066_),
    .Y(_05353_));
 sky130_fd_sc_hd__nand2_1 _41237_ (.A(_09295_),
    .B(_18038_),
    .Y(_19067_));
 sky130_fd_sc_hd__nand2_1 _41238_ (.A(_17834_),
    .B(_09298_),
    .Y(_19068_));
 sky130_fd_sc_hd__nand3_1 _41239_ (.A(_09332_),
    .B(_09273_),
    .C(_09276_),
    .Y(_19069_));
 sky130_fd_sc_hd__nor3_1 _41240_ (.A(_19068_),
    .B(_18036_),
    .C(_19069_),
    .Y(_19070_));
 sky130_fd_sc_hd__nand4_1 _41241_ (.A(_19070_),
    .B(_09269_),
    .C(_09262_),
    .D(_18039_),
    .Y(_19071_));
 sky130_fd_sc_hd__nor3_1 _41242_ (.A(_19067_),
    .B(_17876_),
    .C(_19071_),
    .Y(_19072_));
 sky130_fd_sc_hd__nand2_1 _41243_ (.A(_19072_),
    .B(_19868_),
    .Y(_19073_));
 sky130_fd_sc_hd__inv_1 _41244_ (.A(_19073_),
    .Y(_19074_));
 sky130_fd_sc_hd__nor2_1 _41245_ (.A(_17851_),
    .B(_18136_),
    .Y(_19075_));
 sky130_fd_sc_hd__nand2_1 _41246_ (.A(_19074_),
    .B(_19075_),
    .Y(_19076_));
 sky130_fd_sc_hd__o211ai_1 _41247_ (.A1(\inst$top.soc.uart_0._phy.rx.symbols__valid ),
    .A2(\inst$top.soc.uart_0._phy.rx.lower.rdy ),
    .B1(net2161),
    .C1(_19076_),
    .Y(_19077_));
 sky130_fd_sc_hd__inv_2 _41248_ (.A(_19077_),
    .Y(_05354_));
 sky130_fd_sc_hd__nor2_1 _41249_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[17] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[16] ),
    .Y(_19078_));
 sky130_fd_sc_hd__inv_1 _41250_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[19] ),
    .Y(_19079_));
 sky130_fd_sc_hd__inv_1 _41251_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[18] ),
    .Y(_19080_));
 sky130_fd_sc_hd__nand3_1 _41252_ (.A(_19078_),
    .B(_19079_),
    .C(_19080_),
    .Y(_19081_));
 sky130_fd_sc_hd__nor2_1 _41253_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[23] ),
    .B(_19081_),
    .Y(_19082_));
 sky130_fd_sc_hd__inv_1 _41254_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[20] ),
    .Y(_19083_));
 sky130_fd_sc_hd__nor2_1 _41255_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[21] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[22] ),
    .Y(_19084_));
 sky130_fd_sc_hd__and3_1 _41256_ (.A(_19082_),
    .B(_19083_),
    .C(_19084_),
    .X(_19085_));
 sky130_fd_sc_hd__nor2_1 _41257_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[9] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[8] ),
    .Y(_19086_));
 sky130_fd_sc_hd__inv_1 _41258_ (.A(_19086_),
    .Y(_19087_));
 sky130_fd_sc_hd__nor2_1 _41259_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[14] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[15] ),
    .Y(_19088_));
 sky130_fd_sc_hd__nor2_1 _41260_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[13] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[12] ),
    .Y(_19089_));
 sky130_fd_sc_hd__nand2_1 _41261_ (.A(_19088_),
    .B(_19089_),
    .Y(_19090_));
 sky130_fd_sc_hd__nor4_1 _41262_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[11] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[10] ),
    .C(_19087_),
    .D(_19090_),
    .Y(_19091_));
 sky130_fd_sc_hd__inv_1 _41263_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[2] ),
    .Y(_19092_));
 sky130_fd_sc_hd__nand2_1 _41264_ (.A(_19092_),
    .B(_02712_),
    .Y(_19093_));
 sky130_fd_sc_hd__nor2_1 _41265_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[3] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[4] ),
    .Y(_19094_));
 sky130_fd_sc_hd__inv_1 _41266_ (.A(_19094_),
    .Y(_19095_));
 sky130_fd_sc_hd__nor2_1 _41267_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[7] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[6] ),
    .Y(_19096_));
 sky130_fd_sc_hd__inv_1 _41268_ (.A(_19096_),
    .Y(_19097_));
 sky130_fd_sc_hd__nor4_1 _41269_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[5] ),
    .B(_19093_),
    .C(_19095_),
    .D(_19097_),
    .Y(_19098_));
 sky130_fd_sc_hd__nand4_1 _41271_ (.A(_19085_),
    .B(_19091_),
    .C(_19098_),
    .D(net2567),
    .Y(_19100_));
 sky130_fd_sc_hd__inv_1 _41272_ (.A(net2567),
    .Y(_19101_));
 sky130_fd_sc_hd__nand2_1 _41273_ (.A(net1992),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb$27 ),
    .Y(_19102_));
 sky130_fd_sc_hd__nand2_1 _41274_ (.A(_19100_),
    .B(_19102_),
    .Y(_19103_));
 sky130_fd_sc_hd__clkinv_1 _41275_ (.A(net1079),
    .Y(_19104_));
 sky130_fd_sc_hd__nand2_1 _41276_ (.A(_19104_),
    .B(\inst$top.soc.uart_0._phy.tx.lower.bitno[0] ),
    .Y(_19105_));
 sky130_fd_sc_hd__o21ai_0 _41279_ (.A1(_19101_),
    .A2(_02702_),
    .B1(net1079),
    .Y(_19108_));
 sky130_fd_sc_hd__inv_1 _41280_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.Config.enable._storage ),
    .Y(_19109_));
 sky130_fd_sc_hd__nor2_1 _41281_ (.A(net2986),
    .B(_19109_),
    .Y(_19110_));
 sky130_fd_sc_hd__clkinv_1 _41282_ (.A(net1852),
    .Y(_19111_));
 sky130_fd_sc_hd__a21oi_1 _41284_ (.A1(_19105_),
    .A2(_19108_),
    .B1(net1759),
    .Y(_05355_));
 sky130_fd_sc_hd__nand2_1 _41285_ (.A(_19104_),
    .B(\inst$top.soc.uart_0._phy.tx.lower.bitno[1] ),
    .Y(_19113_));
 sky130_fd_sc_hd__nor2_1 _41286_ (.A(_19097_),
    .B(_19087_),
    .Y(_19114_));
 sky130_fd_sc_hd__nor2_1 _41287_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[3] ),
    .B(_19093_),
    .Y(_19115_));
 sky130_fd_sc_hd__nor2_1 _41288_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[11] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[10] ),
    .Y(_19116_));
 sky130_fd_sc_hd__nor2_1 _41289_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[5] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[4] ),
    .Y(_19117_));
 sky130_fd_sc_hd__nand4_1 _41290_ (.A(_19114_),
    .B(_19115_),
    .C(_19116_),
    .D(_19117_),
    .Y(_19118_));
 sky130_fd_sc_hd__nor2_1 _41291_ (.A(_19090_),
    .B(_19118_),
    .Y(_19119_));
 sky130_fd_sc_hd__inv_1 _41292_ (.A(_19119_),
    .Y(_19120_));
 sky130_fd_sc_hd__inv_1 _41293_ (.A(_19085_),
    .Y(_19121_));
 sky130_fd_sc_hd__nor3_1 _41294_ (.A(net1992),
    .B(_19120_),
    .C(_19121_),
    .Y(_19122_));
 sky130_fd_sc_hd__inv_1 _41295_ (.A(_02705_),
    .Y(_19123_));
 sky130_fd_sc_hd__nand2_1 _41296_ (.A(_19122_),
    .B(_19123_),
    .Y(_19124_));
 sky130_fd_sc_hd__a21oi_1 _41297_ (.A1(_19113_),
    .A2(_19124_),
    .B1(net1759),
    .Y(_05356_));
 sky130_fd_sc_hd__nand2_1 _41298_ (.A(_19104_),
    .B(\inst$top.soc.uart_0._phy.tx.lower.bitno[2] ),
    .Y(_19125_));
 sky130_fd_sc_hd__xor2_1 _41299_ (.A(\inst$top.soc.uart_0._phy.tx.lower.bitno[2] ),
    .B(_02704_),
    .X(_19126_));
 sky130_fd_sc_hd__nand2_1 _41300_ (.A(_19122_),
    .B(_19126_),
    .Y(_19127_));
 sky130_fd_sc_hd__a21oi_1 _41301_ (.A1(_19125_),
    .A2(_19127_),
    .B1(net1759),
    .Y(_05357_));
 sky130_fd_sc_hd__nor3_1 _41302_ (.A(\inst$top.soc.uart_0._phy.tx.lower.bitno[2] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.bitno[0] ),
    .C(\inst$top.soc.uart_0._phy.tx.lower.bitno[1] ),
    .Y(_19128_));
 sky130_fd_sc_hd__nand2_1 _41303_ (.A(net1079),
    .B(_19128_),
    .Y(_19129_));
 sky130_fd_sc_hd__inv_1 _41304_ (.A(_19102_),
    .Y(_19130_));
 sky130_fd_sc_hd__a21oi_1 _41305_ (.A1(_19129_),
    .A2(\inst$top.soc.uart_0._phy.tx.lower.bitno[3] ),
    .B1(_19130_),
    .Y(_19131_));
 sky130_fd_sc_hd__or2_2 _41306_ (.A(\inst$top.soc.uart_0._phy.tx.lower.bitno[3] ),
    .B(_19129_),
    .X(_19132_));
 sky130_fd_sc_hd__a21oi_1 _41307_ (.A1(_19131_),
    .A2(_19132_),
    .B1(net1759),
    .Y(_05358_));
 sky130_fd_sc_hd__nor2_1 _41308_ (.A(\inst$top.soc.uart_0._phy.tx.lower.bitno[2] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.bitno[3] ),
    .Y(_19133_));
 sky130_fd_sc_hd__nor2_1 _41309_ (.A(net2567),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb$27 ),
    .Y(_19134_));
 sky130_fd_sc_hd__a311oi_1 _41311_ (.A1(_19122_),
    .A2(_02704_),
    .A3(_19133_),
    .B1(net1991),
    .C1(net1758),
    .Y(_05359_));
 sky130_fd_sc_hd__nand2_1 _41312_ (.A(_19122_),
    .B(\inst$top.soc.uart_0._phy.tx.lower.shreg.start ),
    .Y(_19136_));
 sky130_fd_sc_hd__nand2_1 _41314_ (.A(_19100_),
    .B(net598),
    .Y(_19138_));
 sky130_fd_sc_hd__nand3_1 _41315_ (.A(_19136_),
    .B(net1853),
    .C(_19138_),
    .Y(_05360_));
 sky130_fd_sc_hd__nand2_1 _41316_ (.A(_19104_),
    .B(\inst$top.soc.uart_0._phy.tx.lower.shreg.start ),
    .Y(_19139_));
 sky130_fd_sc_hd__nand2_1 _41317_ (.A(_19122_),
    .B(\inst$top.soc.uart_0._phy.tx.lower.shreg[1] ),
    .Y(_19140_));
 sky130_fd_sc_hd__a21oi_1 _41318_ (.A1(_19139_),
    .A2(_19140_),
    .B1(net1759),
    .Y(_05361_));
 sky130_fd_sc_hd__nand2_1 _41320_ (.A(_19101_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[0] ),
    .Y(_19142_));
 sky130_fd_sc_hd__nand2_1 _41321_ (.A(\inst$top.soc.uart_0._phy.tx.lower.fsm_state ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.shreg[2] ),
    .Y(_19143_));
 sky130_fd_sc_hd__o21ai_0 _41322_ (.A1(\inst$top.soc.uart_0._phy.tx.lower.shreg[1] ),
    .A2(net1079),
    .B1(net1853),
    .Y(_19144_));
 sky130_fd_sc_hd__a31oi_1 _41323_ (.A1(net1079),
    .A2(_19142_),
    .A3(_19143_),
    .B1(_19144_),
    .Y(_05362_));
 sky130_fd_sc_hd__nand2_1 _41324_ (.A(net1992),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[1] ),
    .Y(_19145_));
 sky130_fd_sc_hd__nand2_1 _41325_ (.A(net2567),
    .B(\inst$top.soc.uart_0._phy.tx.lower.shreg[3] ),
    .Y(_19146_));
 sky130_fd_sc_hd__nor2_1 _41326_ (.A(\inst$top.soc.uart_0._phy.tx.lower.shreg[2] ),
    .B(net1079),
    .Y(_19147_));
 sky130_fd_sc_hd__a311oi_1 _41327_ (.A1(net1079),
    .A2(_19145_),
    .A3(_19146_),
    .B1(net1758),
    .C1(_19147_),
    .Y(_05363_));
 sky130_fd_sc_hd__nand2_1 _41328_ (.A(net1992),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[2] ),
    .Y(_19148_));
 sky130_fd_sc_hd__nand2_1 _41329_ (.A(net2567),
    .B(\inst$top.soc.uart_0._phy.tx.lower.shreg[4] ),
    .Y(_19149_));
 sky130_fd_sc_hd__o21ai_0 _41330_ (.A1(\inst$top.soc.uart_0._phy.tx.lower.shreg[3] ),
    .A2(net1081),
    .B1(net1852),
    .Y(_19150_));
 sky130_fd_sc_hd__a31oi_1 _41331_ (.A1(net1081),
    .A2(_19148_),
    .A3(_19149_),
    .B1(_19150_),
    .Y(_05364_));
 sky130_fd_sc_hd__nand2_1 _41332_ (.A(net1992),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[3] ),
    .Y(_19151_));
 sky130_fd_sc_hd__nand2_1 _41333_ (.A(net2567),
    .B(\inst$top.soc.uart_0._phy.tx.lower.shreg[5] ),
    .Y(_19152_));
 sky130_fd_sc_hd__o21ai_0 _41334_ (.A1(\inst$top.soc.uart_0._phy.tx.lower.shreg[4] ),
    .A2(net1079),
    .B1(net1852),
    .Y(_19153_));
 sky130_fd_sc_hd__a31oi_1 _41335_ (.A1(net1081),
    .A2(_19151_),
    .A3(_19152_),
    .B1(_19153_),
    .Y(_05365_));
 sky130_fd_sc_hd__nand2_1 _41336_ (.A(net1992),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[4] ),
    .Y(_19154_));
 sky130_fd_sc_hd__nand2_1 _41337_ (.A(net2567),
    .B(\inst$top.soc.uart_0._phy.tx.lower.shreg[6] ),
    .Y(_19155_));
 sky130_fd_sc_hd__o21ai_0 _41338_ (.A1(\inst$top.soc.uart_0._phy.tx.lower.shreg[5] ),
    .A2(net1079),
    .B1(net1852),
    .Y(_19156_));
 sky130_fd_sc_hd__a31oi_1 _41339_ (.A1(net1080),
    .A2(_19154_),
    .A3(_19155_),
    .B1(_19156_),
    .Y(_05366_));
 sky130_fd_sc_hd__nand2_1 _41340_ (.A(net1992),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[5] ),
    .Y(_19157_));
 sky130_fd_sc_hd__nand2_1 _41341_ (.A(net2567),
    .B(\inst$top.soc.uart_0._phy.tx.lower.shreg[7] ),
    .Y(_19158_));
 sky130_fd_sc_hd__o21ai_0 _41342_ (.A1(\inst$top.soc.uart_0._phy.tx.lower.shreg[6] ),
    .A2(net1080),
    .B1(net1852),
    .Y(_19159_));
 sky130_fd_sc_hd__a31oi_1 _41343_ (.A1(net1080),
    .A2(_19157_),
    .A3(_19158_),
    .B1(_19159_),
    .Y(_05367_));
 sky130_fd_sc_hd__nand2_1 _41344_ (.A(net1992),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[6] ),
    .Y(_19160_));
 sky130_fd_sc_hd__nand2_1 _41345_ (.A(net2567),
    .B(\inst$top.soc.uart_0._phy.tx.lower.shreg[8] ),
    .Y(_19161_));
 sky130_fd_sc_hd__o21ai_0 _41346_ (.A1(\inst$top.soc.uart_0._phy.tx.lower.shreg[7] ),
    .A2(net1080),
    .B1(net1852),
    .Y(_19162_));
 sky130_fd_sc_hd__a31oi_1 _41347_ (.A1(net1080),
    .A2(_19160_),
    .A3(_19161_),
    .B1(_19162_),
    .Y(_05368_));
 sky130_fd_sc_hd__nand2_1 _41348_ (.A(net1992),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[7] ),
    .Y(_19163_));
 sky130_fd_sc_hd__nand2_1 _41349_ (.A(net2567),
    .B(\inst$top.soc.uart_0._phy.tx.lower.shreg.stop ),
    .Y(_19164_));
 sky130_fd_sc_hd__o21ai_0 _41350_ (.A1(\inst$top.soc.uart_0._phy.tx.lower.shreg[8] ),
    .A2(net1080),
    .B1(net1852),
    .Y(_19165_));
 sky130_fd_sc_hd__a31oi_1 _41351_ (.A1(net1080),
    .A2(_19163_),
    .A3(_19164_),
    .B1(_19165_),
    .Y(_05369_));
 sky130_fd_sc_hd__o21ai_0 _41352_ (.A1(\inst$top.soc.uart_0._phy.tx.lower.shreg.stop ),
    .A2(_19130_),
    .B1(net1852),
    .Y(_19166_));
 sky130_fd_sc_hd__nor2_1 _41353_ (.A(_19166_),
    .B(_19122_),
    .Y(_05370_));
 sky130_fd_sc_hd__inv_1 _41354_ (.A(net1990),
    .Y(_19167_));
 sky130_fd_sc_hd__nor2_1 _41356_ (.A(_19120_),
    .B(_19121_),
    .Y(_19169_));
 sky130_fd_sc_hd__nor2_1 _41357_ (.A(net1992),
    .B(_19169_),
    .Y(_19170_));
 sky130_fd_sc_hd__a21oi_1 _41359_ (.A1(_19170_),
    .A2(\inst$top.soc.uart_0._phy.tx.lower.timer[0] ),
    .B1(net1991),
    .Y(_19172_));
 sky130_fd_sc_hd__o21ai_0 _41360_ (.A1(_02706_),
    .A2(_19170_),
    .B1(_19172_),
    .Y(_19173_));
 sky130_fd_sc_hd__o211ai_1 _41361_ (.A1(_02710_),
    .A2(_19167_),
    .B1(net1852),
    .C1(_19173_),
    .Y(_05371_));
 sky130_fd_sc_hd__inv_1 _41362_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[10] ),
    .Y(_19174_));
 sky130_fd_sc_hd__inv_1 _41363_ (.A(_19114_),
    .Y(_19175_));
 sky130_fd_sc_hd__nor4_1 _41364_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[5] ),
    .B(_19093_),
    .C(_19095_),
    .D(_19175_),
    .Y(_19176_));
 sky130_fd_sc_hd__xor2_1 _41365_ (.A(_19174_),
    .B(_19176_),
    .X(_19177_));
 sky130_fd_sc_hd__inv_1 _41366_ (.A(net881),
    .Y(_19178_));
 sky130_fd_sc_hd__inv_1 _41368_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[10] ),
    .Y(_19180_));
 sky130_fd_sc_hd__nor2_1 _41369_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[6] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[7] ),
    .Y(_19181_));
 sky130_fd_sc_hd__inv_1 _41370_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[8] ),
    .Y(_19182_));
 sky130_fd_sc_hd__nand2_1 _41371_ (.A(_19181_),
    .B(_19182_),
    .Y(_19183_));
 sky130_fd_sc_hd__nor2_1 _41372_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[9] ),
    .B(_19183_),
    .Y(_19184_));
 sky130_fd_sc_hd__inv_1 _41373_ (.A(_19184_),
    .Y(_19185_));
 sky130_fd_sc_hd__inv_1 _41374_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[2] ),
    .Y(_19186_));
 sky130_fd_sc_hd__nand2_1 _41375_ (.A(_19186_),
    .B(_02708_),
    .Y(_19187_));
 sky130_fd_sc_hd__nor2_1 _41376_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[3] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[4] ),
    .Y(_19188_));
 sky130_fd_sc_hd__inv_1 _41377_ (.A(_19188_),
    .Y(_19189_));
 sky130_fd_sc_hd__nor3_1 _41378_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[5] ),
    .B(_19187_),
    .C(_19189_),
    .Y(_19190_));
 sky130_fd_sc_hd__inv_1 _41379_ (.A(_19190_),
    .Y(_19191_));
 sky130_fd_sc_hd__nor2_1 _41380_ (.A(_19185_),
    .B(_19191_),
    .Y(_19192_));
 sky130_fd_sc_hd__nor2_1 _41381_ (.A(_19180_),
    .B(_19192_),
    .Y(_19193_));
 sky130_fd_sc_hd__inv_1 _41382_ (.A(_19192_),
    .Y(_19194_));
 sky130_fd_sc_hd__nor2_1 _41383_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[10] ),
    .B(_19194_),
    .Y(_19195_));
 sky130_fd_sc_hd__o21ai_0 _41385_ (.A1(_19193_),
    .A2(_19195_),
    .B1(net1081),
    .Y(_19197_));
 sky130_fd_sc_hd__o221ai_1 _41386_ (.A1(_19174_),
    .A2(net1850),
    .B1(_19177_),
    .B2(_19178_),
    .C1(_19197_),
    .Y(_19198_));
 sky130_fd_sc_hd__nand2_1 _41388_ (.A(_19198_),
    .B(net1853),
    .Y(_19200_));
 sky130_fd_sc_hd__inv_2 _41389_ (.A(_19200_),
    .Y(_05372_));
 sky130_fd_sc_hd__nor2_1 _41390_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[2] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[1] ),
    .Y(_19201_));
 sky130_fd_sc_hd__inv_1 _41391_ (.A(_19201_),
    .Y(_19202_));
 sky130_fd_sc_hd__nor3_1 _41392_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[0] ),
    .B(_19095_),
    .C(_19202_),
    .Y(_19203_));
 sky130_fd_sc_hd__nor2_1 _41393_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[7] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[8] ),
    .Y(_19204_));
 sky130_fd_sc_hd__nor2_1 _41394_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[5] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[6] ),
    .Y(_19205_));
 sky130_fd_sc_hd__nor2_1 _41395_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[9] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[10] ),
    .Y(_19206_));
 sky130_fd_sc_hd__nand4_1 _41396_ (.A(_19203_),
    .B(_19204_),
    .C(_19205_),
    .D(_19206_),
    .Y(_19207_));
 sky130_fd_sc_hd__xor2_1 _41397_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[11] ),
    .B(_19207_),
    .X(_19208_));
 sky130_fd_sc_hd__nor2_1 _41398_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[2] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[1] ),
    .Y(_19209_));
 sky130_fd_sc_hd__nor2_1 _41399_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[7] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[8] ),
    .Y(_19210_));
 sky130_fd_sc_hd__nand3_1 _41400_ (.A(_19188_),
    .B(_19209_),
    .C(_19210_),
    .Y(_19211_));
 sky130_fd_sc_hd__nor3_1 _41401_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[5] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[6] ),
    .C(_19211_),
    .Y(_19212_));
 sky130_fd_sc_hd__nor2_1 _41402_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[9] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[10] ),
    .Y(_19213_));
 sky130_fd_sc_hd__nand3_1 _41403_ (.A(_19212_),
    .B(_02706_),
    .C(_19213_),
    .Y(_19214_));
 sky130_fd_sc_hd__xor2_1 _41404_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[11] ),
    .B(_19214_),
    .X(_19215_));
 sky130_fd_sc_hd__nand2_1 _41405_ (.A(net1990),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[11] ),
    .Y(_19216_));
 sky130_fd_sc_hd__o221ai_1 _41406_ (.A1(_19208_),
    .A2(net864),
    .B1(_19215_),
    .B2(_19104_),
    .C1(_19216_),
    .Y(_19217_));
 sky130_fd_sc_hd__nand2_1 _41407_ (.A(_19217_),
    .B(net1853),
    .Y(_19218_));
 sky130_fd_sc_hd__inv_2 _41408_ (.A(_19218_),
    .Y(_05373_));
 sky130_fd_sc_hd__inv_1 _41409_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[12] ),
    .Y(_19219_));
 sky130_fd_sc_hd__xor2_1 _41410_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[12] ),
    .B(_19118_),
    .X(_19220_));
 sky130_fd_sc_hd__inv_1 _41411_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[12] ),
    .Y(_19221_));
 sky130_fd_sc_hd__nor2_1 _41412_ (.A(_19183_),
    .B(_19191_),
    .Y(_19222_));
 sky130_fd_sc_hd__inv_1 _41413_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[11] ),
    .Y(_19223_));
 sky130_fd_sc_hd__nand3_1 _41414_ (.A(_19222_),
    .B(_19223_),
    .C(_19213_),
    .Y(_19224_));
 sky130_fd_sc_hd__xor2_1 _41415_ (.A(_19221_),
    .B(_19224_),
    .X(_19225_));
 sky130_fd_sc_hd__nand2_1 _41416_ (.A(_19225_),
    .B(net1081),
    .Y(_19226_));
 sky130_fd_sc_hd__o221ai_1 _41417_ (.A1(_19219_),
    .A2(net1850),
    .B1(_19220_),
    .B2(_19178_),
    .C1(_19226_),
    .Y(_19227_));
 sky130_fd_sc_hd__nand2_1 _41418_ (.A(_19227_),
    .B(net1853),
    .Y(_19228_));
 sky130_fd_sc_hd__inv_2 _41419_ (.A(_19228_),
    .Y(_05374_));
 sky130_fd_sc_hd__inv_1 _41420_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[13] ),
    .Y(_19229_));
 sky130_fd_sc_hd__nor2_1 _41421_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[11] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[12] ),
    .Y(_19230_));
 sky130_fd_sc_hd__nand4_1 _41422_ (.A(_19212_),
    .B(_02706_),
    .C(_19213_),
    .D(_19230_),
    .Y(_19231_));
 sky130_fd_sc_hd__xor2_1 _41423_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[13] ),
    .B(_19231_),
    .X(_19232_));
 sky130_fd_sc_hd__nor2_1 _41424_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[11] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[12] ),
    .Y(_19233_));
 sky130_fd_sc_hd__nand2_1 _41425_ (.A(_19206_),
    .B(_19233_),
    .Y(_19234_));
 sky130_fd_sc_hd__inv_1 _41426_ (.A(_19234_),
    .Y(_19235_));
 sky130_fd_sc_hd__nand4_1 _41427_ (.A(_19203_),
    .B(_19204_),
    .C(_19205_),
    .D(_19235_),
    .Y(_19236_));
 sky130_fd_sc_hd__xor2_1 _41428_ (.A(_19229_),
    .B(_19236_),
    .X(_19237_));
 sky130_fd_sc_hd__nand2_1 _41429_ (.A(net881),
    .B(_19237_),
    .Y(_19238_));
 sky130_fd_sc_hd__o221ai_1 _41430_ (.A1(_19229_),
    .A2(net1850),
    .B1(_19232_),
    .B2(_19104_),
    .C1(_19238_),
    .Y(_19239_));
 sky130_fd_sc_hd__nand2_1 _41431_ (.A(_19239_),
    .B(net1853),
    .Y(_19240_));
 sky130_fd_sc_hd__inv_2 _41432_ (.A(_19240_),
    .Y(_05375_));
 sky130_fd_sc_hd__nand3_1 _41433_ (.A(_19176_),
    .B(_19116_),
    .C(_19089_),
    .Y(_19241_));
 sky130_fd_sc_hd__xor2_1 _41434_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[14] ),
    .B(_19241_),
    .X(_19242_));
 sky130_fd_sc_hd__nand2_1 _41435_ (.A(net1990),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[14] ),
    .Y(_19243_));
 sky130_fd_sc_hd__nor2_1 _41436_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[12] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[13] ),
    .Y(_19244_));
 sky130_fd_sc_hd__nand3_1 _41437_ (.A(_19244_),
    .B(_19180_),
    .C(_19223_),
    .Y(_19245_));
 sky130_fd_sc_hd__nor2_1 _41438_ (.A(_19245_),
    .B(_19194_),
    .Y(_19246_));
 sky130_fd_sc_hd__inv_1 _41439_ (.A(_19246_),
    .Y(_19247_));
 sky130_fd_sc_hd__inv_1 _41440_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[14] ),
    .Y(_19248_));
 sky130_fd_sc_hd__nand2_1 _41441_ (.A(_19247_),
    .B(_19248_),
    .Y(_19249_));
 sky130_fd_sc_hd__nand2_1 _41442_ (.A(_19246_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[14] ),
    .Y(_19250_));
 sky130_fd_sc_hd__nand3_1 _41443_ (.A(net1078),
    .B(_19249_),
    .C(_19250_),
    .Y(_19251_));
 sky130_fd_sc_hd__o211ai_1 _41444_ (.A1(net864),
    .A2(_19242_),
    .B1(_19243_),
    .C1(_19251_),
    .Y(_19252_));
 sky130_fd_sc_hd__nand2_1 _41445_ (.A(_19252_),
    .B(net1851),
    .Y(_19253_));
 sky130_fd_sc_hd__inv_2 _41446_ (.A(_19253_),
    .Y(_05376_));
 sky130_fd_sc_hd__inv_1 _41447_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[15] ),
    .Y(_19254_));
 sky130_fd_sc_hd__nor2_1 _41448_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[13] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[14] ),
    .Y(_19255_));
 sky130_fd_sc_hd__inv_1 _41449_ (.A(_19255_),
    .Y(_19256_));
 sky130_fd_sc_hd__nor3_1 _41450_ (.A(_19254_),
    .B(_19256_),
    .C(_19236_),
    .Y(_19257_));
 sky130_fd_sc_hd__o21ai_0 _41451_ (.A1(_19256_),
    .A2(_19236_),
    .B1(_19254_),
    .Y(_19258_));
 sky130_fd_sc_hd__nand2_1 _41452_ (.A(net881),
    .B(_19258_),
    .Y(_19259_));
 sky130_fd_sc_hd__nor2_1 _41453_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[13] ),
    .B(_19231_),
    .Y(_19260_));
 sky130_fd_sc_hd__inv_1 _41454_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[15] ),
    .Y(_19261_));
 sky130_fd_sc_hd__a21oi_1 _41455_ (.A1(_19260_),
    .A2(_19248_),
    .B1(_19261_),
    .Y(_19262_));
 sky130_fd_sc_hd__nor4_1 _41456_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[13] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[14] ),
    .C(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[15] ),
    .D(_19231_),
    .Y(_19263_));
 sky130_fd_sc_hd__o21ai_0 _41457_ (.A1(_19262_),
    .A2(_19263_),
    .B1(net1078),
    .Y(_19264_));
 sky130_fd_sc_hd__o221ai_1 _41458_ (.A1(_19254_),
    .A2(net1850),
    .B1(_19257_),
    .B2(_19259_),
    .C1(_19264_),
    .Y(_19265_));
 sky130_fd_sc_hd__nand2_1 _41459_ (.A(_19265_),
    .B(net1851),
    .Y(_19266_));
 sky130_fd_sc_hd__inv_2 _41460_ (.A(_19266_),
    .Y(_05377_));
 sky130_fd_sc_hd__inv_1 _41461_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[16] ),
    .Y(_19267_));
 sky130_fd_sc_hd__xor2_1 _41462_ (.A(_19267_),
    .B(_19119_),
    .X(_19268_));
 sky130_fd_sc_hd__nor2_1 _41463_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[14] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[15] ),
    .Y(_19269_));
 sky130_fd_sc_hd__nand2_1 _41464_ (.A(_19244_),
    .B(_19269_),
    .Y(_19270_));
 sky130_fd_sc_hd__nor2_1 _41465_ (.A(_19270_),
    .B(_19224_),
    .Y(_19271_));
 sky130_fd_sc_hd__xor2_1 _41466_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[16] ),
    .B(_19271_),
    .X(_19272_));
 sky130_fd_sc_hd__nand2_1 _41467_ (.A(_19272_),
    .B(net1078),
    .Y(_19273_));
 sky130_fd_sc_hd__o221ai_1 _41468_ (.A1(_19267_),
    .A2(net1850),
    .B1(_19268_),
    .B2(net864),
    .C1(_19273_),
    .Y(_19274_));
 sky130_fd_sc_hd__nand2_1 _41469_ (.A(_19274_),
    .B(net1851),
    .Y(_19275_));
 sky130_fd_sc_hd__inv_2 _41470_ (.A(_19275_),
    .Y(_05378_));
 sky130_fd_sc_hd__inv_1 _41471_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[17] ),
    .Y(_19276_));
 sky130_fd_sc_hd__nand2_1 _41472_ (.A(_19088_),
    .B(_19267_),
    .Y(_19277_));
 sky130_fd_sc_hd__nor3_1 _41473_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[13] ),
    .B(_19277_),
    .C(_19236_),
    .Y(_19278_));
 sky130_fd_sc_hd__xor2_1 _41474_ (.A(_19276_),
    .B(_19278_),
    .X(_19279_));
 sky130_fd_sc_hd__inv_1 _41475_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[16] ),
    .Y(_19280_));
 sky130_fd_sc_hd__nand2_1 _41476_ (.A(_19263_),
    .B(_19280_),
    .Y(_19281_));
 sky130_fd_sc_hd__nor2_1 _41477_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[17] ),
    .B(_19281_),
    .Y(_19282_));
 sky130_fd_sc_hd__inv_1 _41478_ (.A(_19282_),
    .Y(_19283_));
 sky130_fd_sc_hd__nand2_1 _41479_ (.A(_19281_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[17] ),
    .Y(_19284_));
 sky130_fd_sc_hd__nand2_1 _41480_ (.A(_19283_),
    .B(_19284_),
    .Y(_19285_));
 sky130_fd_sc_hd__nand2_1 _41481_ (.A(_19285_),
    .B(net1078),
    .Y(_19286_));
 sky130_fd_sc_hd__o221ai_1 _41482_ (.A1(_19276_),
    .A2(net1850),
    .B1(net864),
    .B2(_19279_),
    .C1(_19286_),
    .Y(_19287_));
 sky130_fd_sc_hd__nand2_1 _41483_ (.A(_19287_),
    .B(net1851),
    .Y(_19288_));
 sky130_fd_sc_hd__inv_2 _41484_ (.A(_19288_),
    .Y(_05379_));
 sky130_fd_sc_hd__nor3_1 _41485_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[17] ),
    .B(_19277_),
    .C(_19241_),
    .Y(_19289_));
 sky130_fd_sc_hd__xor2_1 _41486_ (.A(_19080_),
    .B(_19289_),
    .X(_19290_));
 sky130_fd_sc_hd__nor2_1 _41487_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[16] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[17] ),
    .Y(_19291_));
 sky130_fd_sc_hd__nand2_1 _41488_ (.A(_19269_),
    .B(_19291_),
    .Y(_19292_));
 sky130_fd_sc_hd__nor2_1 _41489_ (.A(_19292_),
    .B(_19247_),
    .Y(_19293_));
 sky130_fd_sc_hd__xor2_1 _41490_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[18] ),
    .B(_19293_),
    .X(_19294_));
 sky130_fd_sc_hd__nand2_1 _41491_ (.A(_19294_),
    .B(net1078),
    .Y(_19295_));
 sky130_fd_sc_hd__o221ai_1 _41492_ (.A1(_19080_),
    .A2(net1850),
    .B1(net864),
    .B2(_19290_),
    .C1(_19295_),
    .Y(_19296_));
 sky130_fd_sc_hd__nand2_1 _41493_ (.A(_19296_),
    .B(net1851),
    .Y(_19297_));
 sky130_fd_sc_hd__inv_2 _41494_ (.A(_19297_),
    .Y(_05380_));
 sky130_fd_sc_hd__inv_1 _41495_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[19] ),
    .Y(_19298_));
 sky130_fd_sc_hd__o21ai_0 _41496_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[18] ),
    .A2(_19283_),
    .B1(_19298_),
    .Y(_19299_));
 sky130_fd_sc_hd__nor2_1 _41497_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[18] ),
    .B(_19283_),
    .Y(_19300_));
 sky130_fd_sc_hd__nand2_1 _41498_ (.A(_19300_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[19] ),
    .Y(_19301_));
 sky130_fd_sc_hd__nand3_1 _41499_ (.A(_19278_),
    .B(_19276_),
    .C(_19080_),
    .Y(_19302_));
 sky130_fd_sc_hd__xor2_1 _41500_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[19] ),
    .B(_19302_),
    .X(_19303_));
 sky130_fd_sc_hd__o22ai_1 _41501_ (.A1(_19079_),
    .A2(net1850),
    .B1(net864),
    .B2(_19303_),
    .Y(_19304_));
 sky130_fd_sc_hd__a31oi_1 _41502_ (.A1(_19299_),
    .A2(_19301_),
    .A3(net1078),
    .B1(_19304_),
    .Y(_19305_));
 sky130_fd_sc_hd__nor2_1 _41503_ (.A(net1758),
    .B(_19305_),
    .Y(_05381_));
 sky130_fd_sc_hd__o21ai_0 _41504_ (.A1(\inst$top.soc.uart_0._phy.tx.lower.timer[1] ),
    .A2(net1850),
    .B1(net1852),
    .Y(_19306_));
 sky130_fd_sc_hd__a221oi_1 _41505_ (.A1(_19170_),
    .A2(_02713_),
    .B1(net1080),
    .B2(_02709_),
    .C1(_19306_),
    .Y(_05382_));
 sky130_fd_sc_hd__nor2_1 _41506_ (.A(_19081_),
    .B(_19120_),
    .Y(_19307_));
 sky130_fd_sc_hd__xor2_1 _41507_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[20] ),
    .B(_19307_),
    .X(_19308_));
 sky130_fd_sc_hd__a22oi_1 _41508_ (.A1(\inst$top.soc.uart_0._phy.tx.lower.timer[20] ),
    .A2(net1990),
    .B1(_19308_),
    .B2(net881),
    .Y(_19309_));
 sky130_fd_sc_hd__inv_1 _41509_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[20] ),
    .Y(_19310_));
 sky130_fd_sc_hd__nor2_1 _41510_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[18] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[19] ),
    .Y(_19311_));
 sky130_fd_sc_hd__nand3_1 _41511_ (.A(_19271_),
    .B(_19291_),
    .C(_19311_),
    .Y(_19312_));
 sky130_fd_sc_hd__xor2_1 _41512_ (.A(_19310_),
    .B(_19312_),
    .X(_19313_));
 sky130_fd_sc_hd__nand2_1 _41513_ (.A(_19313_),
    .B(net1078),
    .Y(_19314_));
 sky130_fd_sc_hd__nand2_1 _41514_ (.A(_19309_),
    .B(_19314_),
    .Y(_19315_));
 sky130_fd_sc_hd__nand2_1 _41515_ (.A(_19315_),
    .B(net1851),
    .Y(_19316_));
 sky130_fd_sc_hd__inv_2 _41516_ (.A(_19316_),
    .Y(_05383_));
 sky130_fd_sc_hd__inv_1 _41517_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[21] ),
    .Y(_19317_));
 sky130_fd_sc_hd__inv_1 _41518_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[18] ),
    .Y(_19318_));
 sky130_fd_sc_hd__nor2_1 _41519_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[19] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[20] ),
    .Y(_19319_));
 sky130_fd_sc_hd__nand3_1 _41520_ (.A(_19282_),
    .B(_19318_),
    .C(_19319_),
    .Y(_19320_));
 sky130_fd_sc_hd__xor2_1 _41521_ (.A(_19317_),
    .B(_19320_),
    .X(_19321_));
 sky130_fd_sc_hd__nand2_1 _41522_ (.A(_19321_),
    .B(net1078),
    .Y(_19322_));
 sky130_fd_sc_hd__nor3_1 _41523_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[19] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[20] ),
    .C(_19302_),
    .Y(_19323_));
 sky130_fd_sc_hd__xor2_1 _41524_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[21] ),
    .B(_19323_),
    .X(_19324_));
 sky130_fd_sc_hd__a22oi_1 _41525_ (.A1(\inst$top.soc.uart_0._phy.tx.lower.timer[21] ),
    .A2(net1990),
    .B1(_19324_),
    .B2(net881),
    .Y(_19325_));
 sky130_fd_sc_hd__nand2_1 _41526_ (.A(_19322_),
    .B(_19325_),
    .Y(_19326_));
 sky130_fd_sc_hd__nand2_1 _41527_ (.A(_19326_),
    .B(net1851),
    .Y(_19327_));
 sky130_fd_sc_hd__inv_2 _41528_ (.A(_19327_),
    .Y(_05384_));
 sky130_fd_sc_hd__inv_1 _41529_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[22] ),
    .Y(_19328_));
 sky130_fd_sc_hd__inv_1 _41530_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[22] ),
    .Y(_19329_));
 sky130_fd_sc_hd__nand4_1 _41531_ (.A(_19293_),
    .B(_19310_),
    .C(_19317_),
    .D(_19311_),
    .Y(_19330_));
 sky130_fd_sc_hd__xor2_1 _41532_ (.A(_19329_),
    .B(_19330_),
    .X(_19331_));
 sky130_fd_sc_hd__nand2_1 _41533_ (.A(_19331_),
    .B(net1078),
    .Y(_19332_));
 sky130_fd_sc_hd__nor3_1 _41534_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[19] ),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[21] ),
    .C(\inst$top.soc.uart_0._phy.tx.lower.timer[20] ),
    .Y(_19333_));
 sky130_fd_sc_hd__nand3_1 _41535_ (.A(_19289_),
    .B(_19080_),
    .C(_19333_),
    .Y(_19334_));
 sky130_fd_sc_hd__xor2_1 _41536_ (.A(_19328_),
    .B(_19334_),
    .X(_19335_));
 sky130_fd_sc_hd__nand2_1 _41537_ (.A(_19335_),
    .B(net881),
    .Y(_19336_));
 sky130_fd_sc_hd__o211ai_1 _41538_ (.A1(_19328_),
    .A2(net1850),
    .B1(_19332_),
    .C1(_19336_),
    .Y(_19337_));
 sky130_fd_sc_hd__nand2_1 _41539_ (.A(_19337_),
    .B(net1851),
    .Y(_19338_));
 sky130_fd_sc_hd__inv_2 _41540_ (.A(_19338_),
    .Y(_05385_));
 sky130_fd_sc_hd__nand2_1 _41541_ (.A(_19323_),
    .B(_19084_),
    .Y(_19339_));
 sky130_fd_sc_hd__xnor2_1 _41542_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[23] ),
    .B(_19339_),
    .Y(_19340_));
 sky130_fd_sc_hd__inv_1 _41543_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[23] ),
    .Y(_19341_));
 sky130_fd_sc_hd__nand4_1 _41544_ (.A(_19300_),
    .B(_19317_),
    .C(_19329_),
    .D(_19319_),
    .Y(_19342_));
 sky130_fd_sc_hd__o21ai_0 _41545_ (.A1(_19341_),
    .A2(_19342_),
    .B1(net1078),
    .Y(_19343_));
 sky130_fd_sc_hd__a21oi_1 _41546_ (.A1(_19341_),
    .A2(_19342_),
    .B1(_19343_),
    .Y(_19344_));
 sky130_fd_sc_hd__a221oi_1 _41547_ (.A1(\inst$top.soc.uart_0._phy.tx.lower.timer[23] ),
    .A2(net1990),
    .B1(net881),
    .B2(_19340_),
    .C1(_19344_),
    .Y(_19345_));
 sky130_fd_sc_hd__nor2_1 _41548_ (.A(net1758),
    .B(_19345_),
    .Y(_05386_));
 sky130_fd_sc_hd__xor2_1 _41549_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[2] ),
    .B(_02712_),
    .X(_19346_));
 sky130_fd_sc_hd__xor2_1 _41550_ (.A(_02708_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[2] ),
    .X(_19347_));
 sky130_fd_sc_hd__nor2_1 _41551_ (.A(_19092_),
    .B(_19167_),
    .Y(_19348_));
 sky130_fd_sc_hd__a221oi_1 _41552_ (.A1(net881),
    .A2(_19346_),
    .B1(net1079),
    .B2(_19347_),
    .C1(_19348_),
    .Y(_19349_));
 sky130_fd_sc_hd__nor2_1 _41553_ (.A(net1758),
    .B(_19349_),
    .Y(_05387_));
 sky130_fd_sc_hd__nor2_1 _41554_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[0] ),
    .B(_19202_),
    .Y(_19350_));
 sky130_fd_sc_hd__xnor2_1 _41555_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[3] ),
    .B(_19350_),
    .Y(_19351_));
 sky130_fd_sc_hd__nand2_1 _41556_ (.A(_19209_),
    .B(_02706_),
    .Y(_19352_));
 sky130_fd_sc_hd__xnor2_1 _41557_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[3] ),
    .B(_19352_),
    .Y(_19353_));
 sky130_fd_sc_hd__nand2_1 _41558_ (.A(net1080),
    .B(_19353_),
    .Y(_19354_));
 sky130_fd_sc_hd__a21oi_1 _41559_ (.A1(net1991),
    .A2(\inst$top.soc.uart_0._phy.tx.lower.timer[3] ),
    .B1(net1758),
    .Y(_19355_));
 sky130_fd_sc_hd__o211ai_1 _41560_ (.A1(_19351_),
    .A2(_19178_),
    .B1(_19354_),
    .C1(_19355_),
    .Y(_05388_));
 sky130_fd_sc_hd__o21ai_0 _41561_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[3] ),
    .A2(_19187_),
    .B1(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[4] ),
    .Y(_19356_));
 sky130_fd_sc_hd__o21ai_0 _41562_ (.A1(_19187_),
    .A2(_19189_),
    .B1(_19356_),
    .Y(_19357_));
 sky130_fd_sc_hd__nand2_1 _41563_ (.A(net1081),
    .B(_19357_),
    .Y(_19358_));
 sky130_fd_sc_hd__xor2_1 _41564_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[4] ),
    .B(_19115_),
    .X(_19359_));
 sky130_fd_sc_hd__nand2_1 _41565_ (.A(net881),
    .B(_19359_),
    .Y(_19360_));
 sky130_fd_sc_hd__a21oi_1 _41566_ (.A1(net1990),
    .A2(\inst$top.soc.uart_0._phy.tx.lower.timer[4] ),
    .B1(net1758),
    .Y(_19361_));
 sky130_fd_sc_hd__nand3_1 _41567_ (.A(_19358_),
    .B(_19360_),
    .C(_19361_),
    .Y(_05389_));
 sky130_fd_sc_hd__nand2_1 _41568_ (.A(_19188_),
    .B(_19209_),
    .Y(_19362_));
 sky130_fd_sc_hd__nor2_1 _41569_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[0] ),
    .B(_19362_),
    .Y(_19363_));
 sky130_fd_sc_hd__xor2_1 _41570_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[5] ),
    .B(_19363_),
    .X(_19364_));
 sky130_fd_sc_hd__nand2_1 _41571_ (.A(net1080),
    .B(_19364_),
    .Y(_19365_));
 sky130_fd_sc_hd__xor2_1 _41572_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[5] ),
    .B(_19203_),
    .X(_19366_));
 sky130_fd_sc_hd__nand2_1 _41573_ (.A(net881),
    .B(_19366_),
    .Y(_19367_));
 sky130_fd_sc_hd__nand2_1 _41574_ (.A(net1990),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[5] ),
    .Y(_19368_));
 sky130_fd_sc_hd__a31oi_1 _41575_ (.A1(_19365_),
    .A2(_19367_),
    .A3(_19368_),
    .B1(net1758),
    .Y(_05390_));
 sky130_fd_sc_hd__nor3_1 _41576_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[5] ),
    .B(_19093_),
    .C(_19095_),
    .Y(_19369_));
 sky130_fd_sc_hd__xnor2_1 _41577_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[6] ),
    .B(_19369_),
    .Y(_19370_));
 sky130_fd_sc_hd__xnor2_1 _41578_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[6] ),
    .B(_19190_),
    .Y(_19371_));
 sky130_fd_sc_hd__a21oi_1 _41579_ (.A1(net1991),
    .A2(\inst$top.soc.uart_0._phy.tx.lower.timer[6] ),
    .B1(net1758),
    .Y(_19372_));
 sky130_fd_sc_hd__o221ai_1 _41580_ (.A1(_19370_),
    .A2(net864),
    .B1(_19371_),
    .B2(_19104_),
    .C1(_19372_),
    .Y(_05391_));
 sky130_fd_sc_hd__nand3_1 _41581_ (.A(_19350_),
    .B(_19094_),
    .C(_19205_),
    .Y(_19373_));
 sky130_fd_sc_hd__xor2_1 _41582_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[7] ),
    .B(_19373_),
    .X(_19374_));
 sky130_fd_sc_hd__nor4_1 _41583_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[0] ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[5] ),
    .C(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[6] ),
    .D(_19362_),
    .Y(_19375_));
 sky130_fd_sc_hd__xnor2_1 _41584_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[7] ),
    .B(_19375_),
    .Y(_19376_));
 sky130_fd_sc_hd__a21oi_1 _41585_ (.A1(net1991),
    .A2(\inst$top.soc.uart_0._phy.tx.lower.timer[7] ),
    .B1(net1758),
    .Y(_19377_));
 sky130_fd_sc_hd__o221ai_1 _41586_ (.A1(_19374_),
    .A2(net864),
    .B1(_19376_),
    .B2(_19104_),
    .C1(_19377_),
    .Y(_05392_));
 sky130_fd_sc_hd__xnor2_1 _41587_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[8] ),
    .B(_19098_),
    .Y(_19378_));
 sky130_fd_sc_hd__nand2_1 _41588_ (.A(net1990),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[8] ),
    .Y(_19379_));
 sky130_fd_sc_hd__a21oi_1 _41589_ (.A1(_19190_),
    .A2(_19181_),
    .B1(_19182_),
    .Y(_19380_));
 sky130_fd_sc_hd__o21ai_0 _41590_ (.A1(_19222_),
    .A2(_19380_),
    .B1(net1081),
    .Y(_19381_));
 sky130_fd_sc_hd__o211ai_1 _41591_ (.A1(_19378_),
    .A2(net864),
    .B1(_19379_),
    .C1(_19381_),
    .Y(_19382_));
 sky130_fd_sc_hd__nand2_1 _41592_ (.A(_19382_),
    .B(net1851),
    .Y(_19383_));
 sky130_fd_sc_hd__inv_2 _41593_ (.A(_19383_),
    .Y(_05393_));
 sky130_fd_sc_hd__nand3_1 _41594_ (.A(_19094_),
    .B(_19204_),
    .C(_19205_),
    .Y(_19384_));
 sky130_fd_sc_hd__nor3_1 _41595_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[0] ),
    .B(_19202_),
    .C(_19384_),
    .Y(_19385_));
 sky130_fd_sc_hd__xnor2_1 _41596_ (.A(\inst$top.soc.uart_0._phy.tx.lower.timer[9] ),
    .B(_19385_),
    .Y(_19386_));
 sky130_fd_sc_hd__nand2_1 _41597_ (.A(_19212_),
    .B(_02706_),
    .Y(_19387_));
 sky130_fd_sc_hd__xor2_1 _41598_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[9] ),
    .B(_19387_),
    .X(_19388_));
 sky130_fd_sc_hd__nand2_1 _41599_ (.A(net1990),
    .B(\inst$top.soc.uart_0._phy.tx.lower.timer[9] ),
    .Y(_19389_));
 sky130_fd_sc_hd__o221ai_1 _41600_ (.A1(_19386_),
    .A2(net864),
    .B1(_19388_),
    .B2(_19104_),
    .C1(_19389_),
    .Y(_19390_));
 sky130_fd_sc_hd__nand2_1 _41601_ (.A(_19390_),
    .B(net1851),
    .Y(_19391_));
 sky130_fd_sc_hd__inv_2 _41602_ (.A(_19391_),
    .Y(_05394_));
 sky130_fd_sc_hd__nor2_1 _41603_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb ),
    .B(_18759_),
    .Y(_19392_));
 sky130_fd_sc_hd__a21oi_1 _41604_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.Config.enable.port__w_data ),
    .A2(\inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb ),
    .B1(_19392_),
    .Y(_19393_));
 sky130_fd_sc_hd__nor2_1 _41605_ (.A(net2997),
    .B(_19393_),
    .Y(_05395_));
 sky130_fd_sc_hd__nand2_1 _41606_ (.A(_18759_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb$34 ),
    .Y(_19394_));
 sky130_fd_sc_hd__inv_2 _41608_ (.A(net1846),
    .Y(_19396_));
 sky130_fd_sc_hd__nand2_1 _41609_ (.A(_19396_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.Config.enable.port__w_data ),
    .Y(_19397_));
 sky130_fd_sc_hd__o211ai_1 _41610_ (.A1(_07464_),
    .A2(_19396_),
    .B1(net2159),
    .C1(_19397_),
    .Y(_05396_));
 sky130_fd_sc_hd__o21ai_0 _41613_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[2] ),
    .A2(net1849),
    .B1(net2166),
    .Y(_19400_));
 sky130_fd_sc_hd__a21oi_1 _41614_ (.A1(_18852_),
    .A2(net1848),
    .B1(_19400_),
    .Y(_05397_));
 sky130_fd_sc_hd__o21ai_0 _41615_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[3] ),
    .A2(net1849),
    .B1(net2166),
    .Y(_19401_));
 sky130_fd_sc_hd__a21oi_1 _41616_ (.A1(_18869_),
    .A2(net1848),
    .B1(_19401_),
    .Y(_05398_));
 sky130_fd_sc_hd__o21ai_0 _41617_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[4] ),
    .A2(net1849),
    .B1(net2166),
    .Y(_19402_));
 sky130_fd_sc_hd__a21oi_1 _41618_ (.A1(_18879_),
    .A2(net1848),
    .B1(_19402_),
    .Y(_05399_));
 sky130_fd_sc_hd__o21ai_0 _41619_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[5] ),
    .A2(net1849),
    .B1(net2165),
    .Y(_19403_));
 sky130_fd_sc_hd__a21oi_1 _41620_ (.A1(_18894_),
    .A2(net1848),
    .B1(_19403_),
    .Y(_05400_));
 sky130_fd_sc_hd__o21ai_0 _41621_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[6] ),
    .A2(net1848),
    .B1(net2162),
    .Y(_19404_));
 sky130_fd_sc_hd__a21oi_1 _41622_ (.A1(_18906_),
    .A2(net1848),
    .B1(_19404_),
    .Y(_05401_));
 sky130_fd_sc_hd__o21ai_0 _41623_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[7] ),
    .A2(net1849),
    .B1(net2165),
    .Y(_19405_));
 sky130_fd_sc_hd__a21oi_1 _41624_ (.A1(_18918_),
    .A2(net1848),
    .B1(_19405_),
    .Y(_05402_));
 sky130_fd_sc_hd__o21ai_0 _41625_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[0] ),
    .A2(net1847),
    .B1(net2161),
    .Y(_19406_));
 sky130_fd_sc_hd__a21oi_1 _41626_ (.A1(_18928_),
    .A2(net1847),
    .B1(_19406_),
    .Y(_05403_));
 sky130_fd_sc_hd__o21ai_0 _41628_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[1] ),
    .A2(net1845),
    .B1(net2134),
    .Y(_19408_));
 sky130_fd_sc_hd__a21oi_1 _41629_ (.A1(_18936_),
    .A2(net1845),
    .B1(_19408_),
    .Y(_05404_));
 sky130_fd_sc_hd__o21ai_0 _41630_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[2] ),
    .A2(net1845),
    .B1(net2134),
    .Y(_19409_));
 sky130_fd_sc_hd__a21oi_1 _41631_ (.A1(_18946_),
    .A2(net1845),
    .B1(_19409_),
    .Y(_05405_));
 sky130_fd_sc_hd__o21ai_0 _41633_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[3] ),
    .A2(net1847),
    .B1(net2162),
    .Y(_19411_));
 sky130_fd_sc_hd__a21oi_1 _41634_ (.A1(_18959_),
    .A2(net1847),
    .B1(_19411_),
    .Y(_05406_));
 sky130_fd_sc_hd__o21ai_0 _41635_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.Status.overflow.port__w_data ),
    .A2(net1846),
    .B1(net2159),
    .Y(_19412_));
 sky130_fd_sc_hd__a21oi_1 _41636_ (.A1(_18824_),
    .A2(net1846),
    .B1(_19412_),
    .Y(_05407_));
 sky130_fd_sc_hd__o21ai_0 _41637_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[4] ),
    .A2(net1847),
    .B1(net2159),
    .Y(_19413_));
 sky130_fd_sc_hd__a21oi_1 _41638_ (.A1(_18965_),
    .A2(net1847),
    .B1(_19413_),
    .Y(_05408_));
 sky130_fd_sc_hd__o21ai_0 _41639_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[5] ),
    .A2(net1845),
    .B1(net2160),
    .Y(_19414_));
 sky130_fd_sc_hd__a21oi_1 _41640_ (.A1(_18981_),
    .A2(net1845),
    .B1(_19414_),
    .Y(_05409_));
 sky130_fd_sc_hd__o21ai_0 _41641_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[6] ),
    .A2(net1845),
    .B1(net2133),
    .Y(_19415_));
 sky130_fd_sc_hd__a21oi_1 _41642_ (.A1(_18987_),
    .A2(net1845),
    .B1(_19415_),
    .Y(_05410_));
 sky130_fd_sc_hd__o21ai_0 _41643_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[7] ),
    .A2(net1845),
    .B1(net2160),
    .Y(_19416_));
 sky130_fd_sc_hd__a21oi_1 _41644_ (.A1(_18997_),
    .A2(net1845),
    .B1(_19416_),
    .Y(_05411_));
 sky130_fd_sc_hd__o21ai_0 _41645_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.Status.error.port__w_data ),
    .A2(net1846),
    .B1(net2159),
    .Y(_19417_));
 sky130_fd_sc_hd__a21oi_1 _41646_ (.A1(_18828_),
    .A2(net1846),
    .B1(_19417_),
    .Y(_05412_));
 sky130_fd_sc_hd__nand2_1 _41647_ (.A(_19396_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[3] ),
    .Y(_19418_));
 sky130_fd_sc_hd__o211ai_1 _41648_ (.A1(_18834_),
    .A2(_19396_),
    .B1(net2160),
    .C1(_19418_),
    .Y(_05413_));
 sky130_fd_sc_hd__nand2_1 _41649_ (.A(_19396_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[4] ),
    .Y(_19419_));
 sky130_fd_sc_hd__o211ai_1 _41650_ (.A1(_18832_),
    .A2(_19396_),
    .B1(net2159),
    .C1(_19419_),
    .Y(_05414_));
 sky130_fd_sc_hd__o21ai_0 _41651_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[5] ),
    .A2(net1846),
    .B1(net2133),
    .Y(_19420_));
 sky130_fd_sc_hd__a21oi_1 _41652_ (.A1(_18837_),
    .A2(net1846),
    .B1(_19420_),
    .Y(_05415_));
 sky130_fd_sc_hd__nand2_1 _41653_ (.A(_19396_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[6] ),
    .Y(_19421_));
 sky130_fd_sc_hd__nand2_1 _41654_ (.A(net1846),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[6] ),
    .Y(_19422_));
 sky130_fd_sc_hd__nand3_1 _41655_ (.A(_19421_),
    .B(_19422_),
    .C(net2160),
    .Y(_05416_));
 sky130_fd_sc_hd__nand2_1 _41656_ (.A(_19396_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[7] ),
    .Y(_19423_));
 sky130_fd_sc_hd__o211ai_1 _41657_ (.A1(_18843_),
    .A2(_19396_),
    .B1(net2159),
    .C1(_19423_),
    .Y(_05417_));
 sky130_fd_sc_hd__o21ai_0 _41659_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[0] ),
    .A2(net1848),
    .B1(net2166),
    .Y(_19425_));
 sky130_fd_sc_hd__a21oi_1 _41660_ (.A1(_19030_),
    .A2(net1849),
    .B1(_19425_),
    .Y(_05418_));
 sky130_fd_sc_hd__o21ai_0 _41661_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[1] ),
    .A2(net1848),
    .B1(net2166),
    .Y(_19426_));
 sky130_fd_sc_hd__a21oi_1 _41662_ (.A1(_19034_),
    .A2(net1848),
    .B1(_19426_),
    .Y(_05419_));
 sky130_fd_sc_hd__nand2_1 _41663_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.Status.error.port__w_data ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb$25 ),
    .Y(_19427_));
 sky130_fd_sc_hd__a21oi_1 _41664_ (.A1(_19427_),
    .A2(\inst$top.soc.uart_0._uart.rx.bridge.Status.error._storage ),
    .B1(\inst$top.soc.uart_0._phy.rx.err.frame ),
    .Y(_19428_));
 sky130_fd_sc_hd__nor2_1 _41665_ (.A(net2995),
    .B(_19428_),
    .Y(_05420_));
 sky130_fd_sc_hd__nand2_1 _41666_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb$25 ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.Status.overflow.port__w_data ),
    .Y(_19429_));
 sky130_fd_sc_hd__a21oi_1 _41667_ (.A1(_19429_),
    .A2(\inst$top.soc.uart_0._uart.rx.bridge.Status.overflow._storage ),
    .B1(\inst$top.soc.uart_0._phy.rx.overflow ),
    .Y(_19430_));
 sky130_fd_sc_hd__nor2_1 _41668_ (.A(net2997),
    .B(_19430_),
    .Y(_05421_));
 sky130_fd_sc_hd__nor2_1 _41669_ (.A(_19067_),
    .B(_19071_),
    .Y(_19431_));
 sky130_fd_sc_hd__nand2_1 _41670_ (.A(_19431_),
    .B(_17866_),
    .Y(_19432_));
 sky130_fd_sc_hd__nor2_1 _41671_ (.A(\inst$top.soc.bus__adr[2] ),
    .B(_19432_),
    .Y(_19433_));
 sky130_fd_sc_hd__inv_1 _41672_ (.A(_19433_),
    .Y(_19434_));
 sky130_fd_sc_hd__nor3_1 _41673_ (.A(net2987),
    .B(_18138_),
    .C(_19434_),
    .Y(_05422_));
 sky130_fd_sc_hd__nand2_1 _41674_ (.A(_17869_),
    .B(_17832_),
    .Y(_19435_));
 sky130_fd_sc_hd__nor2_1 _41675_ (.A(_19435_),
    .B(_19434_),
    .Y(_05423_));
 sky130_fd_sc_hd__nor2_1 _41676_ (.A(_18044_),
    .B(_19434_),
    .Y(_05424_));
 sky130_fd_sc_hd__nor2_1 _41677_ (.A(_17885_),
    .B(_18149_),
    .Y(_19436_));
 sky130_fd_sc_hd__inv_1 _41678_ (.A(_19436_),
    .Y(_19437_));
 sky130_fd_sc_hd__nor2_1 _41679_ (.A(_19437_),
    .B(_19073_),
    .Y(_19438_));
 sky130_fd_sc_hd__nor2_2 _41680_ (.A(_18096_),
    .B(_19073_),
    .Y(_19439_));
 sky130_fd_sc_hd__nand2_1 _41681_ (.A(net804),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[0] ),
    .Y(_19440_));
 sky130_fd_sc_hd__nand3_1 _41682_ (.A(_19074_),
    .B(\inst$top.soc.uart_0._phy.rx.symbols__valid ),
    .C(_18137_),
    .Y(_19441_));
 sky130_fd_sc_hd__o2111ai_1 _41683_ (.A1(_18759_),
    .A2(_17887_),
    .B1(_19438_),
    .C1(_19440_),
    .D1(_19441_),
    .Y(_19442_));
 sky130_fd_sc_hd__o211ai_1 _41684_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[0] ),
    .A2(_19438_),
    .B1(net2159),
    .C1(_19442_),
    .Y(_19443_));
 sky130_fd_sc_hd__inv_2 _41685_ (.A(_19443_),
    .Y(_05425_));
 sky130_fd_sc_hd__nand2_1 _41686_ (.A(_18137_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.Status.overflow._storage ),
    .Y(_19444_));
 sky130_fd_sc_hd__nand2_1 _41687_ (.A(_18095_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[1] ),
    .Y(_19445_));
 sky130_fd_sc_hd__nor3_1 _41688_ (.A(_09314_),
    .B(_09261_),
    .C(_19068_),
    .Y(_19446_));
 sky130_fd_sc_hd__nor2_1 _41689_ (.A(\inst$top.soc.bus__adr[7] ),
    .B(_09317_),
    .Y(_19447_));
 sky130_fd_sc_hd__nand3_1 _41690_ (.A(_19446_),
    .B(_17841_),
    .C(_19447_),
    .Y(_19448_));
 sky130_fd_sc_hd__nor3_1 _41691_ (.A(_18035_),
    .B(_17838_),
    .C(_19069_),
    .Y(_19449_));
 sky130_fd_sc_hd__nor2_1 _41692_ (.A(_09259_),
    .B(_09294_),
    .Y(_19450_));
 sky130_fd_sc_hd__nand4_1 _41693_ (.A(_19449_),
    .B(_09325_),
    .C(_09287_),
    .D(_19450_),
    .Y(_19451_));
 sky130_fd_sc_hd__nor3_1 _41694_ (.A(_17876_),
    .B(_19448_),
    .C(_19451_),
    .Y(_19452_));
 sky130_fd_sc_hd__nand2_1 _41695_ (.A(_19452_),
    .B(_19868_),
    .Y(_19453_));
 sky130_fd_sc_hd__nor2_1 _41696_ (.A(_19437_),
    .B(_19453_),
    .Y(_19454_));
 sky130_fd_sc_hd__o21ai_0 _41697_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[1] ),
    .A2(_19454_),
    .B1(net2135),
    .Y(_19455_));
 sky130_fd_sc_hd__a31oi_1 _41698_ (.A1(_19438_),
    .A2(_19444_),
    .A3(_19445_),
    .B1(_19455_),
    .Y(_05426_));
 sky130_fd_sc_hd__nand2_1 _41699_ (.A(_18137_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.Status.error._storage ),
    .Y(_19456_));
 sky130_fd_sc_hd__nand2_1 _41700_ (.A(_18095_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[2] ),
    .Y(_19457_));
 sky130_fd_sc_hd__o21ai_0 _41701_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[2] ),
    .A2(_19454_),
    .B1(net2135),
    .Y(_19458_));
 sky130_fd_sc_hd__a31oi_1 _41702_ (.A1(_19438_),
    .A2(_19456_),
    .A3(_19457_),
    .B1(_19458_),
    .Y(_05427_));
 sky130_fd_sc_hd__inv_1 _41703_ (.A(_19438_),
    .Y(_19459_));
 sky130_fd_sc_hd__nand2_1 _41704_ (.A(_19459_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[3] ),
    .Y(_19460_));
 sky130_fd_sc_hd__nand2_1 _41706_ (.A(net805),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[3] ),
    .Y(_19462_));
 sky130_fd_sc_hd__a21oi_2 _41707_ (.A1(_19460_),
    .A2(_19462_),
    .B1(net2995),
    .Y(_05428_));
 sky130_fd_sc_hd__nand2_1 _41708_ (.A(_19459_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[4] ),
    .Y(_19463_));
 sky130_fd_sc_hd__nand2_1 _41709_ (.A(net805),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[4] ),
    .Y(_19464_));
 sky130_fd_sc_hd__a21oi_2 _41710_ (.A1(_19463_),
    .A2(_19464_),
    .B1(net2997),
    .Y(_05429_));
 sky130_fd_sc_hd__nand2_1 _41711_ (.A(_19459_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[5] ),
    .Y(_19465_));
 sky130_fd_sc_hd__nand2_1 _41712_ (.A(net804),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[5] ),
    .Y(_19466_));
 sky130_fd_sc_hd__a21oi_1 _41713_ (.A1(_19465_),
    .A2(_19466_),
    .B1(net2995),
    .Y(_05430_));
 sky130_fd_sc_hd__nand2_1 _41714_ (.A(_19459_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[6] ),
    .Y(_19467_));
 sky130_fd_sc_hd__nand2_1 _41715_ (.A(net804),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[6] ),
    .Y(_19468_));
 sky130_fd_sc_hd__a21oi_1 _41716_ (.A1(_19467_),
    .A2(_19468_),
    .B1(net2995),
    .Y(_05431_));
 sky130_fd_sc_hd__nand2_1 _41717_ (.A(_19459_),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[7] ),
    .Y(_19469_));
 sky130_fd_sc_hd__nand2_1 _41718_ (.A(net804),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[7] ),
    .Y(_19470_));
 sky130_fd_sc_hd__a21oi_1 _41719_ (.A1(_19469_),
    .A2(_19470_),
    .B1(net2995),
    .Y(_05432_));
 sky130_fd_sc_hd__nand2_1 _41720_ (.A(_19074_),
    .B(net2135),
    .Y(_19471_));
 sky130_fd_sc_hd__nor2_1 _41721_ (.A(_19437_),
    .B(_19471_),
    .Y(_05433_));
 sky130_fd_sc_hd__nor2_1 _41723_ (.A(_18096_),
    .B(_19453_),
    .Y(_19473_));
 sky130_fd_sc_hd__a31oi_1 _41724_ (.A1(_19868_),
    .A2(_19075_),
    .A3(_19452_),
    .B1(_19473_),
    .Y(_19474_));
 sky130_fd_sc_hd__inv_1 _41725_ (.A(net804),
    .Y(_19475_));
 sky130_fd_sc_hd__o22ai_1 _41726_ (.A1(_19046_),
    .A2(_19076_),
    .B1(_19030_),
    .B2(_19475_),
    .Y(_19476_));
 sky130_fd_sc_hd__a21oi_1 _41727_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[0] ),
    .A2(_19474_),
    .B1(_19476_),
    .Y(_19477_));
 sky130_fd_sc_hd__nor2_1 _41728_ (.A(net2996),
    .B(_19477_),
    .Y(_05434_));
 sky130_fd_sc_hd__o22ai_1 _41729_ (.A1(_19052_),
    .A2(_19076_),
    .B1(_19034_),
    .B2(_19475_),
    .Y(_19478_));
 sky130_fd_sc_hd__a21oi_1 _41730_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[1] ),
    .A2(_19474_),
    .B1(_19478_),
    .Y(_19479_));
 sky130_fd_sc_hd__nor2_1 _41731_ (.A(net2995),
    .B(_19479_),
    .Y(_05435_));
 sky130_fd_sc_hd__o22ai_1 _41732_ (.A1(_19054_),
    .A2(_19076_),
    .B1(_18852_),
    .B2(_19475_),
    .Y(_19480_));
 sky130_fd_sc_hd__a21oi_1 _41733_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[2] ),
    .A2(_19474_),
    .B1(_19480_),
    .Y(_19481_));
 sky130_fd_sc_hd__nor2_1 _41734_ (.A(net2987),
    .B(_19481_),
    .Y(_05436_));
 sky130_fd_sc_hd__o22ai_1 _41735_ (.A1(_19056_),
    .A2(_19076_),
    .B1(_18869_),
    .B2(_19475_),
    .Y(_19482_));
 sky130_fd_sc_hd__a21oi_1 _41736_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[3] ),
    .A2(_19474_),
    .B1(_19482_),
    .Y(_19483_));
 sky130_fd_sc_hd__nor2_1 _41737_ (.A(net2996),
    .B(_19483_),
    .Y(_05437_));
 sky130_fd_sc_hd__o22ai_1 _41738_ (.A1(_19058_),
    .A2(_19076_),
    .B1(_18879_),
    .B2(_19475_),
    .Y(_19484_));
 sky130_fd_sc_hd__a21oi_1 _41739_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[4] ),
    .A2(_19474_),
    .B1(_19484_),
    .Y(_19485_));
 sky130_fd_sc_hd__nor2_1 _41740_ (.A(net2996),
    .B(_19485_),
    .Y(_05438_));
 sky130_fd_sc_hd__o22ai_1 _41741_ (.A1(_19060_),
    .A2(_19076_),
    .B1(_18894_),
    .B2(_19475_),
    .Y(_19486_));
 sky130_fd_sc_hd__a21oi_1 _41742_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[5] ),
    .A2(_19474_),
    .B1(_19486_),
    .Y(_19487_));
 sky130_fd_sc_hd__nor2_1 _41743_ (.A(net2987),
    .B(_19487_),
    .Y(_05439_));
 sky130_fd_sc_hd__o22ai_1 _41744_ (.A1(_19063_),
    .A2(_19076_),
    .B1(_18906_),
    .B2(_19475_),
    .Y(_19488_));
 sky130_fd_sc_hd__a21oi_1 _41745_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[6] ),
    .A2(_19474_),
    .B1(_19488_),
    .Y(_19489_));
 sky130_fd_sc_hd__nor2_1 _41746_ (.A(net2996),
    .B(_19489_),
    .Y(_05440_));
 sky130_fd_sc_hd__o22ai_1 _41747_ (.A1(_19065_),
    .A2(_19076_),
    .B1(_18918_),
    .B2(_19475_),
    .Y(_19490_));
 sky130_fd_sc_hd__a21oi_1 _41748_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[7] ),
    .A2(_19474_),
    .B1(_19490_),
    .Y(_19491_));
 sky130_fd_sc_hd__nor2_2 _41749_ (.A(net2995),
    .B(_19491_),
    .Y(_05441_));
 sky130_fd_sc_hd__inv_1 _41750_ (.A(_19075_),
    .Y(_19492_));
 sky130_fd_sc_hd__nand2_1 _41751_ (.A(_17984_),
    .B(_19492_),
    .Y(_19493_));
 sky130_fd_sc_hd__inv_1 _41752_ (.A(_19493_),
    .Y(_19494_));
 sky130_fd_sc_hd__nor2_1 _41753_ (.A(_19494_),
    .B(_19471_),
    .Y(_05442_));
 sky130_fd_sc_hd__o21ai_0 _41754_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[0] ),
    .A2(_19473_),
    .B1(net2160),
    .Y(_19495_));
 sky130_fd_sc_hd__a21oi_1 _41755_ (.A1(_18928_),
    .A2(net805),
    .B1(_19495_),
    .Y(_05443_));
 sky130_fd_sc_hd__o21ai_0 _41756_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[1] ),
    .A2(_19473_),
    .B1(net2135),
    .Y(_19496_));
 sky130_fd_sc_hd__a21oi_1 _41757_ (.A1(_18936_),
    .A2(net804),
    .B1(_19496_),
    .Y(_05444_));
 sky130_fd_sc_hd__o21ai_0 _41758_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[2] ),
    .A2(_19473_),
    .B1(net2135),
    .Y(_19497_));
 sky130_fd_sc_hd__a21oi_1 _41759_ (.A1(_18946_),
    .A2(net804),
    .B1(_19497_),
    .Y(_05445_));
 sky130_fd_sc_hd__o21ai_0 _41760_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[3] ),
    .A2(_19473_),
    .B1(net2161),
    .Y(_19498_));
 sky130_fd_sc_hd__a21oi_1 _41761_ (.A1(_18959_),
    .A2(net805),
    .B1(_19498_),
    .Y(_05446_));
 sky130_fd_sc_hd__o21ai_0 _41762_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[4] ),
    .A2(_19473_),
    .B1(net2159),
    .Y(_19499_));
 sky130_fd_sc_hd__a21oi_1 _41763_ (.A1(_18965_),
    .A2(net805),
    .B1(_19499_),
    .Y(_05447_));
 sky130_fd_sc_hd__o21ai_0 _41764_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[5] ),
    .A2(_19473_),
    .B1(net2135),
    .Y(_19500_));
 sky130_fd_sc_hd__a21oi_1 _41765_ (.A1(_18981_),
    .A2(net804),
    .B1(_19500_),
    .Y(_05448_));
 sky130_fd_sc_hd__o21ai_0 _41766_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[6] ),
    .A2(_19473_),
    .B1(net2135),
    .Y(_19501_));
 sky130_fd_sc_hd__a21oi_2 _41767_ (.A1(_18987_),
    .A2(net804),
    .B1(_19501_),
    .Y(_05449_));
 sky130_fd_sc_hd__o21ai_0 _41768_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[7] ),
    .A2(_19473_),
    .B1(net2159),
    .Y(_19502_));
 sky130_fd_sc_hd__a21oi_2 _41769_ (.A1(_18997_),
    .A2(net804),
    .B1(_19502_),
    .Y(_05450_));
 sky130_fd_sc_hd__nor2_1 _41770_ (.A(_17856_),
    .B(_17870_),
    .Y(_19503_));
 sky130_fd_sc_hd__inv_1 _41771_ (.A(_19503_),
    .Y(_19504_));
 sky130_fd_sc_hd__nor2_1 _41772_ (.A(_19504_),
    .B(_19471_),
    .Y(_05451_));
 sky130_fd_sc_hd__nor2_1 _41773_ (.A(_19437_),
    .B(_19434_),
    .Y(_19505_));
 sky130_fd_sc_hd__o21ai_0 _41776_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.Config.enable.port__w_data ),
    .A2(net803),
    .B1(net2139),
    .Y(_19508_));
 sky130_fd_sc_hd__a21oi_2 _41777_ (.A1(net900),
    .A2(net803),
    .B1(_19508_),
    .Y(_05452_));
 sky130_fd_sc_hd__o21ai_0 _41778_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.Status.overflow.port__w_data ),
    .A2(net803),
    .B1(net2163),
    .Y(_19509_));
 sky130_fd_sc_hd__a21oi_2 _41779_ (.A1(net868),
    .A2(net803),
    .B1(_19509_),
    .Y(_05453_));
 sky130_fd_sc_hd__o21ai_0 _41780_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.Status.error.port__w_data ),
    .A2(net802),
    .B1(net2159),
    .Y(_19510_));
 sky130_fd_sc_hd__a21oi_2 _41781_ (.A1(_17954_),
    .A2(net803),
    .B1(_19510_),
    .Y(_05454_));
 sky130_fd_sc_hd__o21ai_0 _41782_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[3] ),
    .A2(net802),
    .B1(net2160),
    .Y(_19511_));
 sky130_fd_sc_hd__a21oi_2 _41783_ (.A1(_17960_),
    .A2(net802),
    .B1(_19511_),
    .Y(_05455_));
 sky130_fd_sc_hd__o21ai_0 _41784_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[4] ),
    .A2(net802),
    .B1(net2163),
    .Y(_19512_));
 sky130_fd_sc_hd__a21oi_2 _41785_ (.A1(net867),
    .A2(net803),
    .B1(_19512_),
    .Y(_05456_));
 sky130_fd_sc_hd__o21ai_0 _41786_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[5] ),
    .A2(net802),
    .B1(net2134),
    .Y(_19513_));
 sky130_fd_sc_hd__a21oi_2 _41787_ (.A1(_17972_),
    .A2(net802),
    .B1(_19513_),
    .Y(_05457_));
 sky130_fd_sc_hd__o21ai_0 _41788_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[6] ),
    .A2(net802),
    .B1(net2160),
    .Y(_19514_));
 sky130_fd_sc_hd__a21oi_2 _41789_ (.A1(_17977_),
    .A2(net802),
    .B1(_19514_),
    .Y(_05458_));
 sky130_fd_sc_hd__nor2_1 _41790_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[7] ),
    .B(net802),
    .Y(_19515_));
 sky130_fd_sc_hd__a211oi_2 _41791_ (.A1(net802),
    .A2(_17982_),
    .B1(net2995),
    .C1(_19515_),
    .Y(_05459_));
 sky130_fd_sc_hd__nor3b_1 _41792_ (.A(_19448_),
    .B(_19451_),
    .C_N(_18187_),
    .Y(_19516_));
 sky130_fd_sc_hd__nand2_1 _41793_ (.A(_19516_),
    .B(_19868_),
    .Y(_19517_));
 sky130_fd_sc_hd__nor2_1 _41794_ (.A(_17984_),
    .B(_19517_),
    .Y(_19518_));
 sky130_fd_sc_hd__nor2_1 _41796_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[0] ),
    .B(net825),
    .Y(_19520_));
 sky130_fd_sc_hd__a211oi_2 _41797_ (.A1(net825),
    .A2(net900),
    .B1(net2999),
    .C1(_19520_),
    .Y(_05460_));
 sky130_fd_sc_hd__nor2_1 _41798_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[1] ),
    .B(net826),
    .Y(_19521_));
 sky130_fd_sc_hd__a211oi_2 _41799_ (.A1(net826),
    .A2(net868),
    .B1(net2999),
    .C1(_19521_),
    .Y(_05461_));
 sky130_fd_sc_hd__nor2_1 _41800_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[2] ),
    .B(net825),
    .Y(_19522_));
 sky130_fd_sc_hd__a211oi_2 _41801_ (.A1(net826),
    .A2(_17954_),
    .B1(net2999),
    .C1(_19522_),
    .Y(_05462_));
 sky130_fd_sc_hd__nor2_1 _41802_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[3] ),
    .B(net825),
    .Y(_19523_));
 sky130_fd_sc_hd__a211oi_2 _41803_ (.A1(net825),
    .A2(_17960_),
    .B1(net2999),
    .C1(_19523_),
    .Y(_05463_));
 sky130_fd_sc_hd__nor2_1 _41805_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[4] ),
    .B(net825),
    .Y(_19525_));
 sky130_fd_sc_hd__a211oi_2 _41806_ (.A1(net825),
    .A2(net867),
    .B1(net2999),
    .C1(_19525_),
    .Y(_05464_));
 sky130_fd_sc_hd__nor2_1 _41807_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[5] ),
    .B(net825),
    .Y(_19526_));
 sky130_fd_sc_hd__a211oi_2 _41808_ (.A1(net826),
    .A2(_17972_),
    .B1(net3003),
    .C1(_19526_),
    .Y(_05465_));
 sky130_fd_sc_hd__nor2_1 _41809_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[6] ),
    .B(net826),
    .Y(_19527_));
 sky130_fd_sc_hd__a211oi_2 _41810_ (.A1(net826),
    .A2(_17977_),
    .B1(net2996),
    .C1(_19527_),
    .Y(_05466_));
 sky130_fd_sc_hd__nor2_1 _41811_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[7] ),
    .B(net825),
    .Y(_19528_));
 sky130_fd_sc_hd__a211oi_2 _41812_ (.A1(net825),
    .A2(_17982_),
    .B1(net3000),
    .C1(_19528_),
    .Y(_05467_));
 sky130_fd_sc_hd__nor2_1 _41813_ (.A(_19504_),
    .B(_19434_),
    .Y(_19529_));
 sky130_fd_sc_hd__o21ai_0 _41815_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[0] ),
    .A2(net801),
    .B1(net2161),
    .Y(_19531_));
 sky130_fd_sc_hd__a21oi_2 _41816_ (.A1(net900),
    .A2(net801),
    .B1(_19531_),
    .Y(_05468_));
 sky130_fd_sc_hd__o21ai_0 _41817_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[1] ),
    .A2(net800),
    .B1(net2134),
    .Y(_19532_));
 sky130_fd_sc_hd__a21oi_2 _41818_ (.A1(net868),
    .A2(net800),
    .B1(_19532_),
    .Y(_05469_));
 sky130_fd_sc_hd__o21ai_0 _41819_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[2] ),
    .A2(net800),
    .B1(net2134),
    .Y(_19533_));
 sky130_fd_sc_hd__a21oi_2 _41820_ (.A1(_17954_),
    .A2(net800),
    .B1(_19533_),
    .Y(_05470_));
 sky130_fd_sc_hd__o21ai_0 _41822_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[3] ),
    .A2(net801),
    .B1(net2162),
    .Y(_19535_));
 sky130_fd_sc_hd__a21oi_2 _41823_ (.A1(_17960_),
    .A2(net801),
    .B1(_19535_),
    .Y(_05471_));
 sky130_fd_sc_hd__o21ai_0 _41824_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[4] ),
    .A2(net801),
    .B1(net2160),
    .Y(_19536_));
 sky130_fd_sc_hd__a21oi_2 _41825_ (.A1(net867),
    .A2(net801),
    .B1(_19536_),
    .Y(_05472_));
 sky130_fd_sc_hd__o21ai_0 _41826_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[5] ),
    .A2(net800),
    .B1(net2160),
    .Y(_19537_));
 sky130_fd_sc_hd__a21oi_2 _41827_ (.A1(_17972_),
    .A2(net800),
    .B1(_19537_),
    .Y(_05473_));
 sky130_fd_sc_hd__o21ai_0 _41828_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[6] ),
    .A2(net800),
    .B1(net2134),
    .Y(_19538_));
 sky130_fd_sc_hd__a21oi_2 _41829_ (.A1(_17977_),
    .A2(net800),
    .B1(_19538_),
    .Y(_05474_));
 sky130_fd_sc_hd__nor2_1 _41830_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[7] ),
    .B(net800),
    .Y(_19539_));
 sky130_fd_sc_hd__a211oi_2 _41831_ (.A1(net800),
    .A2(_17982_),
    .B1(net2995),
    .C1(_19539_),
    .Y(_05475_));
 sky130_fd_sc_hd__nor2_1 _41832_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb ),
    .B(_19109_),
    .Y(_19540_));
 sky130_fd_sc_hd__a21oi_1 _41833_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.Config.enable.port__w_data ),
    .A2(\inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb ),
    .B1(_19540_),
    .Y(_19541_));
 sky130_fd_sc_hd__nor2_1 _41834_ (.A(net2987),
    .B(_19541_),
    .Y(_05476_));
 sky130_fd_sc_hd__nand2_1 _41835_ (.A(_19109_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb$32 ),
    .Y(_19542_));
 sky130_fd_sc_hd__clkinv_1 _41836_ (.A(net1844),
    .Y(_19543_));
 sky130_fd_sc_hd__nand2_1 _41837_ (.A(_19543_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.Config.enable.port__w_data ),
    .Y(_19544_));
 sky130_fd_sc_hd__o211ai_1 _41838_ (.A1(_02706_),
    .A2(_19543_),
    .B1(net2132),
    .C1(_19544_),
    .Y(_05477_));
 sky130_fd_sc_hd__o21ai_0 _41842_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[2] ),
    .A2(net1843),
    .B1(net2133),
    .Y(_19548_));
 sky130_fd_sc_hd__a21oi_1 _41843_ (.A1(_19180_),
    .A2(net1842),
    .B1(_19548_),
    .Y(_05478_));
 sky130_fd_sc_hd__o21ai_0 _41844_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[3] ),
    .A2(net1843),
    .B1(net2133),
    .Y(_19549_));
 sky130_fd_sc_hd__a21oi_1 _41845_ (.A1(_19223_),
    .A2(net1842),
    .B1(_19549_),
    .Y(_05479_));
 sky130_fd_sc_hd__o21ai_0 _41846_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[4] ),
    .A2(net1843),
    .B1(net2132),
    .Y(_19550_));
 sky130_fd_sc_hd__a21oi_1 _41847_ (.A1(_19221_),
    .A2(net1844),
    .B1(_19550_),
    .Y(_05480_));
 sky130_fd_sc_hd__nor2_1 _41848_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[13] ),
    .B(_19543_),
    .Y(_19551_));
 sky130_fd_sc_hd__o21ai_0 _41849_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[5] ),
    .A2(net1844),
    .B1(net2132),
    .Y(_19552_));
 sky130_fd_sc_hd__nor2_1 _41850_ (.A(_19551_),
    .B(_19552_),
    .Y(_05481_));
 sky130_fd_sc_hd__o21ai_0 _41851_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[6] ),
    .A2(_19542_),
    .B1(net2122),
    .Y(_19553_));
 sky130_fd_sc_hd__a21oi_1 _41852_ (.A1(_19248_),
    .A2(net1842),
    .B1(_19553_),
    .Y(_05482_));
 sky130_fd_sc_hd__o21ai_0 _41853_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[7] ),
    .A2(net1844),
    .B1(net2132),
    .Y(_19554_));
 sky130_fd_sc_hd__a21oi_1 _41854_ (.A1(_19261_),
    .A2(net1842),
    .B1(_19554_),
    .Y(_05483_));
 sky130_fd_sc_hd__o21ai_0 _41855_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[0] ),
    .A2(_19542_),
    .B1(net2122),
    .Y(_19555_));
 sky130_fd_sc_hd__a21oi_1 _41856_ (.A1(_19280_),
    .A2(net1842),
    .B1(_19555_),
    .Y(_05484_));
 sky130_fd_sc_hd__inv_1 _41857_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[17] ),
    .Y(_19556_));
 sky130_fd_sc_hd__o21ai_0 _41860_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[1] ),
    .A2(net1842),
    .B1(net2123),
    .Y(_19559_));
 sky130_fd_sc_hd__a21oi_1 _41861_ (.A1(_19556_),
    .A2(net1842),
    .B1(_19559_),
    .Y(_05485_));
 sky130_fd_sc_hd__o21ai_0 _41862_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[2] ),
    .A2(net1841),
    .B1(net2121),
    .Y(_19560_));
 sky130_fd_sc_hd__a21oi_1 _41863_ (.A1(_19318_),
    .A2(net1841),
    .B1(_19560_),
    .Y(_05486_));
 sky130_fd_sc_hd__o21ai_0 _41864_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[3] ),
    .A2(net1841),
    .B1(net2121),
    .Y(_19561_));
 sky130_fd_sc_hd__a21oi_1 _41865_ (.A1(_19298_),
    .A2(net1841),
    .B1(_19561_),
    .Y(_05487_));
 sky130_fd_sc_hd__o21ai_0 _41866_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[1] ),
    .A2(net1843),
    .B1(net2132),
    .Y(_19562_));
 sky130_fd_sc_hd__a21oi_1 _41867_ (.A1(_02707_),
    .A2(net1843),
    .B1(_19562_),
    .Y(_05488_));
 sky130_fd_sc_hd__o21ai_0 _41868_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[4] ),
    .A2(net1841),
    .B1(net2121),
    .Y(_19563_));
 sky130_fd_sc_hd__a21oi_1 _41869_ (.A1(_19310_),
    .A2(net1841),
    .B1(_19563_),
    .Y(_05489_));
 sky130_fd_sc_hd__o21ai_0 _41870_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[5] ),
    .A2(net1841),
    .B1(net2123),
    .Y(_19564_));
 sky130_fd_sc_hd__a21oi_1 _41871_ (.A1(_19317_),
    .A2(net1842),
    .B1(_19564_),
    .Y(_05490_));
 sky130_fd_sc_hd__o21ai_0 _41872_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[6] ),
    .A2(net1841),
    .B1(net2121),
    .Y(_19565_));
 sky130_fd_sc_hd__a21oi_1 _41873_ (.A1(_19329_),
    .A2(net1842),
    .B1(_19565_),
    .Y(_05491_));
 sky130_fd_sc_hd__o21ai_0 _41874_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[7] ),
    .A2(net1841),
    .B1(net2123),
    .Y(_19566_));
 sky130_fd_sc_hd__a21oi_1 _41875_ (.A1(_19341_),
    .A2(net1841),
    .B1(_19566_),
    .Y(_05492_));
 sky130_fd_sc_hd__o21ai_0 _41876_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[2] ),
    .A2(net1843),
    .B1(net2133),
    .Y(_19567_));
 sky130_fd_sc_hd__a21oi_1 _41877_ (.A1(_19186_),
    .A2(net1844),
    .B1(_19567_),
    .Y(_05493_));
 sky130_fd_sc_hd__nand2_1 _41878_ (.A(_19543_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[3] ),
    .Y(_19568_));
 sky130_fd_sc_hd__nand2_1 _41879_ (.A(net1844),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[3] ),
    .Y(_19569_));
 sky130_fd_sc_hd__nand3_1 _41880_ (.A(_19568_),
    .B(_19569_),
    .C(net2132),
    .Y(_05494_));
 sky130_fd_sc_hd__nand2_1 _41881_ (.A(_19543_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[4] ),
    .Y(_19570_));
 sky130_fd_sc_hd__nand2_1 _41882_ (.A(net1844),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[4] ),
    .Y(_19571_));
 sky130_fd_sc_hd__nand3_1 _41883_ (.A(_19570_),
    .B(_19571_),
    .C(net2133),
    .Y(_05495_));
 sky130_fd_sc_hd__nor2_1 _41884_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[5] ),
    .B(_19543_),
    .Y(_19572_));
 sky130_fd_sc_hd__o21ai_0 _41885_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[5] ),
    .A2(net1843),
    .B1(net2133),
    .Y(_19573_));
 sky130_fd_sc_hd__nor2_1 _41886_ (.A(_19572_),
    .B(_19573_),
    .Y(_05496_));
 sky130_fd_sc_hd__nand2_1 _41887_ (.A(_19543_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[6] ),
    .Y(_19574_));
 sky130_fd_sc_hd__nand2_1 _41888_ (.A(net1843),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[6] ),
    .Y(_19575_));
 sky130_fd_sc_hd__nand3_1 _41889_ (.A(_19574_),
    .B(_19575_),
    .C(net2133),
    .Y(_05497_));
 sky130_fd_sc_hd__nand2_1 _41890_ (.A(_19543_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[7] ),
    .Y(_19576_));
 sky130_fd_sc_hd__nand2_1 _41891_ (.A(net1844),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[7] ),
    .Y(_19577_));
 sky130_fd_sc_hd__nand3_1 _41892_ (.A(_19576_),
    .B(_19577_),
    .C(net2135),
    .Y(_05498_));
 sky130_fd_sc_hd__o21ai_0 _41893_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[0] ),
    .A2(net1843),
    .B1(net2133),
    .Y(_19578_));
 sky130_fd_sc_hd__a21oi_1 _41894_ (.A1(_19182_),
    .A2(net1844),
    .B1(_19578_),
    .Y(_05499_));
 sky130_fd_sc_hd__nor2_1 _41895_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[9] ),
    .B(_19543_),
    .Y(_19579_));
 sky130_fd_sc_hd__o21ai_0 _41896_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[1] ),
    .A2(net1843),
    .B1(net2133),
    .Y(_19580_));
 sky130_fd_sc_hd__nor2_1 _41897_ (.A(_19579_),
    .B(_19580_),
    .Y(_05500_));
 sky130_fd_sc_hd__nor2_1 _41898_ (.A(_19868_),
    .B(_19432_),
    .Y(_19581_));
 sky130_fd_sc_hd__inv_1 _41899_ (.A(_19581_),
    .Y(_19582_));
 sky130_fd_sc_hd__nor3_1 _41900_ (.A(net2987),
    .B(_19492_),
    .C(_19582_),
    .Y(_05501_));
 sky130_fd_sc_hd__nor2_1 _41901_ (.A(_19435_),
    .B(_19582_),
    .Y(_05502_));
 sky130_fd_sc_hd__nor2_1 _41902_ (.A(_18044_),
    .B(_19582_),
    .Y(_05503_));
 sky130_fd_sc_hd__inv_1 _41903_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[0] ),
    .Y(_19583_));
 sky130_fd_sc_hd__nand2_1 _41904_ (.A(_19072_),
    .B(\inst$top.soc.bus__adr[2] ),
    .Y(_19584_));
 sky130_fd_sc_hd__inv_1 _41905_ (.A(_19584_),
    .Y(_19585_));
 sky130_fd_sc_hd__nand2_1 _41906_ (.A(_19585_),
    .B(_19436_),
    .Y(_19586_));
 sky130_fd_sc_hd__nor2_1 _41907_ (.A(\inst$top.soc.uart_0._phy.tx.lower.fsm_state ),
    .B(_18138_),
    .Y(_19587_));
 sky130_fd_sc_hd__o22ai_1 _41908_ (.A1(_19109_),
    .A2(_17887_),
    .B1(_02706_),
    .B2(_18096_),
    .Y(_19588_));
 sky130_fd_sc_hd__o31ai_1 _41909_ (.A1(_19587_),
    .A2(_19588_),
    .A3(_19586_),
    .B1(net2132),
    .Y(_19589_));
 sky130_fd_sc_hd__a21oi_1 _41910_ (.A1(_19583_),
    .A2(_19586_),
    .B1(_19589_),
    .Y(_05504_));
 sky130_fd_sc_hd__nand2_1 _41911_ (.A(_19586_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[1] ),
    .Y(_19590_));
 sky130_fd_sc_hd__nor2_2 _41912_ (.A(_18096_),
    .B(_19584_),
    .Y(_19591_));
 sky130_fd_sc_hd__nand2_1 _41914_ (.A(_19591_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[1] ),
    .Y(_19593_));
 sky130_fd_sc_hd__a21oi_2 _41915_ (.A1(_19590_),
    .A2(_19593_),
    .B1(net2985),
    .Y(_05505_));
 sky130_fd_sc_hd__nand2_1 _41916_ (.A(_19586_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[2] ),
    .Y(_19594_));
 sky130_fd_sc_hd__nand2_1 _41917_ (.A(net799),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[2] ),
    .Y(_19595_));
 sky130_fd_sc_hd__a21oi_2 _41918_ (.A1(_19594_),
    .A2(_19595_),
    .B1(net2984),
    .Y(_05506_));
 sky130_fd_sc_hd__nand2_1 _41919_ (.A(_19586_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[3] ),
    .Y(_19596_));
 sky130_fd_sc_hd__nand2_1 _41920_ (.A(net799),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[3] ),
    .Y(_19597_));
 sky130_fd_sc_hd__a21oi_2 _41921_ (.A1(_19596_),
    .A2(_19597_),
    .B1(net2984),
    .Y(_05507_));
 sky130_fd_sc_hd__nand2_1 _41922_ (.A(_19586_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[4] ),
    .Y(_19598_));
 sky130_fd_sc_hd__nand2_1 _41923_ (.A(net799),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[4] ),
    .Y(_19599_));
 sky130_fd_sc_hd__a21oi_2 _41924_ (.A1(_19598_),
    .A2(_19599_),
    .B1(net2984),
    .Y(_05508_));
 sky130_fd_sc_hd__nand2_1 _41925_ (.A(_19586_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[5] ),
    .Y(_19600_));
 sky130_fd_sc_hd__nand2_1 _41926_ (.A(net799),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[5] ),
    .Y(_19601_));
 sky130_fd_sc_hd__a21oi_2 _41927_ (.A1(_19600_),
    .A2(_19601_),
    .B1(net2987),
    .Y(_05509_));
 sky130_fd_sc_hd__nand2_1 _41928_ (.A(_19586_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[6] ),
    .Y(_19602_));
 sky130_fd_sc_hd__nand2_1 _41929_ (.A(net799),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[6] ),
    .Y(_19603_));
 sky130_fd_sc_hd__a21oi_2 _41930_ (.A1(_19602_),
    .A2(_19603_),
    .B1(net2984),
    .Y(_05510_));
 sky130_fd_sc_hd__nand2_1 _41931_ (.A(_19586_),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[7] ),
    .Y(_19604_));
 sky130_fd_sc_hd__nand2_1 _41933_ (.A(net799),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[7] ),
    .Y(_19606_));
 sky130_fd_sc_hd__a21oi_2 _41934_ (.A1(_19604_),
    .A2(_19606_),
    .B1(net2984),
    .Y(_05511_));
 sky130_fd_sc_hd__nor2_1 _41935_ (.A(net2987),
    .B(_19586_),
    .Y(_05512_));
 sky130_fd_sc_hd__o21ai_0 _41938_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[0] ),
    .A2(net799),
    .B1(net2132),
    .Y(_19609_));
 sky130_fd_sc_hd__a21oi_2 _41939_ (.A1(_19182_),
    .A2(net799),
    .B1(_19609_),
    .Y(_05513_));
 sky130_fd_sc_hd__inv_1 _41940_ (.A(net798),
    .Y(_19610_));
 sky130_fd_sc_hd__inv_1 _41941_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[1] ),
    .Y(_19611_));
 sky130_fd_sc_hd__nor2_1 _41942_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[9] ),
    .B(_19610_),
    .Y(_19612_));
 sky130_fd_sc_hd__a211oi_2 _41943_ (.A1(_19610_),
    .A2(_19611_),
    .B1(net2984),
    .C1(_19612_),
    .Y(_05514_));
 sky130_fd_sc_hd__o21ai_0 _41944_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[2] ),
    .A2(net798),
    .B1(net2122),
    .Y(_19613_));
 sky130_fd_sc_hd__a21oi_2 _41945_ (.A1(_19180_),
    .A2(_19591_),
    .B1(_19613_),
    .Y(_05515_));
 sky130_fd_sc_hd__o21ai_0 _41946_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[3] ),
    .A2(net798),
    .B1(net2132),
    .Y(_19614_));
 sky130_fd_sc_hd__a21oi_2 _41947_ (.A1(_19223_),
    .A2(net798),
    .B1(_19614_),
    .Y(_05516_));
 sky130_fd_sc_hd__o21ai_0 _41948_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[4] ),
    .A2(net799),
    .B1(net2140),
    .Y(_19615_));
 sky130_fd_sc_hd__a21oi_2 _41949_ (.A1(_19221_),
    .A2(net799),
    .B1(_19615_),
    .Y(_05517_));
 sky130_fd_sc_hd__inv_1 _41950_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[5] ),
    .Y(_19616_));
 sky130_fd_sc_hd__nor2_1 _41951_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[13] ),
    .B(_19610_),
    .Y(_19617_));
 sky130_fd_sc_hd__a211oi_2 _41952_ (.A1(_19610_),
    .A2(_19616_),
    .B1(net2984),
    .C1(_19617_),
    .Y(_05518_));
 sky130_fd_sc_hd__o21ai_0 _41953_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[6] ),
    .A2(net798),
    .B1(net2124),
    .Y(_19618_));
 sky130_fd_sc_hd__a21oi_2 _41954_ (.A1(_19248_),
    .A2(net798),
    .B1(_19618_),
    .Y(_05519_));
 sky130_fd_sc_hd__o21ai_0 _41955_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[7] ),
    .A2(net798),
    .B1(net2124),
    .Y(_19619_));
 sky130_fd_sc_hd__a21oi_2 _41956_ (.A1(_19261_),
    .A2(net798),
    .B1(_19619_),
    .Y(_05520_));
 sky130_fd_sc_hd__nor2_1 _41957_ (.A(_17872_),
    .B(_19584_),
    .Y(_05521_));
 sky130_fd_sc_hd__o21ai_0 _41958_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[0] ),
    .A2(net796),
    .B1(net2122),
    .Y(_19620_));
 sky130_fd_sc_hd__a21oi_2 _41959_ (.A1(_19280_),
    .A2(net796),
    .B1(_19620_),
    .Y(_05522_));
 sky130_fd_sc_hd__o21ai_0 _41960_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[1] ),
    .A2(net797),
    .B1(net2123),
    .Y(_19621_));
 sky130_fd_sc_hd__a21oi_2 _41961_ (.A1(_19556_),
    .A2(net797),
    .B1(_19621_),
    .Y(_05523_));
 sky130_fd_sc_hd__o21ai_0 _41962_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[2] ),
    .A2(net796),
    .B1(net2121),
    .Y(_19622_));
 sky130_fd_sc_hd__a21oi_2 _41963_ (.A1(_19318_),
    .A2(net796),
    .B1(_19622_),
    .Y(_05524_));
 sky130_fd_sc_hd__o21ai_0 _41964_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[3] ),
    .A2(net796),
    .B1(net2121),
    .Y(_19623_));
 sky130_fd_sc_hd__a21oi_1 _41965_ (.A1(_19298_),
    .A2(net796),
    .B1(_19623_),
    .Y(_05525_));
 sky130_fd_sc_hd__o21ai_0 _41967_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[4] ),
    .A2(net796),
    .B1(net2123),
    .Y(_19625_));
 sky130_fd_sc_hd__a21oi_1 _41968_ (.A1(_19310_),
    .A2(net797),
    .B1(_19625_),
    .Y(_05526_));
 sky130_fd_sc_hd__o21ai_0 _41969_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[5] ),
    .A2(net796),
    .B1(net2123),
    .Y(_19626_));
 sky130_fd_sc_hd__a21oi_1 _41970_ (.A1(_19317_),
    .A2(net797),
    .B1(_19626_),
    .Y(_05527_));
 sky130_fd_sc_hd__o21ai_0 _41971_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[6] ),
    .A2(net796),
    .B1(net2124),
    .Y(_19627_));
 sky130_fd_sc_hd__a21oi_1 _41972_ (.A1(_19329_),
    .A2(net796),
    .B1(_19627_),
    .Y(_05528_));
 sky130_fd_sc_hd__o21ai_0 _41973_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[7] ),
    .A2(net797),
    .B1(net2123),
    .Y(_19628_));
 sky130_fd_sc_hd__a21oi_1 _41974_ (.A1(_19341_),
    .A2(net797),
    .B1(_19628_),
    .Y(_05529_));
 sky130_fd_sc_hd__nor3_1 _41975_ (.A(net2985),
    .B(_19504_),
    .C(_19584_),
    .Y(_05530_));
 sky130_fd_sc_hd__nand2_1 _41976_ (.A(_19516_),
    .B(\inst$top.soc.bus__adr[2] ),
    .Y(_19629_));
 sky130_fd_sc_hd__nor2_1 _41977_ (.A(_17932_),
    .B(_19629_),
    .Y(_19630_));
 sky130_fd_sc_hd__nor2_1 _41979_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.Config.enable.port__w_data ),
    .B(net824),
    .Y(_19632_));
 sky130_fd_sc_hd__a211oi_2 _41980_ (.A1(net824),
    .A2(net900),
    .B1(net2992),
    .C1(_19632_),
    .Y(_05531_));
 sky130_fd_sc_hd__nor2_1 _41981_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[1] ),
    .B(net823),
    .Y(_19633_));
 sky130_fd_sc_hd__a211oi_2 _41982_ (.A1(net823),
    .A2(net868),
    .B1(net2986),
    .C1(_19633_),
    .Y(_05532_));
 sky130_fd_sc_hd__nor2_1 _41983_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[2] ),
    .B(net823),
    .Y(_19634_));
 sky130_fd_sc_hd__a211oi_2 _41984_ (.A1(net823),
    .A2(_17954_),
    .B1(net2986),
    .C1(_19634_),
    .Y(_05533_));
 sky130_fd_sc_hd__nor2_1 _41986_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[3] ),
    .B(net823),
    .Y(_19636_));
 sky130_fd_sc_hd__a211oi_2 _41987_ (.A1(net824),
    .A2(_17960_),
    .B1(net2986),
    .C1(_19636_),
    .Y(_05534_));
 sky130_fd_sc_hd__nor2_1 _41988_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[4] ),
    .B(net823),
    .Y(_19637_));
 sky130_fd_sc_hd__a211oi_2 _41989_ (.A1(net824),
    .A2(net867),
    .B1(net2987),
    .C1(_19637_),
    .Y(_05535_));
 sky130_fd_sc_hd__nor2_1 _41990_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[5] ),
    .B(net823),
    .Y(_19638_));
 sky130_fd_sc_hd__a211oi_2 _41991_ (.A1(net823),
    .A2(_17972_),
    .B1(net2987),
    .C1(_19638_),
    .Y(_05536_));
 sky130_fd_sc_hd__nor2_1 _41992_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[6] ),
    .B(net823),
    .Y(_19639_));
 sky130_fd_sc_hd__a211oi_2 _41993_ (.A1(net823),
    .A2(_17977_),
    .B1(net2986),
    .C1(_19639_),
    .Y(_05537_));
 sky130_fd_sc_hd__nor2_1 _41994_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[7] ),
    .B(net824),
    .Y(_19640_));
 sky130_fd_sc_hd__a211oi_2 _41995_ (.A1(net824),
    .A2(_17982_),
    .B1(net2992),
    .C1(_19640_),
    .Y(_05538_));
 sky130_fd_sc_hd__nor2_1 _41996_ (.A(_19494_),
    .B(_19629_),
    .Y(_19641_));
 sky130_fd_sc_hd__nor2_1 _41998_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[0] ),
    .B(net822),
    .Y(_19643_));
 sky130_fd_sc_hd__a211oi_2 _41999_ (.A1(net822),
    .A2(net900),
    .B1(net2986),
    .C1(_19643_),
    .Y(_05539_));
 sky130_fd_sc_hd__nor2_1 _42000_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[1] ),
    .B(net822),
    .Y(_19644_));
 sky130_fd_sc_hd__a211oi_2 _42001_ (.A1(net822),
    .A2(net868),
    .B1(net2986),
    .C1(_19644_),
    .Y(_05540_));
 sky130_fd_sc_hd__nor2_1 _42002_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[2] ),
    .B(net821),
    .Y(_19645_));
 sky130_fd_sc_hd__a211oi_2 _42003_ (.A1(net822),
    .A2(_17954_),
    .B1(net2986),
    .C1(_19645_),
    .Y(_05541_));
 sky130_fd_sc_hd__nor2_1 _42004_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[3] ),
    .B(net821),
    .Y(_19646_));
 sky130_fd_sc_hd__a211oi_2 _42005_ (.A1(net822),
    .A2(_17960_),
    .B1(net2986),
    .C1(_19646_),
    .Y(_05542_));
 sky130_fd_sc_hd__nor2_1 _42006_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[4] ),
    .B(net821),
    .Y(_19647_));
 sky130_fd_sc_hd__a211oi_2 _42007_ (.A1(net821),
    .A2(net867),
    .B1(net2986),
    .C1(_19647_),
    .Y(_05543_));
 sky130_fd_sc_hd__nor2_1 _42009_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[5] ),
    .B(net821),
    .Y(_19649_));
 sky130_fd_sc_hd__a211oi_2 _42010_ (.A1(net821),
    .A2(_17972_),
    .B1(net2985),
    .C1(_19649_),
    .Y(_05544_));
 sky130_fd_sc_hd__nor2_1 _42011_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[6] ),
    .B(net821),
    .Y(_19650_));
 sky130_fd_sc_hd__a211oi_2 _42012_ (.A1(net821),
    .A2(_17977_),
    .B1(net2985),
    .C1(_19650_),
    .Y(_05545_));
 sky130_fd_sc_hd__nor2_1 _42013_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[7] ),
    .B(net821),
    .Y(_19651_));
 sky130_fd_sc_hd__a211oi_2 _42014_ (.A1(net821),
    .A2(_17982_),
    .B1(net2985),
    .C1(_19651_),
    .Y(_05546_));
 sky130_fd_sc_hd__nor2_1 _42015_ (.A(_19504_),
    .B(_19582_),
    .Y(_19652_));
 sky130_fd_sc_hd__o21ai_0 _42017_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[0] ),
    .A2(net795),
    .B1(net2122),
    .Y(_19654_));
 sky130_fd_sc_hd__a21oi_2 _42018_ (.A1(net900),
    .A2(net795),
    .B1(_19654_),
    .Y(_05547_));
 sky130_fd_sc_hd__o21ai_0 _42019_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[1] ),
    .A2(net795),
    .B1(net2124),
    .Y(_19655_));
 sky130_fd_sc_hd__a21oi_2 _42020_ (.A1(net868),
    .A2(net795),
    .B1(_19655_),
    .Y(_05548_));
 sky130_fd_sc_hd__o21ai_0 _42021_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[2] ),
    .A2(net794),
    .B1(net2121),
    .Y(_19656_));
 sky130_fd_sc_hd__a21oi_2 _42022_ (.A1(_17954_),
    .A2(net794),
    .B1(_19656_),
    .Y(_05549_));
 sky130_fd_sc_hd__o21ai_0 _42023_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[3] ),
    .A2(net794),
    .B1(net2121),
    .Y(_19657_));
 sky130_fd_sc_hd__a21oi_2 _42024_ (.A1(_17960_),
    .A2(net794),
    .B1(_19657_),
    .Y(_05550_));
 sky130_fd_sc_hd__o21ai_0 _42025_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[4] ),
    .A2(net794),
    .B1(net2121),
    .Y(_19658_));
 sky130_fd_sc_hd__a21oi_2 _42026_ (.A1(net867),
    .A2(net794),
    .B1(_19658_),
    .Y(_05551_));
 sky130_fd_sc_hd__nor2_1 _42027_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[5] ),
    .B(net794),
    .Y(_19659_));
 sky130_fd_sc_hd__a211oi_2 _42028_ (.A1(net795),
    .A2(_17972_),
    .B1(net2983),
    .C1(_19659_),
    .Y(_05552_));
 sky130_fd_sc_hd__o21ai_0 _42029_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[6] ),
    .A2(net794),
    .B1(net2121),
    .Y(_19660_));
 sky130_fd_sc_hd__a21oi_2 _42030_ (.A1(_17977_),
    .A2(net795),
    .B1(_19660_),
    .Y(_05553_));
 sky130_fd_sc_hd__nor2_1 _42031_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[7] ),
    .B(net794),
    .Y(_19661_));
 sky130_fd_sc_hd__a211oi_2 _42032_ (.A1(net794),
    .A2(_17982_),
    .B1(net2983),
    .C1(_19661_),
    .Y(_05554_));
 sky130_fd_sc_hd__a21oi_1 _42033_ (.A1(_09340_),
    .A2(net2566),
    .B1(\inst$top.soc.cpu.loadstore.dbus__cyc ),
    .Y(_19662_));
 sky130_fd_sc_hd__nor3_1 _42034_ (.A(net2949),
    .B(_09341_),
    .C(_19662_),
    .Y(_05555_));
 sky130_fd_sc_hd__nor2_1 _42035_ (.A(_17849_),
    .B(_17865_),
    .Y(_19663_));
 sky130_fd_sc_hd__nor2_1 _42036_ (.A(net2979),
    .B(\inst$top.soc.wb_to_csr.wb_bus__ack ),
    .Y(_19664_));
 sky130_fd_sc_hd__o21ai_0 _42037_ (.A1(\inst$top.soc.wb_to_csr.cycle[0] ),
    .A2(_17947_),
    .B1(_19664_),
    .Y(_19665_));
 sky130_fd_sc_hd__nor2_1 _42038_ (.A(_19663_),
    .B(_19665_),
    .Y(_05556_));
 sky130_fd_sc_hd__inv_1 _42039_ (.A(_19664_),
    .Y(_19666_));
 sky130_fd_sc_hd__a21oi_1 _42040_ (.A1(_19663_),
    .A2(\inst$top.soc.wb_to_csr.cycle[1] ),
    .B1(_19666_),
    .Y(_19667_));
 sky130_fd_sc_hd__o21a_1 _42041_ (.A1(\inst$top.soc.wb_to_csr.cycle[1] ),
    .A2(_19663_),
    .B1(_19667_),
    .X(_19668_));
 sky130_fd_sc_hd__nor2_1 _42043_ (.A(_17831_),
    .B(_17865_),
    .Y(_19669_));
 sky130_fd_sc_hd__inv_1 _42044_ (.A(_19669_),
    .Y(_19670_));
 sky130_fd_sc_hd__a21oi_1 _42046_ (.A1(net863),
    .A2(_17864_),
    .B1(_19666_),
    .Y(_05558_));
 sky130_fd_sc_hd__nand2_1 _42047_ (.A(_17863_),
    .B(\inst$top.soc.wb_to_csr.cycle[2] ),
    .Y(_19672_));
 sky130_fd_sc_hd__nor2_1 _42049_ (.A(_19666_),
    .B(_19672_),
    .Y(_05559_));
 sky130_fd_sc_hd__nand2_1 _42050_ (.A(_17863_),
    .B(_17852_),
    .Y(_19674_));
 sky130_fd_sc_hd__a22o_1 _42052_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[0] ),
    .B1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__r_en ),
    .B2(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[0] ),
    .X(_19676_));
 sky130_fd_sc_hd__a221oi_1 _42053_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__r_en ),
    .A2(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[0] ),
    .B1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__r_en ),
    .B2(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[0] ),
    .C1(_19676_),
    .Y(_19677_));
 sky130_fd_sc_hd__nand2_1 _42054_ (.A(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[0] ),
    .B(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__r_en ),
    .Y(_19678_));
 sky130_fd_sc_hd__nand2_1 _42055_ (.A(\inst$top.soc.soc_id.bridge.mux.r_shadow__2__r_en ),
    .B(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[1] ),
    .Y(_19679_));
 sky130_fd_sc_hd__nand2_1 _42056_ (.A(_19678_),
    .B(_19679_),
    .Y(_19680_));
 sky130_fd_sc_hd__inv_1 _42057_ (.A(_19680_),
    .Y(_19681_));
 sky130_fd_sc_hd__nand2_1 _42058_ (.A(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[6] ),
    .B(\inst$top.soc.soc_id.bridge.mux.r_shadow__3__r_en ),
    .Y(_19682_));
 sky130_fd_sc_hd__nand2_1 _42059_ (.A(_19681_),
    .B(_19682_),
    .Y(_19683_));
 sky130_fd_sc_hd__inv_1 _42060_ (.A(_19683_),
    .Y(_19684_));
 sky130_fd_sc_hd__inv_1 _42061_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__r_en ),
    .Y(_19685_));
 sky130_fd_sc_hd__nand2_1 _42062_ (.A(\inst$top.soc.soc_id.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[6] ),
    .Y(_19686_));
 sky130_fd_sc_hd__o21ai_0 _42063_ (.A1(_19685_),
    .A2(_19583_),
    .B1(_19686_),
    .Y(_19687_));
 sky130_fd_sc_hd__a221oi_1 _42064_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__r_en ),
    .A2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[0] ),
    .B1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__r_en ),
    .B2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[0] ),
    .C1(_19687_),
    .Y(_19688_));
 sky130_fd_sc_hd__a22o_1 _42065_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[0] ),
    .B1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__r_en ),
    .B2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[0] ),
    .X(_19689_));
 sky130_fd_sc_hd__a21oi_1 _42066_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[0] ),
    .B1(_19689_),
    .Y(_19690_));
 sky130_fd_sc_hd__nand4_1 _42067_ (.A(_19677_),
    .B(_19684_),
    .C(_19688_),
    .D(_19690_),
    .Y(_19691_));
 sky130_fd_sc_hd__o21ai_0 _42069_ (.A1(net897),
    .A2(_19691_),
    .B1(net2051),
    .Y(_19693_));
 sky130_fd_sc_hd__a21oi_1 _42070_ (.A1(_12700_),
    .A2(net897),
    .B1(_19693_),
    .Y(_05560_));
 sky130_fd_sc_hd__nand2_1 _42071_ (.A(_17863_),
    .B(_17857_),
    .Y(_19694_));
 sky130_fd_sc_hd__a22o_1 _42073_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[2] ),
    .B1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__r_en ),
    .B2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[2] ),
    .X(_19696_));
 sky130_fd_sc_hd__a221oi_1 _42074_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[2] ),
    .B1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__r_en ),
    .B2(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[2] ),
    .C1(_19696_),
    .Y(_19697_));
 sky130_fd_sc_hd__nand2_1 _42075_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[2] ),
    .Y(_19698_));
 sky130_fd_sc_hd__nand2_1 _42076_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__r_en ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[2] ),
    .Y(_19699_));
 sky130_fd_sc_hd__nand2_1 _42077_ (.A(_19698_),
    .B(_19699_),
    .Y(_19700_));
 sky130_fd_sc_hd__nand2_1 _42078_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[2] ),
    .Y(_19701_));
 sky130_fd_sc_hd__nand2_1 _42079_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[2] ),
    .Y(_19702_));
 sky130_fd_sc_hd__nand2_1 _42080_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[2] ),
    .Y(_19703_));
 sky130_fd_sc_hd__nand3_1 _42081_ (.A(_19701_),
    .B(_19702_),
    .C(_19703_),
    .Y(_19704_));
 sky130_fd_sc_hd__a211oi_1 _42082_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[2] ),
    .B1(_19700_),
    .C1(_19704_),
    .Y(_19705_));
 sky130_fd_sc_hd__nand3_1 _42083_ (.A(_19697_),
    .B(_19684_),
    .C(_19705_),
    .Y(_19706_));
 sky130_fd_sc_hd__o21ai_0 _42084_ (.A1(net894),
    .A2(_19706_),
    .B1(net2055),
    .Y(_19707_));
 sky130_fd_sc_hd__a21oi_1 _42085_ (.A1(_12718_),
    .A2(net894),
    .B1(_19707_),
    .Y(_05561_));
 sky130_fd_sc_hd__a22o_1 _42086_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[3] ),
    .B1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__r_en ),
    .B2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[3] ),
    .X(_19708_));
 sky130_fd_sc_hd__a221oi_2 _42087_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[3] ),
    .B1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__r_en ),
    .B2(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[3] ),
    .C1(_19708_),
    .Y(_19709_));
 sky130_fd_sc_hd__a221oi_1 _42088_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[3] ),
    .B1(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[1] ),
    .B2(\inst$top.soc.soc_id.bridge.mux.r_shadow__3__r_en ),
    .C1(_19680_),
    .Y(_19710_));
 sky130_fd_sc_hd__nand2_1 _42089_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[3] ),
    .Y(_19711_));
 sky130_fd_sc_hd__nand2_1 _42090_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[3] ),
    .Y(_19712_));
 sky130_fd_sc_hd__nand2_1 _42091_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[3] ),
    .Y(_19713_));
 sky130_fd_sc_hd__nand3_1 _42092_ (.A(_19711_),
    .B(_19712_),
    .C(_19713_),
    .Y(_19714_));
 sky130_fd_sc_hd__a221oi_1 _42093_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__r_en ),
    .A2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[3] ),
    .B1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__r_en ),
    .B2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[3] ),
    .C1(_19714_),
    .Y(_19715_));
 sky130_fd_sc_hd__nand3_1 _42094_ (.A(_19709_),
    .B(_19710_),
    .C(_19715_),
    .Y(_19716_));
 sky130_fd_sc_hd__o21ai_0 _42095_ (.A1(net894),
    .A2(_19716_),
    .B1(net2054),
    .Y(_19717_));
 sky130_fd_sc_hd__a21oi_1 _42096_ (.A1(_12729_),
    .A2(net894),
    .B1(_19717_),
    .Y(_05562_));
 sky130_fd_sc_hd__a22o_1 _42097_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[4] ),
    .B1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__r_en ),
    .B2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[4] ),
    .X(_19718_));
 sky130_fd_sc_hd__a221oi_1 _42098_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[4] ),
    .B1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__r_en ),
    .B2(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[4] ),
    .C1(_19718_),
    .Y(_19719_));
 sky130_fd_sc_hd__a22o_1 _42099_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[4] ),
    .B1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__r_en ),
    .B2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[4] ),
    .X(_19720_));
 sky130_fd_sc_hd__a221oi_1 _42100_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__r_en ),
    .A2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[4] ),
    .B1(\inst$top.soc.soc_id.bridge.mux.r_shadow__1__r_en ),
    .B2(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[1] ),
    .C1(_19720_),
    .Y(_19721_));
 sky130_fd_sc_hd__nand2_1 _42101_ (.A(_19682_),
    .B(_19679_),
    .Y(_19722_));
 sky130_fd_sc_hd__a22o_1 _42102_ (.A1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__r_en ),
    .A2(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[4] ),
    .B1(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__r_en ),
    .B2(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[4] ),
    .X(_19723_));
 sky130_fd_sc_hd__a211oi_1 _42103_ (.A1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[4] ),
    .B1(_19722_),
    .C1(_19723_),
    .Y(_19724_));
 sky130_fd_sc_hd__nand3_1 _42104_ (.A(_19719_),
    .B(_19721_),
    .C(_19724_),
    .Y(_19725_));
 sky130_fd_sc_hd__o21ai_0 _42105_ (.A1(net894),
    .A2(_19725_),
    .B1(net2056),
    .Y(_19726_));
 sky130_fd_sc_hd__a21oi_1 _42106_ (.A1(_12736_),
    .A2(net895),
    .B1(_19726_),
    .Y(_05563_));
 sky130_fd_sc_hd__nand2_1 _42107_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[5] ),
    .Y(_19727_));
 sky130_fd_sc_hd__nand2_1 _42108_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[5] ),
    .Y(_19728_));
 sky130_fd_sc_hd__nand2_1 _42109_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[5] ),
    .Y(_19729_));
 sky130_fd_sc_hd__nand2_1 _42110_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[5] ),
    .Y(_19730_));
 sky130_fd_sc_hd__nand4_1 _42111_ (.A(_19727_),
    .B(_19728_),
    .C(_19729_),
    .D(_19730_),
    .Y(_19731_));
 sky130_fd_sc_hd__nand2_1 _42112_ (.A(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[5] ),
    .Y(_19732_));
 sky130_fd_sc_hd__nand2_1 _42113_ (.A(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[5] ),
    .Y(_19733_));
 sky130_fd_sc_hd__nand2_1 _42114_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[5] ),
    .Y(_19734_));
 sky130_fd_sc_hd__nand3_1 _42115_ (.A(_19732_),
    .B(_19733_),
    .C(_19734_),
    .Y(_19735_));
 sky130_fd_sc_hd__a221o_1 _42116_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__r_en ),
    .A2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[5] ),
    .B1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__r_en ),
    .B2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[5] ),
    .C1(_19722_),
    .X(_19736_));
 sky130_fd_sc_hd__a2111oi_1 _42117_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[5] ),
    .B1(_19731_),
    .C1(_19735_),
    .D1(_19736_),
    .Y(_19737_));
 sky130_fd_sc_hd__inv_1 _42118_ (.A(net1634),
    .Y(_19738_));
 sky130_fd_sc_hd__o21ai_0 _42119_ (.A1(net894),
    .A2(_19738_),
    .B1(net2057),
    .Y(_19739_));
 sky130_fd_sc_hd__a21oi_1 _42120_ (.A1(_12743_),
    .A2(net895),
    .B1(_19739_),
    .Y(_05564_));
 sky130_fd_sc_hd__nand2_1 _42121_ (.A(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[6] ),
    .Y(_19740_));
 sky130_fd_sc_hd__nand2_1 _42122_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[6] ),
    .Y(_19741_));
 sky130_fd_sc_hd__nand2_1 _42123_ (.A(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[6] ),
    .Y(_19742_));
 sky130_fd_sc_hd__nand2_1 _42124_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[6] ),
    .Y(_19743_));
 sky130_fd_sc_hd__nand4_1 _42125_ (.A(_19740_),
    .B(_19741_),
    .C(_19742_),
    .D(_19743_),
    .Y(_19744_));
 sky130_fd_sc_hd__nand2_1 _42126_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__r_en ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[6] ),
    .Y(_19745_));
 sky130_fd_sc_hd__nand2_1 _42127_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[6] ),
    .Y(_19746_));
 sky130_fd_sc_hd__nand2_1 _42128_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[6] ),
    .Y(_19747_));
 sky130_fd_sc_hd__nand2_1 _42129_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[6] ),
    .Y(_19748_));
 sky130_fd_sc_hd__nand4_1 _42130_ (.A(_19745_),
    .B(_19746_),
    .C(_19747_),
    .D(_19748_),
    .Y(_19749_));
 sky130_fd_sc_hd__nor2_1 _42131_ (.A(_19744_),
    .B(_19749_),
    .Y(_19750_));
 sky130_fd_sc_hd__nand2_1 _42132_ (.A(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[1] ),
    .B(\inst$top.soc.soc_id.bridge.mux.r_shadow__3__r_en ),
    .Y(_19751_));
 sky130_fd_sc_hd__nand2_1 _42133_ (.A(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[0] ),
    .B(\inst$top.soc.soc_id.bridge.mux.r_shadow__2__r_en ),
    .Y(_19752_));
 sky130_fd_sc_hd__nand2_1 _42134_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[6] ),
    .Y(_19753_));
 sky130_fd_sc_hd__nand2_1 _42135_ (.A(_19686_),
    .B(_19753_),
    .Y(_19754_));
 sky130_fd_sc_hd__a221oi_1 _42136_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[6] ),
    .B1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__r_en ),
    .B2(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[6] ),
    .C1(_19754_),
    .Y(_19755_));
 sky130_fd_sc_hd__nand4_1 _42137_ (.A(_19750_),
    .B(_19751_),
    .C(_19752_),
    .D(_19755_),
    .Y(_19756_));
 sky130_fd_sc_hd__o21ai_0 _42138_ (.A1(net894),
    .A2(_19756_),
    .B1(net2054),
    .Y(_19757_));
 sky130_fd_sc_hd__a21oi_1 _42139_ (.A1(_12750_),
    .A2(net894),
    .B1(_19757_),
    .Y(_05565_));
 sky130_fd_sc_hd__nand2_1 _42140_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[7] ),
    .Y(_19758_));
 sky130_fd_sc_hd__nand2_1 _42141_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[7] ),
    .Y(_19759_));
 sky130_fd_sc_hd__nand2_1 _42142_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[7] ),
    .Y(_19760_));
 sky130_fd_sc_hd__nand3_1 _42143_ (.A(_19758_),
    .B(_19759_),
    .C(_19760_),
    .Y(_19761_));
 sky130_fd_sc_hd__nand2_1 _42144_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[7] ),
    .Y(_19762_));
 sky130_fd_sc_hd__nand2_1 _42145_ (.A(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[6] ),
    .B(\inst$top.soc.soc_id.bridge.mux.r_shadow__2__r_en ),
    .Y(_19763_));
 sky130_fd_sc_hd__nand2_1 _42146_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__r_en ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[7] ),
    .Y(_19764_));
 sky130_fd_sc_hd__nand3_1 _42147_ (.A(_19762_),
    .B(_19763_),
    .C(_19764_),
    .Y(_19765_));
 sky130_fd_sc_hd__nand2_1 _42148_ (.A(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[7] ),
    .Y(_19766_));
 sky130_fd_sc_hd__nand2_1 _42149_ (.A(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[0] ),
    .B(\inst$top.soc.soc_id.bridge.mux.r_shadow__3__r_en ),
    .Y(_19767_));
 sky130_fd_sc_hd__nand3_1 _42150_ (.A(_19742_),
    .B(_19766_),
    .C(_19767_),
    .Y(_19768_));
 sky130_fd_sc_hd__nand2_1 _42151_ (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[7] ),
    .Y(_19769_));
 sky130_fd_sc_hd__nand2_1 _42152_ (.A(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[7] ),
    .Y(_19770_));
 sky130_fd_sc_hd__nand2_1 _42153_ (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[7] ),
    .Y(_19771_));
 sky130_fd_sc_hd__nand2_1 _42154_ (.A(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[7] ),
    .Y(_19772_));
 sky130_fd_sc_hd__nand4_1 _42155_ (.A(_19769_),
    .B(_19770_),
    .C(_19771_),
    .D(_19772_),
    .Y(_19773_));
 sky130_fd_sc_hd__nor4_1 _42156_ (.A(_19761_),
    .B(_19765_),
    .C(_19768_),
    .D(_19773_),
    .Y(_19774_));
 sky130_fd_sc_hd__inv_1 _42157_ (.A(_19774_),
    .Y(_19775_));
 sky130_fd_sc_hd__o21ai_0 _42158_ (.A1(net894),
    .A2(_19775_),
    .B1(net2054),
    .Y(_19776_));
 sky130_fd_sc_hd__a21oi_1 _42159_ (.A1(_12758_),
    .A2(net894),
    .B1(_19776_),
    .Y(_05566_));
 sky130_fd_sc_hd__nor2_1 _42160_ (.A(_19670_),
    .B(_19691_),
    .Y(_19777_));
 sky130_fd_sc_hd__a211oi_1 _42161_ (.A1(_19670_),
    .A2(_12765_),
    .B1(net2979),
    .C1(_19777_),
    .Y(_05567_));
 sky130_fd_sc_hd__nand2_1 _42162_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[1] ),
    .Y(_19778_));
 sky130_fd_sc_hd__nand2_1 _42163_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[1] ),
    .Y(_19779_));
 sky130_fd_sc_hd__nand2_1 _42164_ (.A(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__r_en ),
    .B(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[1] ),
    .Y(_19780_));
 sky130_fd_sc_hd__nand3_1 _42165_ (.A(_19778_),
    .B(_19779_),
    .C(_19780_),
    .Y(_19781_));
 sky130_fd_sc_hd__a22o_1 _42166_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__r_en ),
    .A2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[1] ),
    .B1(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__r_en ),
    .B2(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[1] ),
    .X(_19782_));
 sky130_fd_sc_hd__a211oi_1 _42167_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[1] ),
    .B1(_19781_),
    .C1(_19782_),
    .Y(_19783_));
 sky130_fd_sc_hd__a22o_1 _42168_ (.A1(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[1] ),
    .B1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__r_en ),
    .B2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[1] ),
    .X(_19784_));
 sky130_fd_sc_hd__a221oi_1 _42169_ (.A1(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__r_en ),
    .A2(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[1] ),
    .B1(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__r_en ),
    .B2(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[1] ),
    .C1(_19784_),
    .Y(_19785_));
 sky130_fd_sc_hd__nand2_1 _42170_ (.A(_19751_),
    .B(_19752_),
    .Y(_19786_));
 sky130_fd_sc_hd__a21oi_1 _42171_ (.A1(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__r_en ),
    .A2(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[1] ),
    .B1(_19786_),
    .Y(_19787_));
 sky130_fd_sc_hd__nand3_1 _42172_ (.A(_19783_),
    .B(_19785_),
    .C(_19787_),
    .Y(_19788_));
 sky130_fd_sc_hd__nor2_1 _42173_ (.A(net863),
    .B(_19788_),
    .Y(_19789_));
 sky130_fd_sc_hd__a211oi_1 _42174_ (.A1(_12772_),
    .A2(net863),
    .B1(net2979),
    .C1(_19789_),
    .Y(_05568_));
 sky130_fd_sc_hd__nor2_1 _42175_ (.A(net863),
    .B(_19706_),
    .Y(_19790_));
 sky130_fd_sc_hd__a211oi_1 _42176_ (.A1(net863),
    .A2(_12780_),
    .B1(net2979),
    .C1(_19790_),
    .Y(_05569_));
 sky130_fd_sc_hd__nor2_1 _42177_ (.A(net863),
    .B(_19716_),
    .Y(_19791_));
 sky130_fd_sc_hd__a211oi_1 _42178_ (.A1(_12788_),
    .A2(net863),
    .B1(net2979),
    .C1(_19791_),
    .Y(_05570_));
 sky130_fd_sc_hd__o21ai_0 _42179_ (.A1(net896),
    .A2(_19788_),
    .B1(net2051),
    .Y(_19792_));
 sky130_fd_sc_hd__a21oi_1 _42180_ (.A1(_12797_),
    .A2(net896),
    .B1(_19792_),
    .Y(_05571_));
 sky130_fd_sc_hd__nor2_1 _42181_ (.A(net863),
    .B(_19725_),
    .Y(_19793_));
 sky130_fd_sc_hd__a211oi_1 _42182_ (.A1(_19670_),
    .A2(_12804_),
    .B1(net2979),
    .C1(_19793_),
    .Y(_05572_));
 sky130_fd_sc_hd__o21ai_0 _42183_ (.A1(\inst$top.soc.wb_to_csr.wb_bus__dat_r[21] ),
    .A2(_19669_),
    .B1(net2119),
    .Y(_19794_));
 sky130_fd_sc_hd__a21oi_1 _42184_ (.A1(net1634),
    .A2(_19669_),
    .B1(_19794_),
    .Y(_05573_));
 sky130_fd_sc_hd__nor2_1 _42185_ (.A(_19756_),
    .B(net863),
    .Y(_19795_));
 sky130_fd_sc_hd__a211oi_1 _42186_ (.A1(net863),
    .A2(_12818_),
    .B1(net2979),
    .C1(_19795_),
    .Y(_05574_));
 sky130_fd_sc_hd__o21ai_0 _42187_ (.A1(\inst$top.soc.wb_to_csr.wb_bus__dat_r[23] ),
    .A2(_19669_),
    .B1(net2119),
    .Y(_19796_));
 sky130_fd_sc_hd__a21oi_1 _42188_ (.A1(_19669_),
    .A2(_19774_),
    .B1(_19796_),
    .Y(_05575_));
 sky130_fd_sc_hd__o21ai_0 _42190_ (.A1(net898),
    .A2(_19691_),
    .B1(net2052),
    .Y(_19798_));
 sky130_fd_sc_hd__a21oi_1 _42191_ (.A1(_12833_),
    .A2(net898),
    .B1(_19798_),
    .Y(_05576_));
 sky130_fd_sc_hd__o21ai_0 _42192_ (.A1(net898),
    .A2(_19788_),
    .B1(net2052),
    .Y(_19799_));
 sky130_fd_sc_hd__a21oi_1 _42193_ (.A1(_12840_),
    .A2(net899),
    .B1(_19799_),
    .Y(_05577_));
 sky130_fd_sc_hd__o21ai_0 _42194_ (.A1(net898),
    .A2(_19706_),
    .B1(net2052),
    .Y(_19800_));
 sky130_fd_sc_hd__a21oi_1 _42195_ (.A1(_12847_),
    .A2(net898),
    .B1(_19800_),
    .Y(_05578_));
 sky130_fd_sc_hd__o21ai_0 _42196_ (.A1(net898),
    .A2(_19716_),
    .B1(net2051),
    .Y(_19801_));
 sky130_fd_sc_hd__a21oi_1 _42197_ (.A1(_12855_),
    .A2(net898),
    .B1(_19801_),
    .Y(_05579_));
 sky130_fd_sc_hd__o21ai_0 _42198_ (.A1(net898),
    .A2(_19725_),
    .B1(net2053),
    .Y(_19802_));
 sky130_fd_sc_hd__a21oi_1 _42199_ (.A1(_12863_),
    .A2(net898),
    .B1(_19802_),
    .Y(_05580_));
 sky130_fd_sc_hd__o21ai_0 _42200_ (.A1(net898),
    .A2(_19738_),
    .B1(net2056),
    .Y(_19803_));
 sky130_fd_sc_hd__a21oi_1 _42201_ (.A1(_12870_),
    .A2(net899),
    .B1(_19803_),
    .Y(_05581_));
 sky130_fd_sc_hd__o21ai_0 _42202_ (.A1(net896),
    .A2(_19706_),
    .B1(net2053),
    .Y(_19804_));
 sky130_fd_sc_hd__a21oi_1 _42203_ (.A1(_12877_),
    .A2(net896),
    .B1(_19804_),
    .Y(_05582_));
 sky130_fd_sc_hd__o21ai_0 _42204_ (.A1(net899),
    .A2(_19756_),
    .B1(net2051),
    .Y(_19805_));
 sky130_fd_sc_hd__a21oi_1 _42205_ (.A1(_12884_),
    .A2(net899),
    .B1(_19805_),
    .Y(_05583_));
 sky130_fd_sc_hd__o21ai_0 _42206_ (.A1(net899),
    .A2(_19775_),
    .B1(net2056),
    .Y(_19806_));
 sky130_fd_sc_hd__a21oi_1 _42207_ (.A1(_12891_),
    .A2(net899),
    .B1(_19806_),
    .Y(_05584_));
 sky130_fd_sc_hd__o21ai_0 _42208_ (.A1(net896),
    .A2(_19716_),
    .B1(net2053),
    .Y(_19807_));
 sky130_fd_sc_hd__a21oi_1 _42209_ (.A1(_12898_),
    .A2(net896),
    .B1(_19807_),
    .Y(_05585_));
 sky130_fd_sc_hd__o21ai_0 _42210_ (.A1(net896),
    .A2(_19725_),
    .B1(net2051),
    .Y(_19808_));
 sky130_fd_sc_hd__a21oi_1 _42211_ (.A1(_12906_),
    .A2(net896),
    .B1(_19808_),
    .Y(_05586_));
 sky130_fd_sc_hd__o21ai_0 _42212_ (.A1(net897),
    .A2(_19738_),
    .B1(net2056),
    .Y(_19809_));
 sky130_fd_sc_hd__a21oi_1 _42213_ (.A1(_12913_),
    .A2(net897),
    .B1(_19809_),
    .Y(_05587_));
 sky130_fd_sc_hd__o21ai_0 _42214_ (.A1(net896),
    .A2(_19756_),
    .B1(net2053),
    .Y(_19810_));
 sky130_fd_sc_hd__a21oi_1 _42215_ (.A1(_12920_),
    .A2(net896),
    .B1(_19810_),
    .Y(_05588_));
 sky130_fd_sc_hd__o21ai_0 _42216_ (.A1(net897),
    .A2(_19775_),
    .B1(net2054),
    .Y(_19811_));
 sky130_fd_sc_hd__a21oi_1 _42217_ (.A1(_12927_),
    .A2(net897),
    .B1(_19811_),
    .Y(_05589_));
 sky130_fd_sc_hd__o21ai_0 _42218_ (.A1(net895),
    .A2(_19691_),
    .B1(net2056),
    .Y(_19812_));
 sky130_fd_sc_hd__a21oi_1 _42219_ (.A1(_12934_),
    .A2(net895),
    .B1(_19812_),
    .Y(_05590_));
 sky130_fd_sc_hd__o21ai_0 _42220_ (.A1(net895),
    .A2(_19788_),
    .B1(net2056),
    .Y(_19813_));
 sky130_fd_sc_hd__a21oi_1 _42221_ (.A1(_12941_),
    .A2(net895),
    .B1(_19813_),
    .Y(_05591_));
 sky130_fd_sc_hd__nand2_1 _42222_ (.A(_18019_),
    .B(_02888_),
    .Y(_19814_));
 sky130_fd_sc_hd__o21ai_4 _42223_ (.A1(_02889_),
    .A2(_02888_),
    .B1(_19814_),
    .Y(net556));
 sky130_fd_sc_hd__inv_2 _42224_ (.A(net1632),
    .Y(net572));
 sky130_fd_sc_hd__inv_2 _42225_ (.A(net2575),
    .Y(net576));
 sky130_fd_sc_hd__inv_2 _42226_ (.A(net2573),
    .Y(net577));
 sky130_fd_sc_hd__inv_2 _42227_ (.A(net2571),
    .Y(net578));
 sky130_fd_sc_hd__inv_2 _42228_ (.A(net2569),
    .Y(net579));
 sky130_fd_sc_hd__nand2_1 _42229_ (.A(_18021_),
    .B(_02885_),
    .Y(_19815_));
 sky130_fd_sc_hd__o21ai_4 _42230_ (.A1(_02886_),
    .A2(_02885_),
    .B1(_19815_),
    .Y(net557));
 sky130_fd_sc_hd__inv_2 _42231_ (.A(net1631),
    .Y(net573));
 sky130_fd_sc_hd__nand2_1 _42232_ (.A(_17796_),
    .B(_02872_),
    .Y(_19816_));
 sky130_fd_sc_hd__o21ai_4 _42233_ (.A1(_02873_),
    .A2(_02872_),
    .B1(_19816_),
    .Y(net564));
 sky130_fd_sc_hd__inv_2 _42234_ (.A(net1628),
    .Y(net580));
 sky130_fd_sc_hd__nand2_1 _42235_ (.A(_17801_),
    .B(_02894_),
    .Y(_19817_));
 sky130_fd_sc_hd__o21ai_4 _42236_ (.A1(_02895_),
    .A2(_02894_),
    .B1(_19817_),
    .Y(net565));
 sky130_fd_sc_hd__inv_2 _42237_ (.A(net1625),
    .Y(net581));
 sky130_fd_sc_hd__nand2_1 _42238_ (.A(_17805_),
    .B(_02869_),
    .Y(_19818_));
 sky130_fd_sc_hd__o21ai_4 _42239_ (.A1(_02870_),
    .A2(_02869_),
    .B1(_19818_),
    .Y(net550));
 sky130_fd_sc_hd__inv_2 _42240_ (.A(net1622),
    .Y(net566));
 sky130_fd_sc_hd__nand2_1 _42241_ (.A(_17810_),
    .B(_02897_),
    .Y(_19819_));
 sky130_fd_sc_hd__o21ai_4 _42242_ (.A1(_02898_),
    .A2(_02897_),
    .B1(_19819_),
    .Y(net551));
 sky130_fd_sc_hd__inv_2 _42243_ (.A(net1619),
    .Y(net567));
 sky130_fd_sc_hd__nand2_1 _42244_ (.A(_17814_),
    .B(_02909_),
    .Y(_19820_));
 sky130_fd_sc_hd__o21ai_4 _42245_ (.A1(_02910_),
    .A2(_02909_),
    .B1(_19820_),
    .Y(net552));
 sky130_fd_sc_hd__inv_2 _42246_ (.A(net1615),
    .Y(net568));
 sky130_fd_sc_hd__nand2_1 _42247_ (.A(_17818_),
    .B(_02906_),
    .Y(_19821_));
 sky130_fd_sc_hd__o21ai_4 _42248_ (.A1(_02907_),
    .A2(_02906_),
    .B1(_19821_),
    .Y(net553));
 sky130_fd_sc_hd__inv_2 _42249_ (.A(net1611),
    .Y(net569));
 sky130_fd_sc_hd__nand2_1 _42250_ (.A(_18025_),
    .B(_02891_),
    .Y(_19822_));
 sky130_fd_sc_hd__o21ai_4 _42251_ (.A1(_02892_),
    .A2(_02891_),
    .B1(_19822_),
    .Y(net558));
 sky130_fd_sc_hd__inv_2 _42252_ (.A(net1610),
    .Y(net574));
 sky130_fd_sc_hd__nand2_1 _42253_ (.A(_17822_),
    .B(_02903_),
    .Y(_19823_));
 sky130_fd_sc_hd__o21ai_4 _42254_ (.A1(_02904_),
    .A2(_02903_),
    .B1(_19823_),
    .Y(net554));
 sky130_fd_sc_hd__inv_2 _42255_ (.A(net1606),
    .Y(net570));
 sky130_fd_sc_hd__nand2_1 _42256_ (.A(_17827_),
    .B(_02900_),
    .Y(_19824_));
 sky130_fd_sc_hd__o21ai_4 _42257_ (.A1(_02901_),
    .A2(_02900_),
    .B1(_19824_),
    .Y(net555));
 sky130_fd_sc_hd__inv_2 _42258_ (.A(net1602),
    .Y(net571));
 sky130_fd_sc_hd__nand2_1 _42259_ (.A(_18029_),
    .B(_02875_),
    .Y(_19825_));
 sky130_fd_sc_hd__o21ai_4 _42260_ (.A1(_02876_),
    .A2(_02875_),
    .B1(_19825_),
    .Y(net559));
 sky130_fd_sc_hd__inv_2 _42261_ (.A(net1601),
    .Y(net575));
 sky130_fd_sc_hd__inv_2 _42262_ (.A(net2577),
    .Y(net589));
 sky130_fd_sc_hd__inv_2 _42263_ (.A(net544),
    .Y(\inst$top.i$88 ));
 sky130_fd_sc_hd__nor2_4 _42264_ (.A(_02872_),
    .B(_17796_),
    .Y(net599));
 sky130_fd_sc_hd__nor2_4 _42265_ (.A(_02894_),
    .B(_17801_),
    .Y(net600));
 sky130_fd_sc_hd__nor2_4 _42266_ (.A(_02869_),
    .B(_17805_),
    .Y(net583));
 sky130_fd_sc_hd__nor2_4 _42267_ (.A(_02897_),
    .B(_17810_),
    .Y(net584));
 sky130_fd_sc_hd__nor2_4 _42268_ (.A(_02909_),
    .B(_17814_),
    .Y(net585));
 sky130_fd_sc_hd__nor2_1 _42269_ (.A(_02906_),
    .B(_17818_),
    .Y(net586));
 sky130_fd_sc_hd__nor2_1 _42270_ (.A(_02903_),
    .B(_17822_),
    .Y(net587));
 sky130_fd_sc_hd__nor2_4 _42271_ (.A(_02900_),
    .B(_17827_),
    .Y(net588));
 sky130_fd_sc_hd__nor2_4 _42272_ (.A(_02888_),
    .B(_18019_),
    .Y(net590));
 sky130_fd_sc_hd__nor2_4 _42273_ (.A(_02885_),
    .B(_18021_),
    .Y(net591));
 sky130_fd_sc_hd__nor2_4 _42274_ (.A(_02891_),
    .B(_18025_),
    .Y(net592));
 sky130_fd_sc_hd__nor2_4 _42275_ (.A(_02875_),
    .B(_18029_),
    .Y(net593));
 sky130_fd_sc_hd__fa_1 _42276_ (.A(_00162_),
    .B(net1698),
    .CIN(net1706),
    .COUT(_00165_),
    .SUM(_00166_));
 sky130_fd_sc_hd__fa_1 _42277_ (.A(_00169_),
    .B(net1385),
    .CIN(net1706),
    .COUT(_00170_),
    .SUM(_00171_));
 sky130_fd_sc_hd__fa_1 _42278_ (.A(_00172_),
    .B(_00173_),
    .CIN(_00174_),
    .COUT(_20825_),
    .SUM(_20826_));
 sky130_fd_sc_hd__fa_1 _42279_ (.A(_00175_),
    .B(_00176_),
    .CIN(_00177_),
    .COUT(_00178_),
    .SUM(_00179_));
 sky130_fd_sc_hd__fa_1 _42280_ (.A(_00180_),
    .B(_20827_),
    .CIN(_20826_),
    .COUT(_20828_),
    .SUM(_20829_));
 sky130_fd_sc_hd__fa_1 _42281_ (.A(_00181_),
    .B(_00182_),
    .CIN(_00183_),
    .COUT(_20827_),
    .SUM(_20830_));
 sky130_fd_sc_hd__fa_1 _42282_ (.A(_00184_),
    .B(_00185_),
    .CIN(_00186_),
    .COUT(_20831_),
    .SUM(_20832_));
 sky130_fd_sc_hd__fa_1 _42283_ (.A(_20831_),
    .B(_20833_),
    .CIN(_20829_),
    .COUT(_00187_),
    .SUM(_00188_));
 sky130_fd_sc_hd__fa_1 _42284_ (.A(_20832_),
    .B(_00189_),
    .CIN(_20830_),
    .COUT(_20833_),
    .SUM(_20834_));
 sky130_fd_sc_hd__fa_1 _42285_ (.A(_00190_),
    .B(_00191_),
    .CIN(_00192_),
    .COUT(_20835_),
    .SUM(_00193_));
 sky130_fd_sc_hd__fa_1 _42286_ (.A(_00194_),
    .B(_00195_),
    .CIN(_00196_),
    .COUT(_20836_),
    .SUM(_00197_));
 sky130_fd_sc_hd__fa_1 _42287_ (.A(_20835_),
    .B(_00198_),
    .CIN(_20834_),
    .COUT(_00199_),
    .SUM(_00200_));
 sky130_fd_sc_hd__fa_1 _42288_ (.A(_20836_),
    .B(_00201_),
    .CIN(_00202_),
    .COUT(_00203_),
    .SUM(_00204_));
 sky130_fd_sc_hd__fa_1 _42289_ (.A(_00205_),
    .B(_00206_),
    .CIN(_00207_),
    .COUT(_00208_),
    .SUM(_00209_));
 sky130_fd_sc_hd__fa_1 _42290_ (.A(_00210_),
    .B(_00211_),
    .CIN(_00212_),
    .COUT(_00213_),
    .SUM(_00214_));
 sky130_fd_sc_hd__fa_1 _42291_ (.A(_00215_),
    .B(_00216_),
    .CIN(_00217_),
    .COUT(_00218_),
    .SUM(_00219_));
 sky130_fd_sc_hd__fa_1 _42292_ (.A(_00220_),
    .B(_20825_),
    .CIN(_00221_),
    .COUT(_20837_),
    .SUM(_20838_));
 sky130_fd_sc_hd__fa_1 _42293_ (.A(_00222_),
    .B(_20828_),
    .CIN(_20838_),
    .COUT(_00223_),
    .SUM(_00224_));
 sky130_fd_sc_hd__fa_1 _42294_ (.A(_00225_),
    .B(_00226_),
    .CIN(_00227_),
    .COUT(_20839_),
    .SUM(_20840_));
 sky130_fd_sc_hd__fa_1 _42295_ (.A(_00228_),
    .B(_00229_),
    .CIN(_00230_),
    .COUT(_00231_),
    .SUM(_00232_));
 sky130_fd_sc_hd__fa_1 _42296_ (.A(_00233_),
    .B(_00234_),
    .CIN(_00235_),
    .COUT(_00236_),
    .SUM(_00237_));
 sky130_fd_sc_hd__fa_1 _42297_ (.A(_00238_),
    .B(_00239_),
    .CIN(_00240_),
    .COUT(_20841_),
    .SUM(_20842_));
 sky130_fd_sc_hd__fa_1 _42298_ (.A(_00241_),
    .B(_20837_),
    .CIN(_20842_),
    .COUT(_00242_),
    .SUM(_00243_));
 sky130_fd_sc_hd__fa_1 _42299_ (.A(_00244_),
    .B(_00245_),
    .CIN(_00246_),
    .COUT(_20843_),
    .SUM(_20844_));
 sky130_fd_sc_hd__fa_1 _42300_ (.A(_00247_),
    .B(_00248_),
    .CIN(_00249_),
    .COUT(_00250_),
    .SUM(_00251_));
 sky130_fd_sc_hd__fa_1 _42301_ (.A(_00252_),
    .B(_00253_),
    .CIN(_00254_),
    .COUT(_00255_),
    .SUM(_00256_));
 sky130_fd_sc_hd__fa_1 _42302_ (.A(_00257_),
    .B(_00258_),
    .CIN(_00259_),
    .COUT(_20845_),
    .SUM(_20846_));
 sky130_fd_sc_hd__fa_1 _42303_ (.A(_00260_),
    .B(_20841_),
    .CIN(_20846_),
    .COUT(_00261_),
    .SUM(_00262_));
 sky130_fd_sc_hd__fa_1 _42304_ (.A(_00263_),
    .B(_00264_),
    .CIN(_00265_),
    .COUT(_00266_),
    .SUM(_00267_));
 sky130_fd_sc_hd__fa_1 _42305_ (.A(_00268_),
    .B(_00269_),
    .CIN(_00270_),
    .COUT(_20847_),
    .SUM(_20848_));
 sky130_fd_sc_hd__fa_1 _42306_ (.A(_00271_),
    .B(_00272_),
    .CIN(_00273_),
    .COUT(_00274_),
    .SUM(_00275_));
 sky130_fd_sc_hd__fa_1 _42307_ (.A(_00276_),
    .B(_00277_),
    .CIN(_00278_),
    .COUT(_00279_),
    .SUM(_00280_));
 sky130_fd_sc_hd__fa_1 _42308_ (.A(_00281_),
    .B(_00282_),
    .CIN(_00283_),
    .COUT(_20849_),
    .SUM(_20850_));
 sky130_fd_sc_hd__fa_1 _42309_ (.A(_00284_),
    .B(_20845_),
    .CIN(_20850_),
    .COUT(_00285_),
    .SUM(_00286_));
 sky130_fd_sc_hd__fa_1 _42310_ (.A(_00287_),
    .B(_20851_),
    .CIN(_20852_),
    .COUT(_20853_),
    .SUM(_20854_));
 sky130_fd_sc_hd__fa_1 _42311_ (.A(_20855_),
    .B(_20856_),
    .CIN(_20857_),
    .COUT(_20858_),
    .SUM(_00288_));
 sky130_fd_sc_hd__fa_1 _42312_ (.A(_00289_),
    .B(_00290_),
    .CIN(_00291_),
    .COUT(_00292_),
    .SUM(_00293_));
 sky130_fd_sc_hd__fa_1 _42313_ (.A(_00294_),
    .B(_00295_),
    .CIN(_00296_),
    .COUT(_20859_),
    .SUM(_00297_));
 sky130_fd_sc_hd__fa_1 _42314_ (.A(_00298_),
    .B(_00299_),
    .CIN(_00300_),
    .COUT(_00301_),
    .SUM(_20860_));
 sky130_fd_sc_hd__fa_1 _42315_ (.A(_20847_),
    .B(_20860_),
    .CIN(_20861_),
    .COUT(_20862_),
    .SUM(_20863_));
 sky130_fd_sc_hd__fa_1 _42316_ (.A(_00302_),
    .B(_00303_),
    .CIN(_00304_),
    .COUT(_00305_),
    .SUM(_00306_));
 sky130_fd_sc_hd__fa_1 _42317_ (.A(_00307_),
    .B(_00308_),
    .CIN(_00309_),
    .COUT(_00310_),
    .SUM(_00311_));
 sky130_fd_sc_hd__fa_1 _42318_ (.A(_00312_),
    .B(_00313_),
    .CIN(_00314_),
    .COUT(_20864_),
    .SUM(_20865_));
 sky130_fd_sc_hd__fa_1 _42319_ (.A(_00315_),
    .B(_20849_),
    .CIN(_20865_),
    .COUT(_00316_),
    .SUM(_00317_));
 sky130_fd_sc_hd__fa_1 _42320_ (.A(_00318_),
    .B(_20866_),
    .CIN(_20867_),
    .COUT(_20868_),
    .SUM(_20869_));
 sky130_fd_sc_hd__fa_1 _42321_ (.A(_20870_),
    .B(_20871_),
    .CIN(_20872_),
    .COUT(_20873_),
    .SUM(_20874_));
 sky130_fd_sc_hd__fa_1 _42322_ (.A(_20875_),
    .B(_20858_),
    .CIN(_20874_),
    .COUT(_20876_),
    .SUM(_20877_));
 sky130_fd_sc_hd__fa_1 _42323_ (.A(_00319_),
    .B(_00320_),
    .CIN(_00321_),
    .COUT(_20878_),
    .SUM(_00322_));
 sky130_fd_sc_hd__fa_1 _42324_ (.A(_00323_),
    .B(_00324_),
    .CIN(_00325_),
    .COUT(_20879_),
    .SUM(_20880_));
 sky130_fd_sc_hd__fa_1 _42325_ (.A(_00326_),
    .B(_20880_),
    .CIN(_20859_),
    .COUT(_00327_),
    .SUM(_00328_));
 sky130_fd_sc_hd__fa_1 _42326_ (.A(_00329_),
    .B(_00330_),
    .CIN(_00331_),
    .COUT(_00332_),
    .SUM(_00333_));
 sky130_fd_sc_hd__fa_1 _42327_ (.A(_00334_),
    .B(_00335_),
    .CIN(_00336_),
    .COUT(_00337_),
    .SUM(_00338_));
 sky130_fd_sc_hd__fa_1 _42328_ (.A(_00339_),
    .B(_00340_),
    .CIN(_00341_),
    .COUT(_20881_),
    .SUM(_20882_));
 sky130_fd_sc_hd__fa_1 _42329_ (.A(_00342_),
    .B(_20864_),
    .CIN(_20882_),
    .COUT(_00343_),
    .SUM(_00344_));
 sky130_fd_sc_hd__fa_1 _42330_ (.A(_00345_),
    .B(_20883_),
    .CIN(_20884_),
    .COUT(_20885_),
    .SUM(_20886_));
 sky130_fd_sc_hd__fa_1 _42331_ (.A(_20887_),
    .B(_20888_),
    .CIN(_20889_),
    .COUT(_20890_),
    .SUM(_20891_));
 sky130_fd_sc_hd__fa_1 _42332_ (.A(_20892_),
    .B(_20873_),
    .CIN(_20891_),
    .COUT(_20893_),
    .SUM(_20894_));
 sky130_fd_sc_hd__fa_1 _42333_ (.A(_00346_),
    .B(_00347_),
    .CIN(_00348_),
    .COUT(_20895_),
    .SUM(_00349_));
 sky130_fd_sc_hd__fa_1 _42334_ (.A(_00350_),
    .B(_00351_),
    .CIN(_00352_),
    .COUT(_00353_),
    .SUM(_00354_));
 sky130_fd_sc_hd__fa_1 _42335_ (.A(_20879_),
    .B(_00355_),
    .CIN(_20878_),
    .COUT(_00356_),
    .SUM(_00357_));
 sky130_fd_sc_hd__fa_1 _42336_ (.A(_00358_),
    .B(_00359_),
    .CIN(_20896_),
    .COUT(_00360_),
    .SUM(_20897_));
 sky130_fd_sc_hd__fa_1 _42337_ (.A(_00361_),
    .B(_00362_),
    .CIN(_00363_),
    .COUT(_00364_),
    .SUM(_00365_));
 sky130_fd_sc_hd__fa_1 _42338_ (.A(_00366_),
    .B(_00367_),
    .CIN(_00368_),
    .COUT(_00369_),
    .SUM(_00370_));
 sky130_fd_sc_hd__fa_1 _42339_ (.A(_00371_),
    .B(_00372_),
    .CIN(_00373_),
    .COUT(_20898_),
    .SUM(_20899_));
 sky130_fd_sc_hd__fa_1 _42340_ (.A(_00374_),
    .B(_20881_),
    .CIN(_20899_),
    .COUT(_00375_),
    .SUM(_00376_));
 sky130_fd_sc_hd__fa_1 _42341_ (.A(_00377_),
    .B(_20900_),
    .CIN(_20897_),
    .COUT(_20901_),
    .SUM(_20902_));
 sky130_fd_sc_hd__fa_1 _42342_ (.A(_20903_),
    .B(_20904_),
    .CIN(_20905_),
    .COUT(_20906_),
    .SUM(_20907_));
 sky130_fd_sc_hd__fa_1 _42343_ (.A(_20908_),
    .B(_20890_),
    .CIN(_20907_),
    .COUT(_20909_),
    .SUM(_20910_));
 sky130_fd_sc_hd__fa_1 _42344_ (.A(_00378_),
    .B(_00379_),
    .CIN(_00380_),
    .COUT(_00381_),
    .SUM(_00382_));
 sky130_fd_sc_hd__fa_1 _42345_ (.A(_00383_),
    .B(_00384_),
    .CIN(_00385_),
    .COUT(_20911_),
    .SUM(_20912_));
 sky130_fd_sc_hd__fa_1 _42346_ (.A(_20912_),
    .B(_00386_),
    .CIN(_00387_),
    .COUT(_20913_),
    .SUM(_00388_));
 sky130_fd_sc_hd__fa_1 _42347_ (.A(_00389_),
    .B(_00390_),
    .CIN(_00391_),
    .COUT(_00392_),
    .SUM(_00393_));
 sky130_fd_sc_hd__fa_1 _42348_ (.A(_00394_),
    .B(_00395_),
    .CIN(_20895_),
    .COUT(_20914_),
    .SUM(_00396_));
 sky130_fd_sc_hd__fa_1 _42349_ (.A(_00397_),
    .B(_00398_),
    .CIN(_20915_),
    .COUT(_00399_),
    .SUM(_00400_));
 sky130_fd_sc_hd__fa_1 _42350_ (.A(_00401_),
    .B(_00402_),
    .CIN(_00403_),
    .COUT(_00404_),
    .SUM(_00405_));
 sky130_fd_sc_hd__fa_1 _42351_ (.A(_00406_),
    .B(_00407_),
    .CIN(_00408_),
    .COUT(_00409_),
    .SUM(_00410_));
 sky130_fd_sc_hd__fa_1 _42352_ (.A(_00411_),
    .B(_00412_),
    .CIN(_00413_),
    .COUT(_20916_),
    .SUM(_20917_));
 sky130_fd_sc_hd__fa_1 _42353_ (.A(_00414_),
    .B(_20898_),
    .CIN(_20917_),
    .COUT(_00415_),
    .SUM(_20918_));
 sky130_fd_sc_hd__fa_1 _42354_ (.A(_20918_),
    .B(_00416_),
    .CIN(_00417_),
    .COUT(_00418_),
    .SUM(_00419_));
 sky130_fd_sc_hd__fa_1 _42355_ (.A(_20919_),
    .B(_20920_),
    .CIN(_20921_),
    .COUT(_20922_),
    .SUM(_20923_));
 sky130_fd_sc_hd__fa_1 _42356_ (.A(_20924_),
    .B(_20906_),
    .CIN(_20923_),
    .COUT(_20925_),
    .SUM(_20926_));
 sky130_fd_sc_hd__fa_1 _42357_ (.A(_00420_),
    .B(_00421_),
    .CIN(_00422_),
    .COUT(_20927_),
    .SUM(_20928_));
 sky130_fd_sc_hd__fa_1 _42358_ (.A(_00423_),
    .B(_00424_),
    .CIN(_00425_),
    .COUT(_20929_),
    .SUM(_20930_));
 sky130_fd_sc_hd__fa_1 _42359_ (.A(_20930_),
    .B(_00426_),
    .CIN(_20928_),
    .COUT(_20931_),
    .SUM(_00427_));
 sky130_fd_sc_hd__fa_1 _42360_ (.A(_00428_),
    .B(_00429_),
    .CIN(_00430_),
    .COUT(_20932_),
    .SUM(_20933_));
 sky130_fd_sc_hd__fa_1 _42361_ (.A(_00431_),
    .B(_20933_),
    .CIN(_20911_),
    .COUT(_20934_),
    .SUM(_20935_));
 sky130_fd_sc_hd__fa_1 _42362_ (.A(_20914_),
    .B(_20935_),
    .CIN(_20913_),
    .COUT(_20936_),
    .SUM(_20937_));
 sky130_fd_sc_hd__fa_1 _42363_ (.A(_00432_),
    .B(_00433_),
    .CIN(_00434_),
    .COUT(_00435_),
    .SUM(_00436_));
 sky130_fd_sc_hd__fa_1 _42364_ (.A(_00437_),
    .B(_00438_),
    .CIN(_00439_),
    .COUT(_00440_),
    .SUM(_00441_));
 sky130_fd_sc_hd__fa_1 _42365_ (.A(_00442_),
    .B(_00443_),
    .CIN(_00444_),
    .COUT(_20938_),
    .SUM(_20939_));
 sky130_fd_sc_hd__fa_1 _42366_ (.A(_00445_),
    .B(_20916_),
    .CIN(_20939_),
    .COUT(_00446_),
    .SUM(_20940_));
 sky130_fd_sc_hd__fa_1 _42367_ (.A(_20940_),
    .B(_00447_),
    .CIN(_20937_),
    .COUT(_00448_),
    .SUM(_00449_));
 sky130_fd_sc_hd__fa_1 _42368_ (.A(_00450_),
    .B(_00451_),
    .CIN(_00452_),
    .COUT(_20941_),
    .SUM(_00453_));
 sky130_fd_sc_hd__fa_1 _42369_ (.A(_20942_),
    .B(_20922_),
    .CIN(_00454_),
    .COUT(_20943_),
    .SUM(_20944_));
 sky130_fd_sc_hd__fa_1 _42370_ (.A(_00455_),
    .B(_00456_),
    .CIN(_00457_),
    .COUT(_20945_),
    .SUM(_20946_));
 sky130_fd_sc_hd__fa_1 _42371_ (.A(_00458_),
    .B(_00459_),
    .CIN(_00460_),
    .COUT(_20947_),
    .SUM(_20948_));
 sky130_fd_sc_hd__fa_1 _42372_ (.A(_20948_),
    .B(_20927_),
    .CIN(_20946_),
    .COUT(_20949_),
    .SUM(_00461_));
 sky130_fd_sc_hd__fa_1 _42373_ (.A(_00462_),
    .B(_00463_),
    .CIN(_00464_),
    .COUT(_20950_),
    .SUM(_20951_));
 sky130_fd_sc_hd__fa_1 _42374_ (.A(_20932_),
    .B(_20951_),
    .CIN(_20929_),
    .COUT(_20952_),
    .SUM(_20953_));
 sky130_fd_sc_hd__fa_1 _42375_ (.A(_20934_),
    .B(_20953_),
    .CIN(_20931_),
    .COUT(_20954_),
    .SUM(_20955_));
 sky130_fd_sc_hd__fa_1 _42376_ (.A(_00466_),
    .B(_00467_),
    .CIN(_00468_),
    .COUT(_20956_),
    .SUM(_20957_));
 sky130_fd_sc_hd__fa_1 _42377_ (.A(_00469_),
    .B(_00470_),
    .CIN(_00471_),
    .COUT(_00472_),
    .SUM(_00473_));
 sky130_fd_sc_hd__fa_1 _42378_ (.A(_00474_),
    .B(_00475_),
    .CIN(_20957_),
    .COUT(_20958_),
    .SUM(_20959_));
 sky130_fd_sc_hd__fa_1 _42379_ (.A(_00476_),
    .B(_20938_),
    .CIN(_20959_),
    .COUT(_00477_),
    .SUM(_20960_));
 sky130_fd_sc_hd__fa_1 _42380_ (.A(_20960_),
    .B(_20936_),
    .CIN(_20955_),
    .COUT(_20961_),
    .SUM(_00478_));
 sky130_fd_sc_hd__fa_1 _42381_ (.A(_00479_),
    .B(_00480_),
    .CIN(_00481_),
    .COUT(_20962_),
    .SUM(_20963_));
 sky130_fd_sc_hd__fa_1 _42382_ (.A(_00482_),
    .B(_20941_),
    .CIN(_20963_),
    .COUT(_00483_),
    .SUM(_00484_));
 sky130_fd_sc_hd__fa_1 _42383_ (.A(_00486_),
    .B(_00487_),
    .CIN(_00488_),
    .COUT(_20964_),
    .SUM(_20965_));
 sky130_fd_sc_hd__fa_1 _42384_ (.A(_00489_),
    .B(_00490_),
    .CIN(_00491_),
    .COUT(_20966_),
    .SUM(_20967_));
 sky130_fd_sc_hd__fa_1 _42385_ (.A(_00492_),
    .B(_00493_),
    .CIN(_00494_),
    .COUT(_20968_),
    .SUM(_20969_));
 sky130_fd_sc_hd__fa_1 _42386_ (.A(_20969_),
    .B(_20945_),
    .CIN(_20967_),
    .COUT(_20970_),
    .SUM(_00495_));
 sky130_fd_sc_hd__fa_1 _42387_ (.A(_00496_),
    .B(_00497_),
    .CIN(_00498_),
    .COUT(_00499_),
    .SUM(_00500_));
 sky130_fd_sc_hd__fa_1 _42388_ (.A(_20950_),
    .B(_00501_),
    .CIN(_20947_),
    .COUT(_20971_),
    .SUM(_20972_));
 sky130_fd_sc_hd__fa_1 _42389_ (.A(_20952_),
    .B(_20972_),
    .CIN(_20949_),
    .COUT(_20973_),
    .SUM(_20974_));
 sky130_fd_sc_hd__fa_1 _42390_ (.A(_00502_),
    .B(_00503_),
    .CIN(_00504_),
    .COUT(_20975_),
    .SUM(_20976_));
 sky130_fd_sc_hd__fa_1 _42391_ (.A(_00505_),
    .B(_00506_),
    .CIN(_00507_),
    .COUT(_00508_),
    .SUM(_00509_));
 sky130_fd_sc_hd__fa_1 _42392_ (.A(_00510_),
    .B(_20956_),
    .CIN(_20976_),
    .COUT(_20977_),
    .SUM(_20978_));
 sky130_fd_sc_hd__fa_1 _42393_ (.A(_00511_),
    .B(_20958_),
    .CIN(_20978_),
    .COUT(_00512_),
    .SUM(_20979_));
 sky130_fd_sc_hd__fa_1 _42394_ (.A(_20979_),
    .B(_20954_),
    .CIN(_20974_),
    .COUT(_20980_),
    .SUM(_20981_));
 sky130_fd_sc_hd__fa_1 _42395_ (.A(_20961_),
    .B(_20981_),
    .CIN(_00513_),
    .COUT(_00514_),
    .SUM(_00515_));
 sky130_fd_sc_hd__fa_1 _42396_ (.A(_20982_),
    .B(_20983_),
    .CIN(_20984_),
    .COUT(_00516_),
    .SUM(_00517_));
 sky130_fd_sc_hd__fa_1 _42397_ (.A(_00518_),
    .B(_20962_),
    .CIN(_00519_),
    .COUT(_00520_),
    .SUM(_00521_));
 sky130_fd_sc_hd__fa_1 _42398_ (.A(_00523_),
    .B(_00524_),
    .CIN(_00525_),
    .COUT(_20985_),
    .SUM(_20986_));
 sky130_fd_sc_hd__fa_1 _42399_ (.A(_00526_),
    .B(_00527_),
    .CIN(_00528_),
    .COUT(_20987_),
    .SUM(_20988_));
 sky130_fd_sc_hd__fa_1 _42400_ (.A(_00529_),
    .B(_00530_),
    .CIN(_00531_),
    .COUT(_00532_),
    .SUM(_00533_));
 sky130_fd_sc_hd__fa_1 _42401_ (.A(_00534_),
    .B(_20966_),
    .CIN(_20988_),
    .COUT(_20989_),
    .SUM(_00535_));
 sky130_fd_sc_hd__fa_1 _42402_ (.A(_00536_),
    .B(_20990_),
    .CIN(_20991_),
    .COUT(_20992_),
    .SUM(_20993_));
 sky130_fd_sc_hd__fa_1 _42403_ (.A(_00537_),
    .B(_00538_),
    .CIN(_00539_),
    .COUT(_00540_),
    .SUM(_00541_));
 sky130_fd_sc_hd__fa_1 _42404_ (.A(_00542_),
    .B(_00543_),
    .CIN(_20968_),
    .COUT(_20994_),
    .SUM(_20995_));
 sky130_fd_sc_hd__fa_1 _42405_ (.A(_20971_),
    .B(_20995_),
    .CIN(_20970_),
    .COUT(_20996_),
    .SUM(_20997_));
 sky130_fd_sc_hd__fa_1 _42406_ (.A(_00544_),
    .B(_00545_),
    .CIN(_00546_),
    .COUT(_20998_),
    .SUM(_20999_));
 sky130_fd_sc_hd__fa_1 _42407_ (.A(_00547_),
    .B(_00548_),
    .CIN(_00549_),
    .COUT(_00550_),
    .SUM(_00551_));
 sky130_fd_sc_hd__fa_1 _42408_ (.A(_00552_),
    .B(_20975_),
    .CIN(_20999_),
    .COUT(_21000_),
    .SUM(_21001_));
 sky130_fd_sc_hd__fa_1 _42409_ (.A(_00553_),
    .B(_20977_),
    .CIN(_21001_),
    .COUT(_00554_),
    .SUM(_21002_));
 sky130_fd_sc_hd__fa_1 _42410_ (.A(_21002_),
    .B(_20973_),
    .CIN(_20997_),
    .COUT(_21003_),
    .SUM(_21004_));
 sky130_fd_sc_hd__fa_1 _42411_ (.A(_20980_),
    .B(_21004_),
    .CIN(_00555_),
    .COUT(_00556_),
    .SUM(_00557_));
 sky130_fd_sc_hd__fa_1 _42412_ (.A(_00558_),
    .B(_00559_),
    .CIN(_00560_),
    .COUT(_21005_),
    .SUM(_21006_));
 sky130_fd_sc_hd__fa_1 _42413_ (.A(_00561_),
    .B(_00562_),
    .CIN(_21006_),
    .COUT(_00563_),
    .SUM(_00564_));
 sky130_fd_sc_hd__fa_1 _42414_ (.A(_00566_),
    .B(_00567_),
    .CIN(_00568_),
    .COUT(_00569_),
    .SUM(_00570_));
 sky130_fd_sc_hd__fa_1 _42415_ (.A(_00571_),
    .B(_00572_),
    .CIN(_00573_),
    .COUT(_21007_),
    .SUM(_21008_));
 sky130_fd_sc_hd__fa_1 _42416_ (.A(_00574_),
    .B(_00575_),
    .CIN(_00576_),
    .COUT(_21009_),
    .SUM(_21010_));
 sky130_fd_sc_hd__fa_1 _42417_ (.A(_21010_),
    .B(_20987_),
    .CIN(_21008_),
    .COUT(_21011_),
    .SUM(_00577_));
 sky130_fd_sc_hd__fa_1 _42418_ (.A(_00578_),
    .B(_21012_),
    .CIN(_21013_),
    .COUT(_21014_),
    .SUM(_21015_));
 sky130_fd_sc_hd__fa_1 _42419_ (.A(_00579_),
    .B(_00580_),
    .CIN(_00581_),
    .COUT(_00582_),
    .SUM(_00583_));
 sky130_fd_sc_hd__fa_1 _42420_ (.A(_00584_),
    .B(_00585_),
    .CIN(_00586_),
    .COUT(_21016_),
    .SUM(_21017_));
 sky130_fd_sc_hd__fa_1 _42421_ (.A(_20994_),
    .B(_21017_),
    .CIN(_20989_),
    .COUT(_21018_),
    .SUM(_21019_));
 sky130_fd_sc_hd__fa_1 _42422_ (.A(_00587_),
    .B(_00588_),
    .CIN(_00589_),
    .COUT(_21020_),
    .SUM(_21021_));
 sky130_fd_sc_hd__fa_1 _42423_ (.A(_00590_),
    .B(_00591_),
    .CIN(_00592_),
    .COUT(_00593_),
    .SUM(_00594_));
 sky130_fd_sc_hd__fa_1 _42424_ (.A(_00595_),
    .B(_20998_),
    .CIN(_21021_),
    .COUT(_21022_),
    .SUM(_21023_));
 sky130_fd_sc_hd__fa_1 _42425_ (.A(_00596_),
    .B(_21000_),
    .CIN(_21023_),
    .COUT(_00597_),
    .SUM(_21024_));
 sky130_fd_sc_hd__fa_1 _42426_ (.A(_21024_),
    .B(_20996_),
    .CIN(_21019_),
    .COUT(_21025_),
    .SUM(_21026_));
 sky130_fd_sc_hd__fa_1 _42427_ (.A(_21003_),
    .B(_21026_),
    .CIN(_00598_),
    .COUT(_00599_),
    .SUM(_00600_));
 sky130_fd_sc_hd__fa_1 _42428_ (.A(_00601_),
    .B(_21027_),
    .CIN(_21028_),
    .COUT(_00602_),
    .SUM(_00603_));
 sky130_fd_sc_hd__fa_1 _42429_ (.A(_00604_),
    .B(_00605_),
    .CIN(_00606_),
    .COUT(_21029_),
    .SUM(_21030_));
 sky130_fd_sc_hd__fa_1 _42430_ (.A(_00607_),
    .B(_21005_),
    .CIN(_21030_),
    .COUT(_00608_),
    .SUM(_00609_));
 sky130_fd_sc_hd__fa_1 _42431_ (.A(_00611_),
    .B(_00612_),
    .CIN(_00613_),
    .COUT(_21031_),
    .SUM(_00614_));
 sky130_fd_sc_hd__fa_1 _42432_ (.A(_00615_),
    .B(_00616_),
    .CIN(_00617_),
    .COUT(_21032_),
    .SUM(_00618_));
 sky130_fd_sc_hd__fa_1 _42433_ (.A(_00619_),
    .B(_00620_),
    .CIN(_21033_),
    .COUT(_00621_),
    .SUM(_21034_));
 sky130_fd_sc_hd__fa_1 _42434_ (.A(_00622_),
    .B(_00623_),
    .CIN(_00624_),
    .COUT(_21035_),
    .SUM(_21036_));
 sky130_fd_sc_hd__fa_1 _42435_ (.A(_00625_),
    .B(_00626_),
    .CIN(_00627_),
    .COUT(_21037_),
    .SUM(_21038_));
 sky130_fd_sc_hd__fa_1 _42436_ (.A(_21038_),
    .B(_21007_),
    .CIN(_21036_),
    .COUT(_21039_),
    .SUM(_00628_));
 sky130_fd_sc_hd__fa_1 _42437_ (.A(_00629_),
    .B(_21040_),
    .CIN(_21034_),
    .COUT(_21041_),
    .SUM(_21042_));
 sky130_fd_sc_hd__fa_1 _42438_ (.A(_00630_),
    .B(_00631_),
    .CIN(_00632_),
    .COUT(_00633_),
    .SUM(_00634_));
 sky130_fd_sc_hd__fa_1 _42439_ (.A(_00635_),
    .B(_00636_),
    .CIN(_21009_),
    .COUT(_21043_),
    .SUM(_21044_));
 sky130_fd_sc_hd__fa_1 _42440_ (.A(_21016_),
    .B(_21044_),
    .CIN(_21011_),
    .COUT(_21045_),
    .SUM(_21046_));
 sky130_fd_sc_hd__fa_1 _42441_ (.A(_00637_),
    .B(_00638_),
    .CIN(_00639_),
    .COUT(_21047_),
    .SUM(_21048_));
 sky130_fd_sc_hd__fa_1 _42442_ (.A(_00640_),
    .B(_00641_),
    .CIN(_00642_),
    .COUT(_00643_),
    .SUM(_00644_));
 sky130_fd_sc_hd__fa_1 _42443_ (.A(_00645_),
    .B(_21020_),
    .CIN(_21048_),
    .COUT(_21049_),
    .SUM(_21050_));
 sky130_fd_sc_hd__fa_1 _42444_ (.A(_00646_),
    .B(_21022_),
    .CIN(_21050_),
    .COUT(_00647_),
    .SUM(_21051_));
 sky130_fd_sc_hd__fa_1 _42445_ (.A(_21051_),
    .B(_21018_),
    .CIN(_21046_),
    .COUT(_21052_),
    .SUM(_21053_));
 sky130_fd_sc_hd__fa_1 _42446_ (.A(_21025_),
    .B(_21053_),
    .CIN(_00648_),
    .COUT(_00649_),
    .SUM(_00650_));
 sky130_fd_sc_hd__fa_1 _42447_ (.A(_00651_),
    .B(_21054_),
    .CIN(_21055_),
    .COUT(_00652_),
    .SUM(_00653_));
 sky130_fd_sc_hd__fa_1 _42448_ (.A(_00654_),
    .B(_00655_),
    .CIN(_00656_),
    .COUT(_21056_),
    .SUM(_21057_));
 sky130_fd_sc_hd__fa_1 _42449_ (.A(_00657_),
    .B(_21029_),
    .CIN(_21057_),
    .COUT(_00658_),
    .SUM(_00659_));
 sky130_fd_sc_hd__fa_1 _42450_ (.A(_00661_),
    .B(_00662_),
    .CIN(_00663_),
    .COUT(_21058_),
    .SUM(_00664_));
 sky130_fd_sc_hd__fa_1 _42451_ (.A(_00665_),
    .B(_00666_),
    .CIN(_00667_),
    .COUT(_21059_),
    .SUM(_21060_));
 sky130_fd_sc_hd__fa_1 _42452_ (.A(_21032_),
    .B(_21060_),
    .CIN(_21031_),
    .COUT(_00668_),
    .SUM(_21061_));
 sky130_fd_sc_hd__fa_1 _42453_ (.A(_00669_),
    .B(_00670_),
    .CIN(_00671_),
    .COUT(_21062_),
    .SUM(_21063_));
 sky130_fd_sc_hd__fa_1 _42454_ (.A(_00672_),
    .B(_00673_),
    .CIN(_00674_),
    .COUT(_21064_),
    .SUM(_21065_));
 sky130_fd_sc_hd__fa_1 _42455_ (.A(_21065_),
    .B(_21035_),
    .CIN(_21063_),
    .COUT(_21066_),
    .SUM(_21067_));
 sky130_fd_sc_hd__fa_1 _42456_ (.A(_21067_),
    .B(_00675_),
    .CIN(_21061_),
    .COUT(_00676_),
    .SUM(_00677_));
 sky130_fd_sc_hd__fa_1 _42457_ (.A(_00678_),
    .B(_00679_),
    .CIN(_00680_),
    .COUT(_00681_),
    .SUM(_00682_));
 sky130_fd_sc_hd__fa_1 _42458_ (.A(_00683_),
    .B(_00684_),
    .CIN(_21037_),
    .COUT(_21068_),
    .SUM(_21069_));
 sky130_fd_sc_hd__fa_1 _42459_ (.A(_21043_),
    .B(_21069_),
    .CIN(_21039_),
    .COUT(_21070_),
    .SUM(_21071_));
 sky130_fd_sc_hd__fa_1 _42460_ (.A(_00685_),
    .B(_00686_),
    .CIN(_00687_),
    .COUT(_21072_),
    .SUM(_21073_));
 sky130_fd_sc_hd__fa_1 _42461_ (.A(_00688_),
    .B(_00689_),
    .CIN(_00690_),
    .COUT(_00691_),
    .SUM(_00692_));
 sky130_fd_sc_hd__fa_1 _42462_ (.A(_00693_),
    .B(_21047_),
    .CIN(_21073_),
    .COUT(_21074_),
    .SUM(_21075_));
 sky130_fd_sc_hd__fa_1 _42463_ (.A(_00694_),
    .B(_21049_),
    .CIN(_21075_),
    .COUT(_00695_),
    .SUM(_21076_));
 sky130_fd_sc_hd__fa_1 _42464_ (.A(_21076_),
    .B(_21045_),
    .CIN(_21071_),
    .COUT(_21077_),
    .SUM(_21078_));
 sky130_fd_sc_hd__fa_1 _42465_ (.A(_21052_),
    .B(_21078_),
    .CIN(_00696_),
    .COUT(_00697_),
    .SUM(_00698_));
 sky130_fd_sc_hd__fa_1 _42466_ (.A(_00699_),
    .B(_21079_),
    .CIN(_21080_),
    .COUT(_00700_),
    .SUM(_00701_));
 sky130_fd_sc_hd__fa_1 _42467_ (.A(_00702_),
    .B(_00703_),
    .CIN(_00704_),
    .COUT(_21081_),
    .SUM(_21082_));
 sky130_fd_sc_hd__fa_1 _42468_ (.A(_00705_),
    .B(_21056_),
    .CIN(_21082_),
    .COUT(_00706_),
    .SUM(_00707_));
 sky130_fd_sc_hd__fa_1 _42469_ (.A(_00709_),
    .B(_00710_),
    .CIN(_00711_),
    .COUT(_21083_),
    .SUM(_00712_));
 sky130_fd_sc_hd__fa_1 _42470_ (.A(_00713_),
    .B(_00714_),
    .CIN(_00715_),
    .COUT(_21084_),
    .SUM(_21085_));
 sky130_fd_sc_hd__fa_1 _42471_ (.A(_21059_),
    .B(_21085_),
    .CIN(_21058_),
    .COUT(_21086_),
    .SUM(_00716_));
 sky130_fd_sc_hd__fa_1 _42472_ (.A(_00717_),
    .B(_00718_),
    .CIN(_00719_),
    .COUT(_21087_),
    .SUM(_21088_));
 sky130_fd_sc_hd__fa_1 _42473_ (.A(_00720_),
    .B(_00721_),
    .CIN(_00722_),
    .COUT(_21089_),
    .SUM(_21090_));
 sky130_fd_sc_hd__fa_1 _42474_ (.A(_21090_),
    .B(_21062_),
    .CIN(_21088_),
    .COUT(_21091_),
    .SUM(_00723_));
 sky130_fd_sc_hd__fa_1 _42475_ (.A(_00724_),
    .B(_00725_),
    .CIN(_00726_),
    .COUT(_00727_),
    .SUM(_21092_));
 sky130_fd_sc_hd__fa_1 _42476_ (.A(_00728_),
    .B(_00729_),
    .CIN(_00730_),
    .COUT(_00731_),
    .SUM(_00732_));
 sky130_fd_sc_hd__fa_1 _42477_ (.A(_00733_),
    .B(_00734_),
    .CIN(_21064_),
    .COUT(_21093_),
    .SUM(_21094_));
 sky130_fd_sc_hd__fa_1 _42478_ (.A(_21068_),
    .B(_21094_),
    .CIN(_21066_),
    .COUT(_21095_),
    .SUM(_21096_));
 sky130_fd_sc_hd__fa_1 _42479_ (.A(_00735_),
    .B(_00736_),
    .CIN(_00737_),
    .COUT(_21097_),
    .SUM(_21098_));
 sky130_fd_sc_hd__fa_1 _42480_ (.A(_00738_),
    .B(_00739_),
    .CIN(_00740_),
    .COUT(_00741_),
    .SUM(_00742_));
 sky130_fd_sc_hd__fa_1 _42481_ (.A(_00743_),
    .B(_21072_),
    .CIN(_21098_),
    .COUT(_21099_),
    .SUM(_21100_));
 sky130_fd_sc_hd__fa_1 _42482_ (.A(_00744_),
    .B(_21074_),
    .CIN(_21100_),
    .COUT(_00745_),
    .SUM(_21101_));
 sky130_fd_sc_hd__fa_1 _42483_ (.A(_21101_),
    .B(_21070_),
    .CIN(_21096_),
    .COUT(_00746_),
    .SUM(_21102_));
 sky130_fd_sc_hd__fa_1 _42484_ (.A(_21077_),
    .B(_21102_),
    .CIN(_00747_),
    .COUT(_00748_),
    .SUM(_21103_));
 sky130_fd_sc_hd__fa_1 _42485_ (.A(_21103_),
    .B(_00749_),
    .CIN(_00750_),
    .COUT(_21104_),
    .SUM(_21105_));
 sky130_fd_sc_hd__fa_1 _42486_ (.A(_00751_),
    .B(_00752_),
    .CIN(_21105_),
    .COUT(_21106_),
    .SUM(_21107_));
 sky130_fd_sc_hd__fa_1 _42487_ (.A(_00753_),
    .B(_21081_),
    .CIN(_21107_),
    .COUT(_00754_),
    .SUM(_00755_));
 sky130_fd_sc_hd__fa_1 _42488_ (.A(_00757_),
    .B(_00758_),
    .CIN(_00759_),
    .COUT(_00760_),
    .SUM(_00761_));
 sky130_fd_sc_hd__fa_1 _42489_ (.A(_00762_),
    .B(_00763_),
    .CIN(_00764_),
    .COUT(_21108_),
    .SUM(_21109_));
 sky130_fd_sc_hd__fa_1 _42490_ (.A(_21109_),
    .B(_00765_),
    .CIN(_00766_),
    .COUT(_00767_),
    .SUM(_00768_));
 sky130_fd_sc_hd__fa_1 _42491_ (.A(_00769_),
    .B(_00770_),
    .CIN(_00771_),
    .COUT(_21110_),
    .SUM(_21111_));
 sky130_fd_sc_hd__fa_1 _42492_ (.A(_21084_),
    .B(_21111_),
    .CIN(_21083_),
    .COUT(_21112_),
    .SUM(_21113_));
 sky130_fd_sc_hd__fa_1 _42493_ (.A(_00772_),
    .B(_00773_),
    .CIN(_00774_),
    .COUT(_21114_),
    .SUM(_21115_));
 sky130_fd_sc_hd__fa_1 _42494_ (.A(_00775_),
    .B(_00776_),
    .CIN(_00777_),
    .COUT(_21116_),
    .SUM(_21117_));
 sky130_fd_sc_hd__fa_1 _42495_ (.A(_21117_),
    .B(_21087_),
    .CIN(_21115_),
    .COUT(_21118_),
    .SUM(_21119_));
 sky130_fd_sc_hd__fa_1 _42496_ (.A(_21119_),
    .B(_21086_),
    .CIN(_21113_),
    .COUT(_21120_),
    .SUM(_21121_));
 sky130_fd_sc_hd__fa_1 _42497_ (.A(_00778_),
    .B(_21121_),
    .CIN(_00779_),
    .COUT(_00780_),
    .SUM(_00781_));
 sky130_fd_sc_hd__fa_1 _42498_ (.A(_00782_),
    .B(_00783_),
    .CIN(_00784_),
    .COUT(_00785_),
    .SUM(_00786_));
 sky130_fd_sc_hd__fa_1 _42499_ (.A(_00787_),
    .B(_00788_),
    .CIN(_21089_),
    .COUT(_21122_),
    .SUM(_21123_));
 sky130_fd_sc_hd__fa_1 _42500_ (.A(_21093_),
    .B(_21123_),
    .CIN(_21091_),
    .COUT(_21124_),
    .SUM(_21125_));
 sky130_fd_sc_hd__fa_1 _42501_ (.A(_00789_),
    .B(_00790_),
    .CIN(_00791_),
    .COUT(_21126_),
    .SUM(_21127_));
 sky130_fd_sc_hd__fa_1 _42502_ (.A(_00792_),
    .B(_00793_),
    .CIN(_00794_),
    .COUT(_00795_),
    .SUM(_00796_));
 sky130_fd_sc_hd__fa_1 _42503_ (.A(_00797_),
    .B(_21097_),
    .CIN(_21127_),
    .COUT(_21128_),
    .SUM(_21129_));
 sky130_fd_sc_hd__fa_1 _42504_ (.A(_00798_),
    .B(_21099_),
    .CIN(_21129_),
    .COUT(_00799_),
    .SUM(_21130_));
 sky130_fd_sc_hd__fa_1 _42505_ (.A(_21130_),
    .B(_21095_),
    .CIN(_21125_),
    .COUT(_00800_),
    .SUM(_00801_));
 sky130_fd_sc_hd__fa_1 _42506_ (.A(_00802_),
    .B(_00803_),
    .CIN(_21131_),
    .COUT(_21132_),
    .SUM(_21133_));
 sky130_fd_sc_hd__fa_1 _42507_ (.A(_21133_),
    .B(_21134_),
    .CIN(_21135_),
    .COUT(_00804_),
    .SUM(_00805_));
 sky130_fd_sc_hd__fa_1 _42508_ (.A(_00806_),
    .B(_21104_),
    .CIN(_00807_),
    .COUT(_21136_),
    .SUM(_21137_));
 sky130_fd_sc_hd__fa_1 _42509_ (.A(_00808_),
    .B(_21106_),
    .CIN(_21137_),
    .COUT(_00809_),
    .SUM(_00810_));
 sky130_fd_sc_hd__fa_1 _42510_ (.A(_00812_),
    .B(_00813_),
    .CIN(_00814_),
    .COUT(_21138_),
    .SUM(_21139_));
 sky130_fd_sc_hd__fa_1 _42511_ (.A(_00815_),
    .B(_00816_),
    .CIN(_00817_),
    .COUT(_21140_),
    .SUM(_21141_));
 sky130_fd_sc_hd__fa_1 _42512_ (.A(_21141_),
    .B(_00818_),
    .CIN(_21139_),
    .COUT(_00819_),
    .SUM(_00820_));
 sky130_fd_sc_hd__fa_1 _42513_ (.A(_00821_),
    .B(_00822_),
    .CIN(_00823_),
    .COUT(_21142_),
    .SUM(_21143_));
 sky130_fd_sc_hd__fa_1 _42514_ (.A(_21110_),
    .B(_21143_),
    .CIN(_21108_),
    .COUT(_21144_),
    .SUM(_21145_));
 sky130_fd_sc_hd__fa_1 _42515_ (.A(_00824_),
    .B(_00825_),
    .CIN(_00826_),
    .COUT(_00827_),
    .SUM(_00828_));
 sky130_fd_sc_hd__fa_1 _42516_ (.A(_00829_),
    .B(_00830_),
    .CIN(_00831_),
    .COUT(_21146_),
    .SUM(_21147_));
 sky130_fd_sc_hd__fa_1 _42517_ (.A(_21147_),
    .B(_21114_),
    .CIN(_00832_),
    .COUT(_21148_),
    .SUM(_21149_));
 sky130_fd_sc_hd__fa_1 _42518_ (.A(_21149_),
    .B(_21112_),
    .CIN(_21145_),
    .COUT(_21150_),
    .SUM(_21151_));
 sky130_fd_sc_hd__fa_1 _42519_ (.A(_21120_),
    .B(_21151_),
    .CIN(_00833_),
    .COUT(_00834_),
    .SUM(_00835_));
 sky130_fd_sc_hd__fa_1 _42520_ (.A(_00836_),
    .B(_00837_),
    .CIN(_00838_),
    .COUT(_00839_),
    .SUM(_00840_));
 sky130_fd_sc_hd__fa_1 _42521_ (.A(_00841_),
    .B(_00842_),
    .CIN(_21116_),
    .COUT(_21152_),
    .SUM(_21153_));
 sky130_fd_sc_hd__fa_1 _42522_ (.A(_21122_),
    .B(_21153_),
    .CIN(_21118_),
    .COUT(_21154_),
    .SUM(_21155_));
 sky130_fd_sc_hd__fa_1 _42523_ (.A(_00843_),
    .B(_00844_),
    .CIN(_00845_),
    .COUT(_21156_),
    .SUM(_21157_));
 sky130_fd_sc_hd__fa_1 _42524_ (.A(_00846_),
    .B(_00847_),
    .CIN(_00848_),
    .COUT(_00849_),
    .SUM(_00850_));
 sky130_fd_sc_hd__fa_1 _42525_ (.A(_00851_),
    .B(_21126_),
    .CIN(_21157_),
    .COUT(_21158_),
    .SUM(_21159_));
 sky130_fd_sc_hd__fa_1 _42526_ (.A(_00852_),
    .B(_21128_),
    .CIN(_21159_),
    .COUT(_00853_),
    .SUM(_21160_));
 sky130_fd_sc_hd__fa_1 _42527_ (.A(_21160_),
    .B(_21124_),
    .CIN(_21155_),
    .COUT(_00854_),
    .SUM(_00855_));
 sky130_fd_sc_hd__fa_1 _42528_ (.A(_00856_),
    .B(_00857_),
    .CIN(_00858_),
    .COUT(_21161_),
    .SUM(_00859_));
 sky130_fd_sc_hd__fa_1 _42529_ (.A(_00860_),
    .B(_00861_),
    .CIN(_00862_),
    .COUT(_21162_),
    .SUM(_21163_));
 sky130_fd_sc_hd__fa_1 _42530_ (.A(_00863_),
    .B(_00864_),
    .CIN(_21163_),
    .COUT(_21164_),
    .SUM(_21165_));
 sky130_fd_sc_hd__fa_1 _42531_ (.A(_00865_),
    .B(_21136_),
    .CIN(_21165_),
    .COUT(_00866_),
    .SUM(_00867_));
 sky130_fd_sc_hd__fa_1 _42532_ (.A(_00869_),
    .B(_00870_),
    .CIN(_00871_),
    .COUT(_21166_),
    .SUM(_21167_));
 sky130_fd_sc_hd__fa_1 _42533_ (.A(_00872_),
    .B(_00873_),
    .CIN(_00874_),
    .COUT(_21168_),
    .SUM(_21169_));
 sky130_fd_sc_hd__fa_1 _42534_ (.A(_21169_),
    .B(_21138_),
    .CIN(_21167_),
    .COUT(_00875_),
    .SUM(_00876_));
 sky130_fd_sc_hd__fa_1 _42535_ (.A(_00877_),
    .B(_00878_),
    .CIN(_00879_),
    .COUT(_21170_),
    .SUM(_21171_));
 sky130_fd_sc_hd__fa_1 _42536_ (.A(_21142_),
    .B(_21171_),
    .CIN(_21140_),
    .COUT(_21172_),
    .SUM(_21173_));
 sky130_fd_sc_hd__fa_1 _42537_ (.A(_00880_),
    .B(_00881_),
    .CIN(_00882_),
    .COUT(_21174_),
    .SUM(_21175_));
 sky130_fd_sc_hd__fa_1 _42538_ (.A(_00883_),
    .B(_00884_),
    .CIN(_00885_),
    .COUT(_21176_),
    .SUM(_21177_));
 sky130_fd_sc_hd__fa_1 _42539_ (.A(_21177_),
    .B(_00886_),
    .CIN(_21175_),
    .COUT(_21178_),
    .SUM(_21179_));
 sky130_fd_sc_hd__fa_1 _42540_ (.A(_21179_),
    .B(_21144_),
    .CIN(_21173_),
    .COUT(_21180_),
    .SUM(_21181_));
 sky130_fd_sc_hd__fa_1 _42541_ (.A(_21150_),
    .B(_21181_),
    .CIN(_00887_),
    .COUT(_00888_),
    .SUM(_00889_));
 sky130_fd_sc_hd__fa_1 _42542_ (.A(_00890_),
    .B(_21182_),
    .CIN(_21183_),
    .COUT(_00891_),
    .SUM(_00892_));
 sky130_fd_sc_hd__fa_1 _42543_ (.A(_00893_),
    .B(_00894_),
    .CIN(_00895_),
    .COUT(_00896_),
    .SUM(_00897_));
 sky130_fd_sc_hd__fa_1 _42544_ (.A(_00898_),
    .B(_00899_),
    .CIN(_21146_),
    .COUT(_21184_),
    .SUM(_21185_));
 sky130_fd_sc_hd__fa_1 _42545_ (.A(_21152_),
    .B(_21185_),
    .CIN(_21148_),
    .COUT(_21186_),
    .SUM(_21187_));
 sky130_fd_sc_hd__fa_1 _42546_ (.A(_00900_),
    .B(_00901_),
    .CIN(_00902_),
    .COUT(_21188_),
    .SUM(_21189_));
 sky130_fd_sc_hd__fa_1 _42547_ (.A(_00903_),
    .B(_00904_),
    .CIN(_00905_),
    .COUT(_00906_),
    .SUM(_00907_));
 sky130_fd_sc_hd__fa_1 _42548_ (.A(_00908_),
    .B(_21156_),
    .CIN(_21189_),
    .COUT(_21190_),
    .SUM(_21191_));
 sky130_fd_sc_hd__fa_1 _42549_ (.A(_00909_),
    .B(_21158_),
    .CIN(_21191_),
    .COUT(_00910_),
    .SUM(_21192_));
 sky130_fd_sc_hd__fa_1 _42550_ (.A(_21192_),
    .B(_21154_),
    .CIN(_21187_),
    .COUT(_00911_),
    .SUM(_00912_));
 sky130_fd_sc_hd__fa_1 _42551_ (.A(_00913_),
    .B(_00914_),
    .CIN(_00915_),
    .COUT(_21193_),
    .SUM(_00916_));
 sky130_fd_sc_hd__fa_1 _42552_ (.A(_00917_),
    .B(_00918_),
    .CIN(_00919_),
    .COUT(_21194_),
    .SUM(_21195_));
 sky130_fd_sc_hd__fa_1 _42553_ (.A(_00920_),
    .B(_21162_),
    .CIN(_21195_),
    .COUT(_21196_),
    .SUM(_21197_));
 sky130_fd_sc_hd__fa_1 _42554_ (.A(_00921_),
    .B(_21164_),
    .CIN(_21197_),
    .COUT(_00922_),
    .SUM(_00923_));
 sky130_fd_sc_hd__fa_1 _42555_ (.A(_00925_),
    .B(_00926_),
    .CIN(_00927_),
    .COUT(_21198_),
    .SUM(_21199_));
 sky130_fd_sc_hd__fa_1 _42556_ (.A(_00928_),
    .B(_00929_),
    .CIN(_00930_),
    .COUT(_21200_),
    .SUM(_21201_));
 sky130_fd_sc_hd__fa_1 _42557_ (.A(_00931_),
    .B(_00932_),
    .CIN(_00933_),
    .COUT(_21202_),
    .SUM(_21203_));
 sky130_fd_sc_hd__fa_1 _42558_ (.A(_21203_),
    .B(_21166_),
    .CIN(_21201_),
    .COUT(_21204_),
    .SUM(_00934_));
 sky130_fd_sc_hd__fa_1 _42559_ (.A(_00935_),
    .B(_00936_),
    .CIN(_00937_),
    .COUT(_21205_),
    .SUM(_21206_));
 sky130_fd_sc_hd__fa_1 _42560_ (.A(_21170_),
    .B(_21206_),
    .CIN(_21168_),
    .COUT(_21207_),
    .SUM(_21208_));
 sky130_fd_sc_hd__fa_1 _42561_ (.A(_00938_),
    .B(_00939_),
    .CIN(_00940_),
    .COUT(_21209_),
    .SUM(_21210_));
 sky130_fd_sc_hd__fa_1 _42562_ (.A(_00941_),
    .B(_00942_),
    .CIN(_00943_),
    .COUT(_21211_),
    .SUM(_21212_));
 sky130_fd_sc_hd__fa_1 _42563_ (.A(_21212_),
    .B(_21174_),
    .CIN(_21210_),
    .COUT(_21213_),
    .SUM(_21214_));
 sky130_fd_sc_hd__fa_1 _42564_ (.A(_21214_),
    .B(_21172_),
    .CIN(_21208_),
    .COUT(_21215_),
    .SUM(_21216_));
 sky130_fd_sc_hd__fa_1 _42565_ (.A(_21180_),
    .B(_21216_),
    .CIN(_00944_),
    .COUT(_00945_),
    .SUM(_21217_));
 sky130_fd_sc_hd__fa_1 _42566_ (.A(_21217_),
    .B(_00946_),
    .CIN(_00947_),
    .COUT(_21218_),
    .SUM(_21219_));
 sky130_fd_sc_hd__fa_1 _42567_ (.A(_00948_),
    .B(_00949_),
    .CIN(_00950_),
    .COUT(_00951_),
    .SUM(_00952_));
 sky130_fd_sc_hd__fa_1 _42568_ (.A(_00953_),
    .B(_00954_),
    .CIN(_21176_),
    .COUT(_21220_),
    .SUM(_21221_));
 sky130_fd_sc_hd__fa_1 _42569_ (.A(_21184_),
    .B(_21221_),
    .CIN(_21178_),
    .COUT(_21222_),
    .SUM(_21223_));
 sky130_fd_sc_hd__fa_1 _42570_ (.A(_00955_),
    .B(_00956_),
    .CIN(_00957_),
    .COUT(_21224_),
    .SUM(_21225_));
 sky130_fd_sc_hd__fa_1 _42571_ (.A(_00958_),
    .B(_00959_),
    .CIN(_00960_),
    .COUT(_00961_),
    .SUM(_00962_));
 sky130_fd_sc_hd__fa_1 _42572_ (.A(_00963_),
    .B(_21188_),
    .CIN(_21225_),
    .COUT(_21226_),
    .SUM(_21227_));
 sky130_fd_sc_hd__fa_1 _42573_ (.A(_00964_),
    .B(_21190_),
    .CIN(_21227_),
    .COUT(_00965_),
    .SUM(_21228_));
 sky130_fd_sc_hd__fa_1 _42574_ (.A(_21228_),
    .B(_21186_),
    .CIN(_21223_),
    .COUT(_00966_),
    .SUM(_00967_));
 sky130_fd_sc_hd__fa_1 _42575_ (.A(_00968_),
    .B(_00969_),
    .CIN(_00970_),
    .COUT(_21229_),
    .SUM(_00971_));
 sky130_fd_sc_hd__fa_1 _42576_ (.A(_00972_),
    .B(_00973_),
    .CIN(_21219_),
    .COUT(_21230_),
    .SUM(_21231_));
 sky130_fd_sc_hd__fa_1 _42577_ (.A(_00974_),
    .B(_21194_),
    .CIN(_21231_),
    .COUT(_21232_),
    .SUM(_21233_));
 sky130_fd_sc_hd__fa_1 _42578_ (.A(_00975_),
    .B(_21196_),
    .CIN(_21233_),
    .COUT(_00976_),
    .SUM(_00977_));
 sky130_fd_sc_hd__fa_1 _42579_ (.A(_00979_),
    .B(_00980_),
    .CIN(_00981_),
    .COUT(_00982_),
    .SUM(_00983_));
 sky130_fd_sc_hd__fa_1 _42580_ (.A(_00984_),
    .B(_00985_),
    .CIN(_00986_),
    .COUT(_21234_),
    .SUM(_21235_));
 sky130_fd_sc_hd__fa_1 _42581_ (.A(_00987_),
    .B(_00988_),
    .CIN(_00989_),
    .COUT(_21236_),
    .SUM(_21237_));
 sky130_fd_sc_hd__fa_1 _42582_ (.A(_21237_),
    .B(_21200_),
    .CIN(_21235_),
    .COUT(_21238_),
    .SUM(_21239_));
 sky130_fd_sc_hd__fa_1 _42583_ (.A(_21204_),
    .B(_21239_),
    .CIN(_00990_),
    .COUT(_21240_),
    .SUM(_00991_));
 sky130_fd_sc_hd__fa_1 _42584_ (.A(_00992_),
    .B(_00993_),
    .CIN(_00994_),
    .COUT(_00995_),
    .SUM(_00996_));
 sky130_fd_sc_hd__fa_1 _42585_ (.A(_21205_),
    .B(_00997_),
    .CIN(_21202_),
    .COUT(_21241_),
    .SUM(_21242_));
 sky130_fd_sc_hd__fa_1 _42586_ (.A(_00998_),
    .B(_00999_),
    .CIN(_01000_),
    .COUT(_21243_),
    .SUM(_21244_));
 sky130_fd_sc_hd__fa_1 _42587_ (.A(_01001_),
    .B(_01002_),
    .CIN(_01003_),
    .COUT(_21245_),
    .SUM(_21246_));
 sky130_fd_sc_hd__fa_1 _42588_ (.A(_21246_),
    .B(_21209_),
    .CIN(_21244_),
    .COUT(_21247_),
    .SUM(_21248_));
 sky130_fd_sc_hd__fa_1 _42589_ (.A(_21248_),
    .B(_21207_),
    .CIN(_21242_),
    .COUT(_21249_),
    .SUM(_21250_));
 sky130_fd_sc_hd__fa_1 _42590_ (.A(_21215_),
    .B(_21250_),
    .CIN(_01004_),
    .COUT(_01005_),
    .SUM(_21251_));
 sky130_fd_sc_hd__fa_1 _42591_ (.A(_21251_),
    .B(_01006_),
    .CIN(_01007_),
    .COUT(_21252_),
    .SUM(_21253_));
 sky130_fd_sc_hd__fa_1 _42592_ (.A(_01008_),
    .B(_01009_),
    .CIN(_01010_),
    .COUT(_01011_),
    .SUM(_01012_));
 sky130_fd_sc_hd__fa_1 _42593_ (.A(_01013_),
    .B(_01014_),
    .CIN(_21211_),
    .COUT(_21254_),
    .SUM(_21255_));
 sky130_fd_sc_hd__fa_1 _42594_ (.A(_21220_),
    .B(_21255_),
    .CIN(_21213_),
    .COUT(_21256_),
    .SUM(_21257_));
 sky130_fd_sc_hd__fa_1 _42595_ (.A(_01015_),
    .B(_01016_),
    .CIN(_01017_),
    .COUT(_21258_),
    .SUM(_21259_));
 sky130_fd_sc_hd__fa_1 _42596_ (.A(_01018_),
    .B(_01019_),
    .CIN(_01020_),
    .COUT(_01021_),
    .SUM(_01022_));
 sky130_fd_sc_hd__fa_1 _42597_ (.A(_01023_),
    .B(_21224_),
    .CIN(_21259_),
    .COUT(_21260_),
    .SUM(_21261_));
 sky130_fd_sc_hd__fa_1 _42598_ (.A(_01024_),
    .B(_21226_),
    .CIN(_21261_),
    .COUT(_01025_),
    .SUM(_21262_));
 sky130_fd_sc_hd__fa_1 _42599_ (.A(_21262_),
    .B(_21222_),
    .CIN(_21257_),
    .COUT(_01026_),
    .SUM(_01027_));
 sky130_fd_sc_hd__fa_1 _42600_ (.A(_01028_),
    .B(_01029_),
    .CIN(_01030_),
    .COUT(_21263_),
    .SUM(_01031_));
 sky130_fd_sc_hd__fa_1 _42601_ (.A(_01032_),
    .B(_21218_),
    .CIN(_21253_),
    .COUT(_21264_),
    .SUM(_21265_));
 sky130_fd_sc_hd__fa_1 _42602_ (.A(_01033_),
    .B(_21230_),
    .CIN(_21265_),
    .COUT(_21266_),
    .SUM(_21267_));
 sky130_fd_sc_hd__fa_1 _42603_ (.A(_01034_),
    .B(_21232_),
    .CIN(_21267_),
    .COUT(_01035_),
    .SUM(_01036_));
 sky130_fd_sc_hd__fa_1 _42604_ (.A(_01038_),
    .B(_01039_),
    .CIN(_01040_),
    .COUT(_21268_),
    .SUM(_01041_));
 sky130_fd_sc_hd__fa_1 _42605_ (.A(_01042_),
    .B(_01043_),
    .CIN(_01044_),
    .COUT(_21269_),
    .SUM(_21270_));
 sky130_fd_sc_hd__fa_1 _42606_ (.A(_01045_),
    .B(_01046_),
    .CIN(_01047_),
    .COUT(_21271_),
    .SUM(_21272_));
 sky130_fd_sc_hd__fa_1 _42607_ (.A(_21272_),
    .B(_21234_),
    .CIN(_21270_),
    .COUT(_21273_),
    .SUM(_21274_));
 sky130_fd_sc_hd__fa_1 _42608_ (.A(_21238_),
    .B(_21274_),
    .CIN(_01048_),
    .COUT(_21275_),
    .SUM(_01049_));
 sky130_fd_sc_hd__fa_1 _42609_ (.A(_01050_),
    .B(_21276_),
    .CIN(_21277_),
    .COUT(_01051_),
    .SUM(_01052_));
 sky130_fd_sc_hd__fa_1 _42610_ (.A(_01053_),
    .B(_01054_),
    .CIN(_01055_),
    .COUT(_01056_),
    .SUM(_01057_));
 sky130_fd_sc_hd__fa_1 _42611_ (.A(_01058_),
    .B(_01059_),
    .CIN(_21236_),
    .COUT(_21278_),
    .SUM(_21279_));
 sky130_fd_sc_hd__fa_1 _42612_ (.A(_01060_),
    .B(_01061_),
    .CIN(_01062_),
    .COUT(_21280_),
    .SUM(_21281_));
 sky130_fd_sc_hd__fa_1 _42613_ (.A(_01063_),
    .B(_01064_),
    .CIN(_01065_),
    .COUT(_21282_),
    .SUM(_21283_));
 sky130_fd_sc_hd__fa_1 _42614_ (.A(_21283_),
    .B(_21243_),
    .CIN(_21281_),
    .COUT(_21284_),
    .SUM(_21285_));
 sky130_fd_sc_hd__fa_1 _42615_ (.A(_21285_),
    .B(_21241_),
    .CIN(_21279_),
    .COUT(_21286_),
    .SUM(_21287_));
 sky130_fd_sc_hd__fa_1 _42616_ (.A(_21249_),
    .B(_21287_),
    .CIN(_21240_),
    .COUT(_01066_),
    .SUM(_21288_));
 sky130_fd_sc_hd__fa_1 _42617_ (.A(_21288_),
    .B(_01067_),
    .CIN(_01068_),
    .COUT(_21289_),
    .SUM(_21290_));
 sky130_fd_sc_hd__fa_1 _42618_ (.A(_01069_),
    .B(_01070_),
    .CIN(_01071_),
    .COUT(_21291_),
    .SUM(_21292_));
 sky130_fd_sc_hd__fa_1 _42619_ (.A(_01072_),
    .B(_21292_),
    .CIN(_21245_),
    .COUT(_21293_),
    .SUM(_21294_));
 sky130_fd_sc_hd__fa_1 _42620_ (.A(_21254_),
    .B(_21294_),
    .CIN(_21247_),
    .COUT(_21295_),
    .SUM(_21296_));
 sky130_fd_sc_hd__fa_1 _42621_ (.A(_01073_),
    .B(_01074_),
    .CIN(_01075_),
    .COUT(_01076_),
    .SUM(_01077_));
 sky130_fd_sc_hd__fa_1 _42622_ (.A(_01078_),
    .B(_01079_),
    .CIN(_01080_),
    .COUT(_01081_),
    .SUM(_01082_));
 sky130_fd_sc_hd__fa_1 _42623_ (.A(_01083_),
    .B(_21258_),
    .CIN(_01084_),
    .COUT(_21297_),
    .SUM(_21298_));
 sky130_fd_sc_hd__fa_1 _42624_ (.A(_01085_),
    .B(_21260_),
    .CIN(_21298_),
    .COUT(_01086_),
    .SUM(_21299_));
 sky130_fd_sc_hd__fa_1 _42625_ (.A(_21299_),
    .B(_21256_),
    .CIN(_21296_),
    .COUT(_01087_),
    .SUM(_01088_));
 sky130_fd_sc_hd__fa_1 _42626_ (.A(_01089_),
    .B(_01090_),
    .CIN(_01091_),
    .COUT(_21300_),
    .SUM(_01092_));
 sky130_fd_sc_hd__fa_1 _42627_ (.A(_01093_),
    .B(_21252_),
    .CIN(_21290_),
    .COUT(_21301_),
    .SUM(_21302_));
 sky130_fd_sc_hd__fa_1 _42628_ (.A(_01094_),
    .B(_21264_),
    .CIN(_21302_),
    .COUT(_21303_),
    .SUM(_21304_));
 sky130_fd_sc_hd__fa_1 _42629_ (.A(_01095_),
    .B(_21266_),
    .CIN(_21304_),
    .COUT(_01096_),
    .SUM(_01097_));
 sky130_fd_sc_hd__fa_1 _42630_ (.A(_01099_),
    .B(_01100_),
    .CIN(_01101_),
    .COUT(_21305_),
    .SUM(_01102_));
 sky130_fd_sc_hd__fa_1 _42631_ (.A(_01103_),
    .B(_01104_),
    .CIN(_01105_),
    .COUT(_21306_),
    .SUM(_21307_));
 sky130_fd_sc_hd__fa_1 _42632_ (.A(_21268_),
    .B(_21307_),
    .CIN(_01106_),
    .COUT(_21308_),
    .SUM(_01107_));
 sky130_fd_sc_hd__fa_1 _42633_ (.A(_01108_),
    .B(_01109_),
    .CIN(_01110_),
    .COUT(_21309_),
    .SUM(_21310_));
 sky130_fd_sc_hd__fa_1 _42634_ (.A(_01111_),
    .B(_01112_),
    .CIN(_01113_),
    .COUT(_21311_),
    .SUM(_21312_));
 sky130_fd_sc_hd__fa_1 _42635_ (.A(_21312_),
    .B(_21269_),
    .CIN(_21310_),
    .COUT(_21313_),
    .SUM(_21314_));
 sky130_fd_sc_hd__fa_1 _42636_ (.A(_21273_),
    .B(_21314_),
    .CIN(_01114_),
    .COUT(_21315_),
    .SUM(_21316_));
 sky130_fd_sc_hd__fa_1 _42637_ (.A(_21316_),
    .B(_01115_),
    .CIN(_01116_),
    .COUT(_21317_),
    .SUM(_21318_));
 sky130_fd_sc_hd__fa_1 _42638_ (.A(_01117_),
    .B(_01118_),
    .CIN(_01119_),
    .COUT(_01120_),
    .SUM(_01121_));
 sky130_fd_sc_hd__fa_1 _42639_ (.A(_01122_),
    .B(_01123_),
    .CIN(_21271_),
    .COUT(_21319_),
    .SUM(_21320_));
 sky130_fd_sc_hd__fa_1 _42640_ (.A(_01124_),
    .B(_01125_),
    .CIN(_01126_),
    .COUT(_21321_),
    .SUM(_21322_));
 sky130_fd_sc_hd__fa_1 _42641_ (.A(_01127_),
    .B(_01128_),
    .CIN(_01129_),
    .COUT(_21323_),
    .SUM(_21324_));
 sky130_fd_sc_hd__fa_1 _42642_ (.A(_21324_),
    .B(_21280_),
    .CIN(_21322_),
    .COUT(_21325_),
    .SUM(_21326_));
 sky130_fd_sc_hd__fa_1 _42643_ (.A(_21326_),
    .B(_21278_),
    .CIN(_21320_),
    .COUT(_21327_),
    .SUM(_21328_));
 sky130_fd_sc_hd__fa_1 _42644_ (.A(_21286_),
    .B(_21328_),
    .CIN(_21275_),
    .COUT(_01130_),
    .SUM(_21329_));
 sky130_fd_sc_hd__fa_1 _42645_ (.A(_21329_),
    .B(_01131_),
    .CIN(_21318_),
    .COUT(_21330_),
    .SUM(_21331_));
 sky130_fd_sc_hd__fa_1 _42646_ (.A(_01132_),
    .B(_01133_),
    .CIN(_01134_),
    .COUT(_01135_),
    .SUM(_01136_));
 sky130_fd_sc_hd__fa_1 _42647_ (.A(_21291_),
    .B(_01137_),
    .CIN(_21282_),
    .COUT(_21332_),
    .SUM(_21333_));
 sky130_fd_sc_hd__fa_1 _42648_ (.A(_21293_),
    .B(_21333_),
    .CIN(_21284_),
    .COUT(_21334_),
    .SUM(_21335_));
 sky130_fd_sc_hd__fa_1 _42649_ (.A(_01138_),
    .B(_01139_),
    .CIN(_01140_),
    .COUT(_01141_),
    .SUM(_01142_));
 sky130_fd_sc_hd__fa_1 _42650_ (.A(_01143_),
    .B(_01144_),
    .CIN(_01145_),
    .COUT(_01146_),
    .SUM(_01147_));
 sky130_fd_sc_hd__fa_1 _42651_ (.A(_01148_),
    .B(_01149_),
    .CIN(_01150_),
    .COUT(_21336_),
    .SUM(_21337_));
 sky130_fd_sc_hd__fa_1 _42652_ (.A(_01151_),
    .B(_21297_),
    .CIN(_21337_),
    .COUT(_01152_),
    .SUM(_21338_));
 sky130_fd_sc_hd__fa_1 _42653_ (.A(_21338_),
    .B(_21295_),
    .CIN(_21335_),
    .COUT(_01153_),
    .SUM(_01154_));
 sky130_fd_sc_hd__fa_1 _42654_ (.A(_01155_),
    .B(_01156_),
    .CIN(_01157_),
    .COUT(_21339_),
    .SUM(_01158_));
 sky130_fd_sc_hd__fa_1 _42655_ (.A(_01159_),
    .B(_21289_),
    .CIN(_21331_),
    .COUT(_21340_),
    .SUM(_21341_));
 sky130_fd_sc_hd__fa_1 _42656_ (.A(_01160_),
    .B(_21301_),
    .CIN(_21341_),
    .COUT(_21342_),
    .SUM(_21343_));
 sky130_fd_sc_hd__fa_1 _42657_ (.A(_01161_),
    .B(_21303_),
    .CIN(_21343_),
    .COUT(_01162_),
    .SUM(_01163_));
 sky130_fd_sc_hd__fa_1 _42658_ (.A(_01165_),
    .B(_01166_),
    .CIN(_01167_),
    .COUT(_21344_),
    .SUM(_01168_));
 sky130_fd_sc_hd__fa_1 _42659_ (.A(_01169_),
    .B(_01170_),
    .CIN(_01171_),
    .COUT(_21345_),
    .SUM(_21346_));
 sky130_fd_sc_hd__fa_1 _42660_ (.A(_21306_),
    .B(_21346_),
    .CIN(_21305_),
    .COUT(_21347_),
    .SUM(_01172_));
 sky130_fd_sc_hd__fa_1 _42661_ (.A(_01173_),
    .B(_01174_),
    .CIN(_01175_),
    .COUT(_21348_),
    .SUM(_21349_));
 sky130_fd_sc_hd__fa_1 _42662_ (.A(_01176_),
    .B(_01177_),
    .CIN(_01178_),
    .COUT(_21350_),
    .SUM(_21351_));
 sky130_fd_sc_hd__fa_1 _42663_ (.A(_21351_),
    .B(_21309_),
    .CIN(_21349_),
    .COUT(_21352_),
    .SUM(_21353_));
 sky130_fd_sc_hd__fa_1 _42664_ (.A(_21313_),
    .B(_21353_),
    .CIN(_21308_),
    .COUT(_21354_),
    .SUM(_01179_));
 sky130_fd_sc_hd__fa_1 _42665_ (.A(_01180_),
    .B(_21355_),
    .CIN(_21356_),
    .COUT(_01181_),
    .SUM(_01182_));
 sky130_fd_sc_hd__fa_1 _42666_ (.A(_01183_),
    .B(_01184_),
    .CIN(_01185_),
    .COUT(_21357_),
    .SUM(_21358_));
 sky130_fd_sc_hd__fa_1 _42667_ (.A(_01186_),
    .B(_21358_),
    .CIN(_21311_),
    .COUT(_21359_),
    .SUM(_21360_));
 sky130_fd_sc_hd__fa_1 _42668_ (.A(_01187_),
    .B(_01188_),
    .CIN(_01189_),
    .COUT(_21361_),
    .SUM(_21362_));
 sky130_fd_sc_hd__fa_1 _42669_ (.A(_01190_),
    .B(_01191_),
    .CIN(_01192_),
    .COUT(_21363_),
    .SUM(_21364_));
 sky130_fd_sc_hd__fa_1 _42670_ (.A(_21364_),
    .B(_21321_),
    .CIN(_21362_),
    .COUT(_21365_),
    .SUM(_21366_));
 sky130_fd_sc_hd__fa_1 _42671_ (.A(_21366_),
    .B(_21319_),
    .CIN(_21360_),
    .COUT(_21367_),
    .SUM(_21368_));
 sky130_fd_sc_hd__fa_1 _42672_ (.A(_21327_),
    .B(_21368_),
    .CIN(_21315_),
    .COUT(_21369_),
    .SUM(_21370_));
 sky130_fd_sc_hd__fa_1 _42673_ (.A(_21370_),
    .B(_21317_),
    .CIN(_01193_),
    .COUT(_21371_),
    .SUM(_21372_));
 sky130_fd_sc_hd__fa_1 _42674_ (.A(_01194_),
    .B(_01195_),
    .CIN(_01196_),
    .COUT(_01197_),
    .SUM(_01198_));
 sky130_fd_sc_hd__fa_1 _42675_ (.A(_01199_),
    .B(_01200_),
    .CIN(_21323_),
    .COUT(_21373_),
    .SUM(_21374_));
 sky130_fd_sc_hd__fa_1 _42676_ (.A(_21332_),
    .B(_21374_),
    .CIN(_21325_),
    .COUT(_21375_),
    .SUM(_21376_));
 sky130_fd_sc_hd__fa_1 _42677_ (.A(_01201_),
    .B(_01202_),
    .CIN(_01203_),
    .COUT(_01204_),
    .SUM(_01205_));
 sky130_fd_sc_hd__fa_1 _42678_ (.A(_01206_),
    .B(_01207_),
    .CIN(_01208_),
    .COUT(_01209_),
    .SUM(_01210_));
 sky130_fd_sc_hd__fa_1 _42679_ (.A(_01211_),
    .B(_01212_),
    .CIN(_01213_),
    .COUT(_21377_),
    .SUM(_21378_));
 sky130_fd_sc_hd__fa_1 _42680_ (.A(_01214_),
    .B(_21336_),
    .CIN(_21378_),
    .COUT(_01215_),
    .SUM(_21379_));
 sky130_fd_sc_hd__fa_1 _42681_ (.A(_21379_),
    .B(_21334_),
    .CIN(_21376_),
    .COUT(_21380_),
    .SUM(_01216_));
 sky130_fd_sc_hd__fa_1 _42682_ (.A(_01217_),
    .B(_01218_),
    .CIN(_01219_),
    .COUT(_21381_),
    .SUM(_01220_));
 sky130_fd_sc_hd__fa_1 _42683_ (.A(_01221_),
    .B(_21330_),
    .CIN(_21372_),
    .COUT(_21382_),
    .SUM(_21383_));
 sky130_fd_sc_hd__fa_1 _42684_ (.A(_01222_),
    .B(_21340_),
    .CIN(_21383_),
    .COUT(_21384_),
    .SUM(_21385_));
 sky130_fd_sc_hd__fa_1 _42685_ (.A(_01223_),
    .B(_21342_),
    .CIN(_21385_),
    .COUT(_01224_),
    .SUM(_01225_));
 sky130_fd_sc_hd__fa_1 _42686_ (.A(_01227_),
    .B(_01228_),
    .CIN(_01229_),
    .COUT(_21386_),
    .SUM(_01230_));
 sky130_fd_sc_hd__fa_1 _42687_ (.A(_01231_),
    .B(_01232_),
    .CIN(_01233_),
    .COUT(_21387_),
    .SUM(_21388_));
 sky130_fd_sc_hd__fa_1 _42688_ (.A(_21345_),
    .B(_21388_),
    .CIN(_21344_),
    .COUT(_21389_),
    .SUM(_21390_));
 sky130_fd_sc_hd__fa_1 _42689_ (.A(_21390_),
    .B(_01234_),
    .CIN(_01235_),
    .COUT(_21391_),
    .SUM(_21392_));
 sky130_fd_sc_hd__fa_1 _42690_ (.A(_01236_),
    .B(_01237_),
    .CIN(_01238_),
    .COUT(_21393_),
    .SUM(_21394_));
 sky130_fd_sc_hd__fa_1 _42691_ (.A(_01239_),
    .B(_01240_),
    .CIN(_01241_),
    .COUT(_21395_),
    .SUM(_21396_));
 sky130_fd_sc_hd__fa_1 _42692_ (.A(_21396_),
    .B(_21348_),
    .CIN(_21394_),
    .COUT(_21397_),
    .SUM(_21398_));
 sky130_fd_sc_hd__fa_1 _42693_ (.A(_21352_),
    .B(_21398_),
    .CIN(_21347_),
    .COUT(_21399_),
    .SUM(_21400_));
 sky130_fd_sc_hd__fa_1 _42694_ (.A(_21400_),
    .B(_01242_),
    .CIN(_21392_),
    .COUT(_21401_),
    .SUM(_21402_));
 sky130_fd_sc_hd__fa_1 _42695_ (.A(_01243_),
    .B(_01244_),
    .CIN(_01245_),
    .COUT(_01246_),
    .SUM(_01247_));
 sky130_fd_sc_hd__fa_1 _42696_ (.A(_21357_),
    .B(_01248_),
    .CIN(_21350_),
    .COUT(_21403_),
    .SUM(_21404_));
 sky130_fd_sc_hd__fa_1 _42697_ (.A(_01249_),
    .B(_01250_),
    .CIN(_01251_),
    .COUT(_21405_),
    .SUM(_21406_));
 sky130_fd_sc_hd__fa_1 _42698_ (.A(_01252_),
    .B(_01253_),
    .CIN(_01254_),
    .COUT(_21407_),
    .SUM(_21408_));
 sky130_fd_sc_hd__fa_1 _42699_ (.A(_21408_),
    .B(_21361_),
    .CIN(_21406_),
    .COUT(_21409_),
    .SUM(_21410_));
 sky130_fd_sc_hd__fa_1 _42700_ (.A(_21410_),
    .B(_21359_),
    .CIN(_21404_),
    .COUT(_21411_),
    .SUM(_21412_));
 sky130_fd_sc_hd__fa_1 _42701_ (.A(_21367_),
    .B(_21412_),
    .CIN(_21354_),
    .COUT(_01255_),
    .SUM(_21413_));
 sky130_fd_sc_hd__fa_1 _42702_ (.A(_21413_),
    .B(_01256_),
    .CIN(_21402_),
    .COUT(_21414_),
    .SUM(_21415_));
 sky130_fd_sc_hd__fa_1 _42703_ (.A(_01257_),
    .B(_01258_),
    .CIN(_01259_),
    .COUT(_01260_),
    .SUM(_01261_));
 sky130_fd_sc_hd__fa_1 _42704_ (.A(_01262_),
    .B(_01263_),
    .CIN(_21363_),
    .COUT(_21416_),
    .SUM(_21417_));
 sky130_fd_sc_hd__fa_1 _42705_ (.A(_21373_),
    .B(_21417_),
    .CIN(_21365_),
    .COUT(_21418_),
    .SUM(_21419_));
 sky130_fd_sc_hd__fa_1 _42706_ (.A(_01264_),
    .B(_01265_),
    .CIN(_01266_),
    .COUT(_01267_),
    .SUM(_01268_));
 sky130_fd_sc_hd__fa_1 _42707_ (.A(_01269_),
    .B(_01270_),
    .CIN(_01271_),
    .COUT(_01272_),
    .SUM(_01273_));
 sky130_fd_sc_hd__fa_1 _42708_ (.A(_01274_),
    .B(_01275_),
    .CIN(_01276_),
    .COUT(_21420_),
    .SUM(_21421_));
 sky130_fd_sc_hd__fa_1 _42709_ (.A(_01277_),
    .B(_21377_),
    .CIN(_21421_),
    .COUT(_01278_),
    .SUM(_21422_));
 sky130_fd_sc_hd__fa_1 _42710_ (.A(_21422_),
    .B(_21375_),
    .CIN(_21419_),
    .COUT(_01279_),
    .SUM(_21423_));
 sky130_fd_sc_hd__fa_1 _42711_ (.A(_21380_),
    .B(_21423_),
    .CIN(_21369_),
    .COUT(_01280_),
    .SUM(_21424_));
 sky130_fd_sc_hd__fa_1 _42712_ (.A(_21424_),
    .B(_21371_),
    .CIN(_21415_),
    .COUT(_21425_),
    .SUM(_21426_));
 sky130_fd_sc_hd__fa_1 _42713_ (.A(_01281_),
    .B(_21382_),
    .CIN(_21426_),
    .COUT(_21427_),
    .SUM(_21428_));
 sky130_fd_sc_hd__fa_1 _42714_ (.A(_01282_),
    .B(_21384_),
    .CIN(_21428_),
    .COUT(_01283_),
    .SUM(_01284_));
 sky130_fd_sc_hd__fa_1 _42715_ (.A(_01286_),
    .B(_01287_),
    .CIN(_01288_),
    .COUT(_21429_),
    .SUM(_21430_));
 sky130_fd_sc_hd__fa_1 _42716_ (.A(_21430_),
    .B(_01289_),
    .CIN(_01290_),
    .COUT(_21431_),
    .SUM(_21432_));
 sky130_fd_sc_hd__fa_1 _42717_ (.A(_01291_),
    .B(_01292_),
    .CIN(_01293_),
    .COUT(_21433_),
    .SUM(_21434_));
 sky130_fd_sc_hd__fa_1 _42718_ (.A(_21387_),
    .B(_21434_),
    .CIN(_21386_),
    .COUT(_21435_),
    .SUM(_21436_));
 sky130_fd_sc_hd__fa_1 _42719_ (.A(_21436_),
    .B(_01294_),
    .CIN(_21432_),
    .COUT(_21437_),
    .SUM(_21438_));
 sky130_fd_sc_hd__fa_1 _42720_ (.A(_01295_),
    .B(_01296_),
    .CIN(_01297_),
    .COUT(_21439_),
    .SUM(_21440_));
 sky130_fd_sc_hd__fa_1 _42721_ (.A(_01298_),
    .B(_01299_),
    .CIN(_01300_),
    .COUT(_21441_),
    .SUM(_21442_));
 sky130_fd_sc_hd__fa_1 _42722_ (.A(_21442_),
    .B(_21393_),
    .CIN(_21440_),
    .COUT(_21443_),
    .SUM(_21444_));
 sky130_fd_sc_hd__fa_1 _42723_ (.A(_21397_),
    .B(_21444_),
    .CIN(_21389_),
    .COUT(_21445_),
    .SUM(_21446_));
 sky130_fd_sc_hd__fa_1 _42724_ (.A(_21446_),
    .B(_21391_),
    .CIN(_21438_),
    .COUT(_21447_),
    .SUM(_21448_));
 sky130_fd_sc_hd__fa_1 _42725_ (.A(_01301_),
    .B(_01302_),
    .CIN(_01303_),
    .COUT(_21449_),
    .SUM(_21450_));
 sky130_fd_sc_hd__fa_1 _42726_ (.A(_01304_),
    .B(_21450_),
    .CIN(_21395_),
    .COUT(_21451_),
    .SUM(_21452_));
 sky130_fd_sc_hd__fa_1 _42727_ (.A(_01305_),
    .B(_01306_),
    .CIN(_01307_),
    .COUT(_21453_),
    .SUM(_21454_));
 sky130_fd_sc_hd__fa_1 _42728_ (.A(_01308_),
    .B(_01309_),
    .CIN(_01310_),
    .COUT(_21455_),
    .SUM(_21456_));
 sky130_fd_sc_hd__fa_1 _42729_ (.A(_21456_),
    .B(_21405_),
    .CIN(_21454_),
    .COUT(_21457_),
    .SUM(_21458_));
 sky130_fd_sc_hd__fa_1 _42730_ (.A(_21458_),
    .B(_21403_),
    .CIN(_21452_),
    .COUT(_21459_),
    .SUM(_21460_));
 sky130_fd_sc_hd__fa_1 _42731_ (.A(_21411_),
    .B(_21460_),
    .CIN(_21399_),
    .COUT(_01311_),
    .SUM(_21461_));
 sky130_fd_sc_hd__fa_1 _42732_ (.A(_21461_),
    .B(_21401_),
    .CIN(_21448_),
    .COUT(_21462_),
    .SUM(_21463_));
 sky130_fd_sc_hd__fa_1 _42733_ (.A(_01312_),
    .B(_01313_),
    .CIN(_01314_),
    .COUT(_01315_),
    .SUM(_01316_));
 sky130_fd_sc_hd__fa_1 _42734_ (.A(_01317_),
    .B(_01318_),
    .CIN(_21407_),
    .COUT(_21464_),
    .SUM(_21465_));
 sky130_fd_sc_hd__fa_1 _42735_ (.A(_21416_),
    .B(_21465_),
    .CIN(_21409_),
    .COUT(_21466_),
    .SUM(_21467_));
 sky130_fd_sc_hd__fa_1 _42736_ (.A(_01319_),
    .B(_01320_),
    .CIN(_01321_),
    .COUT(_01322_),
    .SUM(_01323_));
 sky130_fd_sc_hd__fa_1 _42737_ (.A(_01324_),
    .B(_01325_),
    .CIN(_01326_),
    .COUT(_01327_),
    .SUM(_01328_));
 sky130_fd_sc_hd__fa_1 _42738_ (.A(_01329_),
    .B(_01330_),
    .CIN(_01331_),
    .COUT(_21468_),
    .SUM(_21469_));
 sky130_fd_sc_hd__fa_1 _42739_ (.A(_01332_),
    .B(_21420_),
    .CIN(_21469_),
    .COUT(_01333_),
    .SUM(_21470_));
 sky130_fd_sc_hd__fa_1 _42740_ (.A(_21470_),
    .B(_21418_),
    .CIN(_21467_),
    .COUT(_01334_),
    .SUM(_01335_));
 sky130_fd_sc_hd__fa_1 _42741_ (.A(_01336_),
    .B(_01337_),
    .CIN(_01338_),
    .COUT(_21471_),
    .SUM(_01339_));
 sky130_fd_sc_hd__fa_1 _42742_ (.A(_01340_),
    .B(_21414_),
    .CIN(_21463_),
    .COUT(_21472_),
    .SUM(_21473_));
 sky130_fd_sc_hd__fa_1 _42743_ (.A(_01341_),
    .B(_01342_),
    .CIN(_01343_),
    .COUT(_01344_),
    .SUM(_01345_));
 sky130_fd_sc_hd__fa_1 _42744_ (.A(_01346_),
    .B(_21425_),
    .CIN(_21473_),
    .COUT(_21474_),
    .SUM(_21475_));
 sky130_fd_sc_hd__fa_1 _42745_ (.A(_01347_),
    .B(_21427_),
    .CIN(_21475_),
    .COUT(_01348_),
    .SUM(_01349_));
 sky130_fd_sc_hd__fa_1 _42746_ (.A(_01351_),
    .B(_01352_),
    .CIN(_01353_),
    .COUT(_21476_),
    .SUM(_21477_));
 sky130_fd_sc_hd__fa_1 _42747_ (.A(_01354_),
    .B(_01355_),
    .CIN(_01356_),
    .COUT(_21478_),
    .SUM(_21479_));
 sky130_fd_sc_hd__fa_1 _42748_ (.A(_21479_),
    .B(_01357_),
    .CIN(_21477_),
    .COUT(_21480_),
    .SUM(_21481_));
 sky130_fd_sc_hd__fa_1 _42749_ (.A(_01358_),
    .B(_01359_),
    .CIN(_01360_),
    .COUT(_21482_),
    .SUM(_21483_));
 sky130_fd_sc_hd__fa_1 _42750_ (.A(_21433_),
    .B(_21483_),
    .CIN(_21429_),
    .COUT(_21484_),
    .SUM(_21485_));
 sky130_fd_sc_hd__fa_1 _42751_ (.A(_21485_),
    .B(_21431_),
    .CIN(_21481_),
    .COUT(_21486_),
    .SUM(_21487_));
 sky130_fd_sc_hd__fa_1 _42752_ (.A(_01361_),
    .B(_01362_),
    .CIN(_01363_),
    .COUT(_21488_),
    .SUM(_21489_));
 sky130_fd_sc_hd__fa_1 _42753_ (.A(_01364_),
    .B(_01365_),
    .CIN(_01366_),
    .COUT(_21490_),
    .SUM(_21491_));
 sky130_fd_sc_hd__fa_1 _42754_ (.A(_21491_),
    .B(_21439_),
    .CIN(_21489_),
    .COUT(_21492_),
    .SUM(_21493_));
 sky130_fd_sc_hd__fa_1 _42755_ (.A(_21443_),
    .B(_21493_),
    .CIN(_21435_),
    .COUT(_21494_),
    .SUM(_21495_));
 sky130_fd_sc_hd__fa_1 _42756_ (.A(_21495_),
    .B(_21437_),
    .CIN(_21487_),
    .COUT(_21496_),
    .SUM(_21497_));
 sky130_fd_sc_hd__fa_1 _42757_ (.A(_01367_),
    .B(_01368_),
    .CIN(_01369_),
    .COUT(_01370_),
    .SUM(_01371_));
 sky130_fd_sc_hd__fa_1 _42758_ (.A(_21449_),
    .B(_01372_),
    .CIN(_21441_),
    .COUT(_21498_),
    .SUM(_21499_));
 sky130_fd_sc_hd__fa_1 _42759_ (.A(_01373_),
    .B(_01374_),
    .CIN(_01375_),
    .COUT(_21500_),
    .SUM(_21501_));
 sky130_fd_sc_hd__fa_1 _42760_ (.A(_01376_),
    .B(_01377_),
    .CIN(_01378_),
    .COUT(_21502_),
    .SUM(_21503_));
 sky130_fd_sc_hd__fa_1 _42761_ (.A(_21503_),
    .B(_21453_),
    .CIN(_21501_),
    .COUT(_21504_),
    .SUM(_21505_));
 sky130_fd_sc_hd__fa_1 _42762_ (.A(_21505_),
    .B(_21451_),
    .CIN(_21499_),
    .COUT(_21506_),
    .SUM(_21507_));
 sky130_fd_sc_hd__fa_1 _42763_ (.A(_21459_),
    .B(_21507_),
    .CIN(_21445_),
    .COUT(_01379_),
    .SUM(_21508_));
 sky130_fd_sc_hd__fa_1 _42764_ (.A(_21508_),
    .B(_21447_),
    .CIN(_21497_),
    .COUT(_21509_),
    .SUM(_21510_));
 sky130_fd_sc_hd__fa_1 _42765_ (.A(_01380_),
    .B(_01381_),
    .CIN(_01382_),
    .COUT(_01383_),
    .SUM(_01384_));
 sky130_fd_sc_hd__fa_1 _42766_ (.A(_01385_),
    .B(_01386_),
    .CIN(_21455_),
    .COUT(_21511_),
    .SUM(_21512_));
 sky130_fd_sc_hd__fa_1 _42767_ (.A(_21464_),
    .B(_21512_),
    .CIN(_21457_),
    .COUT(_21513_),
    .SUM(_21514_));
 sky130_fd_sc_hd__fa_1 _42768_ (.A(_01387_),
    .B(_01388_),
    .CIN(_01389_),
    .COUT(_01390_),
    .SUM(_01391_));
 sky130_fd_sc_hd__fa_1 _42769_ (.A(_01392_),
    .B(_01393_),
    .CIN(_01394_),
    .COUT(_21515_),
    .SUM(_21516_));
 sky130_fd_sc_hd__fa_1 _42770_ (.A(_21516_),
    .B(_01395_),
    .CIN(_01396_),
    .COUT(_21517_),
    .SUM(_21518_));
 sky130_fd_sc_hd__fa_1 _42771_ (.A(_01397_),
    .B(_21468_),
    .CIN(_21518_),
    .COUT(_01398_),
    .SUM(_21519_));
 sky130_fd_sc_hd__fa_1 _42772_ (.A(_21519_),
    .B(_21466_),
    .CIN(_21514_),
    .COUT(_01399_),
    .SUM(_01400_));
 sky130_fd_sc_hd__fa_1 _42773_ (.A(_01401_),
    .B(_01402_),
    .CIN(_01403_),
    .COUT(_21520_),
    .SUM(_01404_));
 sky130_fd_sc_hd__fa_1 _42774_ (.A(_01405_),
    .B(_21462_),
    .CIN(_21510_),
    .COUT(_21521_),
    .SUM(_21522_));
 sky130_fd_sc_hd__fa_1 _42775_ (.A(_01406_),
    .B(_21472_),
    .CIN(_21522_),
    .COUT(_21523_),
    .SUM(_21524_));
 sky130_fd_sc_hd__fa_1 _42776_ (.A(_01407_),
    .B(_21474_),
    .CIN(_21524_),
    .COUT(_01408_),
    .SUM(_01409_));
 sky130_fd_sc_hd__fa_1 _42777_ (.A(_01410_),
    .B(_01411_),
    .CIN(_01412_),
    .COUT(_21525_),
    .SUM(_21526_));
 sky130_fd_sc_hd__fa_1 _42778_ (.A(_01413_),
    .B(_01414_),
    .CIN(_01415_),
    .COUT(_21527_),
    .SUM(_21528_));
 sky130_fd_sc_hd__fa_1 _42779_ (.A(_21528_),
    .B(_21476_),
    .CIN(_21526_),
    .COUT(_21529_),
    .SUM(_21530_));
 sky130_fd_sc_hd__fa_1 _42780_ (.A(_01416_),
    .B(_01417_),
    .CIN(_01418_),
    .COUT(_21531_),
    .SUM(_21532_));
 sky130_fd_sc_hd__fa_1 _42781_ (.A(_21482_),
    .B(_21532_),
    .CIN(_21478_),
    .COUT(_21533_),
    .SUM(_21534_));
 sky130_fd_sc_hd__fa_1 _42782_ (.A(_21534_),
    .B(_21480_),
    .CIN(_21530_),
    .COUT(_21535_),
    .SUM(_21536_));
 sky130_fd_sc_hd__fa_1 _42783_ (.A(_01419_),
    .B(_01420_),
    .CIN(_01421_),
    .COUT(_21537_),
    .SUM(_21538_));
 sky130_fd_sc_hd__fa_1 _42784_ (.A(_01422_),
    .B(_01423_),
    .CIN(_01424_),
    .COUT(_21539_),
    .SUM(_21540_));
 sky130_fd_sc_hd__fa_1 _42785_ (.A(_21540_),
    .B(_21488_),
    .CIN(_21538_),
    .COUT(_21541_),
    .SUM(_21542_));
 sky130_fd_sc_hd__fa_1 _42786_ (.A(_21492_),
    .B(_21542_),
    .CIN(_21484_),
    .COUT(_21543_),
    .SUM(_21544_));
 sky130_fd_sc_hd__fa_1 _42787_ (.A(_21544_),
    .B(_21486_),
    .CIN(_21536_),
    .COUT(_21545_),
    .SUM(_21546_));
 sky130_fd_sc_hd__fa_1 _42788_ (.A(_01425_),
    .B(_01426_),
    .CIN(_01427_),
    .COUT(_21547_),
    .SUM(_21548_));
 sky130_fd_sc_hd__fa_1 _42789_ (.A(_01429_),
    .B(_21548_),
    .CIN(_21490_),
    .COUT(_21549_),
    .SUM(_21550_));
 sky130_fd_sc_hd__fa_1 _42790_ (.A(_01430_),
    .B(_01431_),
    .CIN(_01432_),
    .COUT(_21551_),
    .SUM(_21552_));
 sky130_fd_sc_hd__fa_1 _42791_ (.A(_01433_),
    .B(_01434_),
    .CIN(_01435_),
    .COUT(_21553_),
    .SUM(_21554_));
 sky130_fd_sc_hd__fa_1 _42792_ (.A(_21554_),
    .B(_21500_),
    .CIN(_21552_),
    .COUT(_21555_),
    .SUM(_21556_));
 sky130_fd_sc_hd__fa_1 _42793_ (.A(_21556_),
    .B(_21498_),
    .CIN(_21550_),
    .COUT(_21557_),
    .SUM(_21558_));
 sky130_fd_sc_hd__fa_1 _42794_ (.A(_21506_),
    .B(_21558_),
    .CIN(_21494_),
    .COUT(_01436_),
    .SUM(_21559_));
 sky130_fd_sc_hd__fa_1 _42795_ (.A(_21559_),
    .B(_21496_),
    .CIN(_21546_),
    .COUT(_21560_),
    .SUM(_21561_));
 sky130_fd_sc_hd__fa_1 _42796_ (.A(_01437_),
    .B(_01438_),
    .CIN(_01439_),
    .COUT(_01440_),
    .SUM(_01441_));
 sky130_fd_sc_hd__fa_1 _42797_ (.A(_01442_),
    .B(_01443_),
    .CIN(_21502_),
    .COUT(_21562_),
    .SUM(_21563_));
 sky130_fd_sc_hd__fa_1 _42798_ (.A(_21511_),
    .B(_21563_),
    .CIN(_21504_),
    .COUT(_21564_),
    .SUM(_21565_));
 sky130_fd_sc_hd__fa_1 _42799_ (.A(_01444_),
    .B(_01445_),
    .CIN(_01446_),
    .COUT(_01447_),
    .SUM(_01448_));
 sky130_fd_sc_hd__fa_1 _42800_ (.A(_01449_),
    .B(_01450_),
    .CIN(_01341_),
    .COUT(_01451_),
    .SUM(_01452_));
 sky130_fd_sc_hd__fa_1 _42801_ (.A(_01453_),
    .B(_01454_),
    .CIN(_01455_),
    .COUT(_21566_),
    .SUM(_21567_));
 sky130_fd_sc_hd__fa_1 _42802_ (.A(_21515_),
    .B(_21517_),
    .CIN(_21567_),
    .COUT(_01456_),
    .SUM(_21568_));
 sky130_fd_sc_hd__fa_1 _42803_ (.A(_21568_),
    .B(_21513_),
    .CIN(_21565_),
    .COUT(_01457_),
    .SUM(_01458_));
 sky130_fd_sc_hd__fa_1 _42804_ (.A(_01459_),
    .B(_01460_),
    .CIN(_01461_),
    .COUT(_21569_),
    .SUM(_01462_));
 sky130_fd_sc_hd__fa_1 _42805_ (.A(_01463_),
    .B(_21509_),
    .CIN(_21561_),
    .COUT(_21570_),
    .SUM(_21571_));
 sky130_fd_sc_hd__fa_1 _42806_ (.A(_01464_),
    .B(_21521_),
    .CIN(_21571_),
    .COUT(_21572_),
    .SUM(_21573_));
 sky130_fd_sc_hd__fa_1 _42807_ (.A(_01465_),
    .B(_21523_),
    .CIN(_21573_),
    .COUT(_01466_),
    .SUM(_01467_));
 sky130_fd_sc_hd__fa_1 _42808_ (.A(_01469_),
    .B(_01470_),
    .CIN(_01471_),
    .COUT(_21574_),
    .SUM(_21575_));
 sky130_fd_sc_hd__fa_1 _42809_ (.A(_01472_),
    .B(_01473_),
    .CIN(_01474_),
    .COUT(_21576_),
    .SUM(_21577_));
 sky130_fd_sc_hd__fa_1 _42810_ (.A(_21577_),
    .B(_21525_),
    .CIN(_21575_),
    .COUT(_21578_),
    .SUM(_21579_));
 sky130_fd_sc_hd__fa_1 _42811_ (.A(_01475_),
    .B(_01476_),
    .CIN(_01477_),
    .COUT(_21580_),
    .SUM(_21581_));
 sky130_fd_sc_hd__fa_1 _42812_ (.A(_21531_),
    .B(_21581_),
    .CIN(_21527_),
    .COUT(_21582_),
    .SUM(_21583_));
 sky130_fd_sc_hd__fa_1 _42813_ (.A(_21583_),
    .B(_21529_),
    .CIN(_21579_),
    .COUT(_21584_),
    .SUM(_21585_));
 sky130_fd_sc_hd__fa_1 _42814_ (.A(_01478_),
    .B(_01479_),
    .CIN(_01480_),
    .COUT(_21586_),
    .SUM(_21587_));
 sky130_fd_sc_hd__fa_1 _42815_ (.A(_01481_),
    .B(_01482_),
    .CIN(_01483_),
    .COUT(_21588_),
    .SUM(_21589_));
 sky130_fd_sc_hd__fa_1 _42816_ (.A(_21589_),
    .B(_21537_),
    .CIN(_21587_),
    .COUT(_21590_),
    .SUM(_21591_));
 sky130_fd_sc_hd__fa_1 _42817_ (.A(_21541_),
    .B(_21591_),
    .CIN(_21533_),
    .COUT(_21592_),
    .SUM(_21593_));
 sky130_fd_sc_hd__fa_1 _42818_ (.A(_21593_),
    .B(_21535_),
    .CIN(_21585_),
    .COUT(_21594_),
    .SUM(_21595_));
 sky130_fd_sc_hd__fa_1 _42819_ (.A(_01484_),
    .B(_01485_),
    .CIN(_01486_),
    .COUT(_01487_),
    .SUM(_01488_));
 sky130_fd_sc_hd__fa_1 _42820_ (.A(_21547_),
    .B(_01489_),
    .CIN(_21539_),
    .COUT(_21596_),
    .SUM(_21597_));
 sky130_fd_sc_hd__fa_1 _42821_ (.A(_01490_),
    .B(_01491_),
    .CIN(_01492_),
    .COUT(_21598_),
    .SUM(_21599_));
 sky130_fd_sc_hd__fa_1 _42822_ (.A(_01493_),
    .B(_01494_),
    .CIN(_01495_),
    .COUT(_21600_),
    .SUM(_21601_));
 sky130_fd_sc_hd__fa_1 _42823_ (.A(_21601_),
    .B(_21551_),
    .CIN(_21599_),
    .COUT(_21602_),
    .SUM(_21603_));
 sky130_fd_sc_hd__fa_1 _42824_ (.A(_21603_),
    .B(_21549_),
    .CIN(_21597_),
    .COUT(_21604_),
    .SUM(_21605_));
 sky130_fd_sc_hd__fa_1 _42825_ (.A(_21557_),
    .B(_21605_),
    .CIN(_21543_),
    .COUT(_01496_),
    .SUM(_21606_));
 sky130_fd_sc_hd__fa_1 _42826_ (.A(_21606_),
    .B(_21545_),
    .CIN(_21595_),
    .COUT(_21607_),
    .SUM(_21608_));
 sky130_fd_sc_hd__fa_1 _42827_ (.A(_01497_),
    .B(_01498_),
    .CIN(_01499_),
    .COUT(_01500_),
    .SUM(_01501_));
 sky130_fd_sc_hd__fa_1 _42828_ (.A(_01502_),
    .B(_01503_),
    .CIN(_21553_),
    .COUT(_21609_),
    .SUM(_21610_));
 sky130_fd_sc_hd__fa_1 _42829_ (.A(_21562_),
    .B(_21610_),
    .CIN(_21555_),
    .COUT(_21611_),
    .SUM(_21612_));
 sky130_fd_sc_hd__fa_1 _42830_ (.A(_01504_),
    .B(_01505_),
    .CIN(_01506_),
    .COUT(_01507_),
    .SUM(_01508_));
 sky130_fd_sc_hd__fa_1 _42831_ (.A(_01509_),
    .B(_01510_),
    .CIN(_01453_),
    .COUT(_21613_),
    .SUM(_21614_));
 sky130_fd_sc_hd__fa_1 _42832_ (.A(_01511_),
    .B(_21566_),
    .CIN(_21614_),
    .COUT(_01512_),
    .SUM(_21615_));
 sky130_fd_sc_hd__fa_1 _42833_ (.A(_21615_),
    .B(_21564_),
    .CIN(_21612_),
    .COUT(_01513_),
    .SUM(_01514_));
 sky130_fd_sc_hd__fa_1 _42834_ (.A(_01515_),
    .B(_01516_),
    .CIN(_01517_),
    .COUT(_21616_),
    .SUM(_01518_));
 sky130_fd_sc_hd__fa_1 _42835_ (.A(_01519_),
    .B(_21560_),
    .CIN(_21608_),
    .COUT(_21617_),
    .SUM(_21618_));
 sky130_fd_sc_hd__fa_1 _42836_ (.A(_01520_),
    .B(_21570_),
    .CIN(_21618_),
    .COUT(_21619_),
    .SUM(_21620_));
 sky130_fd_sc_hd__fa_1 _42837_ (.A(_01521_),
    .B(_21572_),
    .CIN(_21620_),
    .COUT(_01522_),
    .SUM(_01523_));
 sky130_fd_sc_hd__fa_1 _42838_ (.A(_01525_),
    .B(_01526_),
    .CIN(_01527_),
    .COUT(_21621_),
    .SUM(_21622_));
 sky130_fd_sc_hd__fa_1 _42839_ (.A(_01528_),
    .B(_01529_),
    .CIN(_01530_),
    .COUT(_21623_),
    .SUM(_21624_));
 sky130_fd_sc_hd__fa_1 _42840_ (.A(_21624_),
    .B(_21574_),
    .CIN(_21622_),
    .COUT(_21625_),
    .SUM(_21626_));
 sky130_fd_sc_hd__fa_1 _42841_ (.A(_01531_),
    .B(_01532_),
    .CIN(_01533_),
    .COUT(_21627_),
    .SUM(_21628_));
 sky130_fd_sc_hd__fa_1 _42842_ (.A(_21580_),
    .B(_21628_),
    .CIN(_21576_),
    .COUT(_21629_),
    .SUM(_21630_));
 sky130_fd_sc_hd__fa_1 _42843_ (.A(_21630_),
    .B(_21578_),
    .CIN(_21626_),
    .COUT(_21631_),
    .SUM(_21632_));
 sky130_fd_sc_hd__fa_1 _42844_ (.A(_01534_),
    .B(_01535_),
    .CIN(_01536_),
    .COUT(_21633_),
    .SUM(_21634_));
 sky130_fd_sc_hd__fa_1 _42845_ (.A(_01537_),
    .B(_01538_),
    .CIN(_01539_),
    .COUT(_01540_),
    .SUM(_01541_));
 sky130_fd_sc_hd__fa_1 _42846_ (.A(_01542_),
    .B(_21586_),
    .CIN(_21634_),
    .COUT(_21635_),
    .SUM(_21636_));
 sky130_fd_sc_hd__fa_1 _42847_ (.A(_21590_),
    .B(_21636_),
    .CIN(_21582_),
    .COUT(_21637_),
    .SUM(_21638_));
 sky130_fd_sc_hd__fa_1 _42848_ (.A(_21638_),
    .B(_21584_),
    .CIN(_21632_),
    .COUT(_21639_),
    .SUM(_21640_));
 sky130_fd_sc_hd__fa_1 _42849_ (.A(_01543_),
    .B(_01544_),
    .CIN(_01545_),
    .COUT(_01546_),
    .SUM(_01547_));
 sky130_fd_sc_hd__fa_1 _42850_ (.A(_01548_),
    .B(_01549_),
    .CIN(_21588_),
    .COUT(_21641_),
    .SUM(_21642_));
 sky130_fd_sc_hd__fa_1 _42851_ (.A(_01550_),
    .B(_01551_),
    .CIN(_01552_),
    .COUT(_21643_),
    .SUM(_21644_));
 sky130_fd_sc_hd__fa_1 _42852_ (.A(_01553_),
    .B(_01554_),
    .CIN(_01555_),
    .COUT(_21645_),
    .SUM(_21646_));
 sky130_fd_sc_hd__fa_1 _42853_ (.A(_21646_),
    .B(_21598_),
    .CIN(_21644_),
    .COUT(_21647_),
    .SUM(_21648_));
 sky130_fd_sc_hd__fa_1 _42854_ (.A(_21648_),
    .B(_21596_),
    .CIN(_21642_),
    .COUT(_21649_),
    .SUM(_21650_));
 sky130_fd_sc_hd__fa_1 _42855_ (.A(_21604_),
    .B(_21650_),
    .CIN(_21592_),
    .COUT(_01556_),
    .SUM(_21651_));
 sky130_fd_sc_hd__fa_1 _42856_ (.A(_21651_),
    .B(_21594_),
    .CIN(_21640_),
    .COUT(_21652_),
    .SUM(_21653_));
 sky130_fd_sc_hd__fa_1 _42857_ (.A(_01557_),
    .B(_01558_),
    .CIN(_01559_),
    .COUT(_01560_),
    .SUM(_01561_));
 sky130_fd_sc_hd__fa_1 _42858_ (.A(_01562_),
    .B(_01563_),
    .CIN(_21600_),
    .COUT(_21654_),
    .SUM(_21655_));
 sky130_fd_sc_hd__fa_1 _42859_ (.A(_21609_),
    .B(_21655_),
    .CIN(_21602_),
    .COUT(_21656_),
    .SUM(_21657_));
 sky130_fd_sc_hd__fa_1 _42860_ (.A(_01564_),
    .B(_01565_),
    .CIN(_01504_),
    .COUT(_01566_),
    .SUM(_01567_));
 sky130_fd_sc_hd__fa_1 _42861_ (.A(_01568_),
    .B(_01569_),
    .CIN(_01453_),
    .COUT(_21658_),
    .SUM(_21659_));
 sky130_fd_sc_hd__fa_1 _42862_ (.A(_21613_),
    .B(_21659_),
    .CIN(_01511_),
    .COUT(_01570_),
    .SUM(_21660_));
 sky130_fd_sc_hd__fa_1 _42863_ (.A(_21660_),
    .B(_21611_),
    .CIN(_21657_),
    .COUT(_01571_),
    .SUM(_01572_));
 sky130_fd_sc_hd__fa_1 _42864_ (.A(_01573_),
    .B(_01574_),
    .CIN(_01575_),
    .COUT(_21661_),
    .SUM(_01576_));
 sky130_fd_sc_hd__fa_1 _42865_ (.A(_01577_),
    .B(_21607_),
    .CIN(_21653_),
    .COUT(_21662_),
    .SUM(_21663_));
 sky130_fd_sc_hd__fa_1 _42866_ (.A(_01578_),
    .B(_21617_),
    .CIN(_21663_),
    .COUT(_21664_),
    .SUM(_21665_));
 sky130_fd_sc_hd__fa_1 _42867_ (.A(_01579_),
    .B(_21619_),
    .CIN(_21665_),
    .COUT(_01580_),
    .SUM(_01581_));
 sky130_fd_sc_hd__fa_1 _42868_ (.A(_01583_),
    .B(_01584_),
    .CIN(_01585_),
    .COUT(_21666_),
    .SUM(_21667_));
 sky130_fd_sc_hd__fa_1 _42869_ (.A(_01586_),
    .B(_01587_),
    .CIN(_01588_),
    .COUT(_21668_),
    .SUM(_21669_));
 sky130_fd_sc_hd__fa_1 _42870_ (.A(_21669_),
    .B(_21621_),
    .CIN(_21667_),
    .COUT(_21670_),
    .SUM(_21671_));
 sky130_fd_sc_hd__fa_1 _42871_ (.A(_01589_),
    .B(_01590_),
    .CIN(_01591_),
    .COUT(_21672_),
    .SUM(_21673_));
 sky130_fd_sc_hd__fa_1 _42872_ (.A(_21627_),
    .B(_21673_),
    .CIN(_21623_),
    .COUT(_21674_),
    .SUM(_21675_));
 sky130_fd_sc_hd__fa_1 _42873_ (.A(_21675_),
    .B(_21625_),
    .CIN(_21671_),
    .COUT(_21676_),
    .SUM(_21677_));
 sky130_fd_sc_hd__fa_1 _42874_ (.A(_01592_),
    .B(_01593_),
    .CIN(_01594_),
    .COUT(_21678_),
    .SUM(_21679_));
 sky130_fd_sc_hd__fa_1 _42875_ (.A(_01595_),
    .B(_01596_),
    .CIN(_01597_),
    .COUT(_21680_),
    .SUM(_21681_));
 sky130_fd_sc_hd__fa_1 _42876_ (.A(_21681_),
    .B(_21633_),
    .CIN(_21679_),
    .COUT(_21682_),
    .SUM(_21683_));
 sky130_fd_sc_hd__fa_1 _42877_ (.A(_21635_),
    .B(_21683_),
    .CIN(_21629_),
    .COUT(_21684_),
    .SUM(_21685_));
 sky130_fd_sc_hd__fa_1 _42878_ (.A(_21685_),
    .B(_21631_),
    .CIN(_21677_),
    .COUT(_21686_),
    .SUM(_21687_));
 sky130_fd_sc_hd__fa_1 _42879_ (.A(_01598_),
    .B(_01599_),
    .CIN(_01600_),
    .COUT(_01601_),
    .SUM(_01602_));
 sky130_fd_sc_hd__fa_1 _42880_ (.A(_01603_),
    .B(_01604_),
    .CIN(_01605_),
    .COUT(_21688_),
    .SUM(_21689_));
 sky130_fd_sc_hd__fa_1 _42881_ (.A(_01606_),
    .B(_01607_),
    .CIN(_01608_),
    .COUT(_21690_),
    .SUM(_21691_));
 sky130_fd_sc_hd__fa_1 _42882_ (.A(_01609_),
    .B(_01610_),
    .CIN(_01611_),
    .COUT(_21692_),
    .SUM(_21693_));
 sky130_fd_sc_hd__fa_1 _42883_ (.A(_21693_),
    .B(_21643_),
    .CIN(_21691_),
    .COUT(_21694_),
    .SUM(_21695_));
 sky130_fd_sc_hd__fa_1 _42884_ (.A(_21695_),
    .B(_21641_),
    .CIN(_21689_),
    .COUT(_21696_),
    .SUM(_21697_));
 sky130_fd_sc_hd__fa_1 _42885_ (.A(_21649_),
    .B(_21697_),
    .CIN(_21637_),
    .COUT(_01612_),
    .SUM(_21698_));
 sky130_fd_sc_hd__fa_1 _42886_ (.A(_21698_),
    .B(_21639_),
    .CIN(_21687_),
    .COUT(_21699_),
    .SUM(_21700_));
 sky130_fd_sc_hd__fa_1 _42887_ (.A(_01613_),
    .B(_01614_),
    .CIN(_01615_),
    .COUT(_01616_),
    .SUM(_01617_));
 sky130_fd_sc_hd__fa_1 _42888_ (.A(_01618_),
    .B(_01619_),
    .CIN(_21645_),
    .COUT(_21701_),
    .SUM(_21702_));
 sky130_fd_sc_hd__fa_1 _42889_ (.A(_21654_),
    .B(_21702_),
    .CIN(_21647_),
    .COUT(_21703_),
    .SUM(_21704_));
 sky130_fd_sc_hd__fa_1 _42890_ (.A(_01620_),
    .B(_01621_),
    .CIN(_01622_),
    .COUT(_21705_),
    .SUM(_21706_));
 sky130_fd_sc_hd__fa_1 _42891_ (.A(_01623_),
    .B(_21706_),
    .CIN(_01453_),
    .COUT(_21707_),
    .SUM(_21708_));
 sky130_fd_sc_hd__fa_1 _42892_ (.A(_21658_),
    .B(_21708_),
    .CIN(_01511_),
    .COUT(_01624_),
    .SUM(_21709_));
 sky130_fd_sc_hd__fa_1 _42893_ (.A(_21709_),
    .B(_21656_),
    .CIN(_21704_),
    .COUT(_01625_),
    .SUM(_01626_));
 sky130_fd_sc_hd__fa_1 _42894_ (.A(_01627_),
    .B(_01628_),
    .CIN(_01629_),
    .COUT(_21710_),
    .SUM(_01630_));
 sky130_fd_sc_hd__fa_1 _42895_ (.A(_01631_),
    .B(_21652_),
    .CIN(_21700_),
    .COUT(_21711_),
    .SUM(_21712_));
 sky130_fd_sc_hd__fa_1 _42896_ (.A(_01632_),
    .B(_21662_),
    .CIN(_21712_),
    .COUT(_21713_),
    .SUM(_21714_));
 sky130_fd_sc_hd__fa_1 _42897_ (.A(_01633_),
    .B(_21664_),
    .CIN(_21714_),
    .COUT(_01634_),
    .SUM(_01635_));
 sky130_fd_sc_hd__fa_1 _42898_ (.A(_01637_),
    .B(_01638_),
    .CIN(_01639_),
    .COUT(_21715_),
    .SUM(_21716_));
 sky130_fd_sc_hd__fa_1 _42899_ (.A(_01640_),
    .B(_01641_),
    .CIN(_01642_),
    .COUT(_21717_),
    .SUM(_21718_));
 sky130_fd_sc_hd__fa_1 _42900_ (.A(_21718_),
    .B(_21666_),
    .CIN(_21716_),
    .COUT(_21719_),
    .SUM(_21720_));
 sky130_fd_sc_hd__fa_1 _42901_ (.A(_01643_),
    .B(_01644_),
    .CIN(_01645_),
    .COUT(_21721_),
    .SUM(_21722_));
 sky130_fd_sc_hd__fa_1 _42902_ (.A(_21672_),
    .B(_21722_),
    .CIN(_21668_),
    .COUT(_21723_),
    .SUM(_21724_));
 sky130_fd_sc_hd__fa_1 _42903_ (.A(_21724_),
    .B(_21670_),
    .CIN(_21720_),
    .COUT(_21725_),
    .SUM(_21726_));
 sky130_fd_sc_hd__fa_1 _42904_ (.A(_01646_),
    .B(_01647_),
    .CIN(_01648_),
    .COUT(_21727_),
    .SUM(_21728_));
 sky130_fd_sc_hd__fa_1 _42905_ (.A(_01649_),
    .B(_01650_),
    .CIN(_01651_),
    .COUT(_21729_),
    .SUM(_21730_));
 sky130_fd_sc_hd__fa_1 _42906_ (.A(_21730_),
    .B(_21678_),
    .CIN(_21728_),
    .COUT(_21731_),
    .SUM(_21732_));
 sky130_fd_sc_hd__fa_1 _42907_ (.A(_21682_),
    .B(_21732_),
    .CIN(_21674_),
    .COUT(_21733_),
    .SUM(_21734_));
 sky130_fd_sc_hd__fa_1 _42908_ (.A(_21734_),
    .B(_21676_),
    .CIN(_21726_),
    .COUT(_21735_),
    .SUM(_21736_));
 sky130_fd_sc_hd__fa_1 _42909_ (.A(_01652_),
    .B(_01653_),
    .CIN(_01654_),
    .COUT(_01655_),
    .SUM(_01656_));
 sky130_fd_sc_hd__fa_1 _42910_ (.A(_01657_),
    .B(_01658_),
    .CIN(_21680_),
    .COUT(_21737_),
    .SUM(_21738_));
 sky130_fd_sc_hd__fa_1 _42911_ (.A(_01659_),
    .B(_01660_),
    .CIN(_01661_),
    .COUT(_21739_),
    .SUM(_21740_));
 sky130_fd_sc_hd__fa_1 _42912_ (.A(_01662_),
    .B(_01663_),
    .CIN(_01664_),
    .COUT(_21741_),
    .SUM(_21742_));
 sky130_fd_sc_hd__fa_1 _42913_ (.A(_21742_),
    .B(_21690_),
    .CIN(_21740_),
    .COUT(_21743_),
    .SUM(_21744_));
 sky130_fd_sc_hd__fa_1 _42914_ (.A(_21744_),
    .B(_21688_),
    .CIN(_21738_),
    .COUT(_21745_),
    .SUM(_21746_));
 sky130_fd_sc_hd__fa_1 _42915_ (.A(_21696_),
    .B(_21746_),
    .CIN(_21684_),
    .COUT(_01665_),
    .SUM(_21747_));
 sky130_fd_sc_hd__fa_1 _42916_ (.A(_21747_),
    .B(_21686_),
    .CIN(_21736_),
    .COUT(_21748_),
    .SUM(_21749_));
 sky130_fd_sc_hd__fa_1 _42917_ (.A(_01666_),
    .B(_01667_),
    .CIN(_01668_),
    .COUT(_01669_),
    .SUM(_01670_));
 sky130_fd_sc_hd__fa_1 _42918_ (.A(_01671_),
    .B(_01672_),
    .CIN(_21692_),
    .COUT(_21750_),
    .SUM(_21751_));
 sky130_fd_sc_hd__fa_1 _42919_ (.A(_21701_),
    .B(_21751_),
    .CIN(_21694_),
    .COUT(_21752_),
    .SUM(_21753_));
 sky130_fd_sc_hd__fa_1 _42920_ (.A(_21705_),
    .B(_21706_),
    .CIN(_01453_),
    .COUT(_01673_),
    .SUM(_01674_));
 sky130_fd_sc_hd__fa_1 _42921_ (.A(_21707_),
    .B(_01674_),
    .CIN(_01511_),
    .COUT(_01675_),
    .SUM(_21754_));
 sky130_fd_sc_hd__fa_1 _42922_ (.A(_21754_),
    .B(_21703_),
    .CIN(_21753_),
    .COUT(_01677_),
    .SUM(_01678_));
 sky130_fd_sc_hd__fa_1 _42923_ (.A(_01679_),
    .B(_01680_),
    .CIN(_01681_),
    .COUT(_21755_),
    .SUM(_01682_));
 sky130_fd_sc_hd__fa_1 _42924_ (.A(_01683_),
    .B(_21699_),
    .CIN(_21749_),
    .COUT(_21756_),
    .SUM(_21757_));
 sky130_fd_sc_hd__fa_1 _42925_ (.A(_01684_),
    .B(_21711_),
    .CIN(_21757_),
    .COUT(_21758_),
    .SUM(_21759_));
 sky130_fd_sc_hd__fa_1 _42926_ (.A(_01685_),
    .B(_21713_),
    .CIN(_21759_),
    .COUT(_01686_),
    .SUM(_01687_));
 sky130_fd_sc_hd__fa_1 _42927_ (.A(_01689_),
    .B(_01690_),
    .CIN(_01691_),
    .COUT(_21760_),
    .SUM(_21761_));
 sky130_fd_sc_hd__fa_1 _42928_ (.A(_01692_),
    .B(_01693_),
    .CIN(_01694_),
    .COUT(_21762_),
    .SUM(_21763_));
 sky130_fd_sc_hd__fa_1 _42929_ (.A(_21763_),
    .B(_21715_),
    .CIN(_21761_),
    .COUT(_21764_),
    .SUM(_21765_));
 sky130_fd_sc_hd__fa_1 _42930_ (.A(_01695_),
    .B(_01696_),
    .CIN(_01697_),
    .COUT(_21766_),
    .SUM(_21767_));
 sky130_fd_sc_hd__fa_1 _42931_ (.A(_21721_),
    .B(_21767_),
    .CIN(_21717_),
    .COUT(_21768_),
    .SUM(_21769_));
 sky130_fd_sc_hd__fa_1 _42932_ (.A(_21769_),
    .B(_21719_),
    .CIN(_21765_),
    .COUT(_21770_),
    .SUM(_21771_));
 sky130_fd_sc_hd__fa_1 _42933_ (.A(_01698_),
    .B(_01699_),
    .CIN(_01700_),
    .COUT(_21772_),
    .SUM(_21773_));
 sky130_fd_sc_hd__fa_1 _42934_ (.A(_01701_),
    .B(_01702_),
    .CIN(_01703_),
    .COUT(_21774_),
    .SUM(_21775_));
 sky130_fd_sc_hd__fa_1 _42935_ (.A(_21775_),
    .B(_21727_),
    .CIN(_21773_),
    .COUT(_21776_),
    .SUM(_21777_));
 sky130_fd_sc_hd__fa_1 _42936_ (.A(_21731_),
    .B(_21777_),
    .CIN(_21723_),
    .COUT(_21778_),
    .SUM(_21779_));
 sky130_fd_sc_hd__fa_1 _42937_ (.A(_21779_),
    .B(_21725_),
    .CIN(_21771_),
    .COUT(_21780_),
    .SUM(_21781_));
 sky130_fd_sc_hd__fa_1 _42938_ (.A(_01704_),
    .B(_01705_),
    .CIN(_01706_),
    .COUT(_01707_),
    .SUM(_01708_));
 sky130_fd_sc_hd__fa_1 _42939_ (.A(_01709_),
    .B(_01710_),
    .CIN(_21729_),
    .COUT(_21782_),
    .SUM(_21783_));
 sky130_fd_sc_hd__fa_1 _42940_ (.A(_01711_),
    .B(_01712_),
    .CIN(_01713_),
    .COUT(_21784_),
    .SUM(_21785_));
 sky130_fd_sc_hd__fa_1 _42941_ (.A(_01714_),
    .B(_01715_),
    .CIN(_01716_),
    .COUT(_21786_),
    .SUM(_21787_));
 sky130_fd_sc_hd__fa_1 _42942_ (.A(_21787_),
    .B(_21739_),
    .CIN(_21785_),
    .COUT(_01717_),
    .SUM(_21788_));
 sky130_fd_sc_hd__fa_1 _42943_ (.A(_21788_),
    .B(_21737_),
    .CIN(_21783_),
    .COUT(_21789_),
    .SUM(_21790_));
 sky130_fd_sc_hd__fa_1 _42944_ (.A(_21745_),
    .B(_21790_),
    .CIN(_21733_),
    .COUT(_21791_),
    .SUM(_21792_));
 sky130_fd_sc_hd__fa_1 _42945_ (.A(_21792_),
    .B(_21735_),
    .CIN(_21781_),
    .COUT(_21793_),
    .SUM(_21794_));
 sky130_fd_sc_hd__fa_1 _42946_ (.A(_01718_),
    .B(_01719_),
    .CIN(_01720_),
    .COUT(_21795_),
    .SUM(_21796_));
 sky130_fd_sc_hd__fa_1 _42947_ (.A(_01721_),
    .B(_21796_),
    .CIN(_21741_),
    .COUT(_01722_),
    .SUM(_21797_));
 sky130_fd_sc_hd__fa_1 _42948_ (.A(_21750_),
    .B(_21797_),
    .CIN(_21743_),
    .COUT(_01723_),
    .SUM(_21798_));
 sky130_fd_sc_hd__fa_1 _42949_ (.A(_01724_),
    .B(_01676_),
    .CIN(_01451_),
    .COUT(_01725_),
    .SUM(_01726_));
 sky130_fd_sc_hd__fa_1 _42950_ (.A(_01727_),
    .B(_21752_),
    .CIN(_21798_),
    .COUT(_21799_),
    .SUM(_01728_));
 sky130_fd_sc_hd__fa_1 _42951_ (.A(_01729_),
    .B(_01730_),
    .CIN(_01731_),
    .COUT(_21800_),
    .SUM(_01732_));
 sky130_fd_sc_hd__fa_1 _42952_ (.A(_01733_),
    .B(_21748_),
    .CIN(_21794_),
    .COUT(_21801_),
    .SUM(_21802_));
 sky130_fd_sc_hd__fa_1 _42953_ (.A(_01734_),
    .B(_21756_),
    .CIN(_21802_),
    .COUT(_21803_),
    .SUM(_21804_));
 sky130_fd_sc_hd__fa_1 _42954_ (.A(_01735_),
    .B(_21758_),
    .CIN(_21804_),
    .COUT(_01736_),
    .SUM(_01737_));
 sky130_fd_sc_hd__fa_1 _42955_ (.A(_01739_),
    .B(_01740_),
    .CIN(_01741_),
    .COUT(_21805_),
    .SUM(_21806_));
 sky130_fd_sc_hd__fa_1 _42956_ (.A(_01742_),
    .B(_01743_),
    .CIN(_01744_),
    .COUT(_21807_),
    .SUM(_21808_));
 sky130_fd_sc_hd__fa_1 _42957_ (.A(_21808_),
    .B(_21760_),
    .CIN(_21806_),
    .COUT(_21809_),
    .SUM(_21810_));
 sky130_fd_sc_hd__fa_1 _42958_ (.A(_01745_),
    .B(_01746_),
    .CIN(_01747_),
    .COUT(_21811_),
    .SUM(_21812_));
 sky130_fd_sc_hd__fa_1 _42959_ (.A(_21766_),
    .B(_21812_),
    .CIN(_21762_),
    .COUT(_21813_),
    .SUM(_21814_));
 sky130_fd_sc_hd__fa_1 _42960_ (.A(_21814_),
    .B(_21764_),
    .CIN(_21810_),
    .COUT(_21815_),
    .SUM(_21816_));
 sky130_fd_sc_hd__fa_1 _42961_ (.A(_01748_),
    .B(_01749_),
    .CIN(_01750_),
    .COUT(_21817_),
    .SUM(_21818_));
 sky130_fd_sc_hd__fa_1 _42962_ (.A(_01751_),
    .B(_01752_),
    .CIN(_01753_),
    .COUT(_21819_),
    .SUM(_21820_));
 sky130_fd_sc_hd__fa_1 _42963_ (.A(_21820_),
    .B(_21772_),
    .CIN(_21818_),
    .COUT(_21821_),
    .SUM(_21822_));
 sky130_fd_sc_hd__fa_1 _42964_ (.A(_21776_),
    .B(_21822_),
    .CIN(_21768_),
    .COUT(_21823_),
    .SUM(_21824_));
 sky130_fd_sc_hd__fa_1 _42965_ (.A(_21824_),
    .B(_21770_),
    .CIN(_21816_),
    .COUT(_21825_),
    .SUM(_21826_));
 sky130_fd_sc_hd__fa_1 _42966_ (.A(_01754_),
    .B(_01755_),
    .CIN(_01756_),
    .COUT(_01757_),
    .SUM(_01758_));
 sky130_fd_sc_hd__fa_1 _42967_ (.A(_01759_),
    .B(_01760_),
    .CIN(_21774_),
    .COUT(_21827_),
    .SUM(_21828_));
 sky130_fd_sc_hd__fa_1 _42968_ (.A(_01761_),
    .B(_01762_),
    .CIN(_01763_),
    .COUT(_21829_),
    .SUM(_21830_));
 sky130_fd_sc_hd__fa_1 _42969_ (.A(_01764_),
    .B(_01765_),
    .CIN(_01766_),
    .COUT(_21831_),
    .SUM(_21832_));
 sky130_fd_sc_hd__fa_1 _42970_ (.A(_21832_),
    .B(_21784_),
    .CIN(_21830_),
    .COUT(_01767_),
    .SUM(_21833_));
 sky130_fd_sc_hd__fa_1 _42971_ (.A(_21833_),
    .B(_21782_),
    .CIN(_21828_),
    .COUT(_21834_),
    .SUM(_21835_));
 sky130_fd_sc_hd__fa_1 _42972_ (.A(_21789_),
    .B(_21835_),
    .CIN(_21778_),
    .COUT(_21836_),
    .SUM(_21837_));
 sky130_fd_sc_hd__fa_1 _42973_ (.A(_21837_),
    .B(_21780_),
    .CIN(_21826_),
    .COUT(_21838_),
    .SUM(_21839_));
 sky130_fd_sc_hd__fa_1 _42974_ (.A(_01768_),
    .B(_01769_),
    .CIN(_01666_),
    .COUT(_01770_),
    .SUM(_01771_));
 sky130_fd_sc_hd__fa_1 _42975_ (.A(_21795_),
    .B(_01772_),
    .CIN(_21786_),
    .COUT(_01773_),
    .SUM(_01774_));
 sky130_fd_sc_hd__fa_1 _42976_ (.A(_01775_),
    .B(_01776_),
    .CIN(_01777_),
    .COUT(_21840_),
    .SUM(_21841_));
 sky130_fd_sc_hd__fa_1 _42977_ (.A(_01778_),
    .B(_21841_),
    .CIN(_01726_),
    .COUT(_01779_),
    .SUM(_01780_));
 sky130_fd_sc_hd__fa_1 _42978_ (.A(_21799_),
    .B(_01781_),
    .CIN(_21791_),
    .COUT(_01782_),
    .SUM(_21842_));
 sky130_fd_sc_hd__fa_1 _42979_ (.A(_21842_),
    .B(_21793_),
    .CIN(_21839_),
    .COUT(_21843_),
    .SUM(_21844_));
 sky130_fd_sc_hd__fa_1 _42980_ (.A(_01783_),
    .B(_21801_),
    .CIN(_21844_),
    .COUT(_21845_),
    .SUM(_21846_));
 sky130_fd_sc_hd__fa_1 _42981_ (.A(_01784_),
    .B(_21803_),
    .CIN(_21846_),
    .COUT(_01785_),
    .SUM(_01786_));
 sky130_fd_sc_hd__fa_1 _42982_ (.A(_01788_),
    .B(_01789_),
    .CIN(_01790_),
    .COUT(_21847_),
    .SUM(_21848_));
 sky130_fd_sc_hd__fa_1 _42983_ (.A(_01791_),
    .B(_01792_),
    .CIN(_01793_),
    .COUT(_21849_),
    .SUM(_21850_));
 sky130_fd_sc_hd__fa_1 _42984_ (.A(_21850_),
    .B(_21805_),
    .CIN(_21848_),
    .COUT(_21851_),
    .SUM(_21852_));
 sky130_fd_sc_hd__fa_1 _42985_ (.A(_01794_),
    .B(_01795_),
    .CIN(_01796_),
    .COUT(_21853_),
    .SUM(_21854_));
 sky130_fd_sc_hd__fa_1 _42986_ (.A(_21811_),
    .B(_21854_),
    .CIN(_21807_),
    .COUT(_21855_),
    .SUM(_21856_));
 sky130_fd_sc_hd__fa_1 _42987_ (.A(_21856_),
    .B(_21809_),
    .CIN(_21852_),
    .COUT(_21857_),
    .SUM(_21858_));
 sky130_fd_sc_hd__fa_1 _42988_ (.A(_01797_),
    .B(_01798_),
    .CIN(_01799_),
    .COUT(_21859_),
    .SUM(_21860_));
 sky130_fd_sc_hd__fa_1 _42989_ (.A(_01800_),
    .B(_01801_),
    .CIN(_01802_),
    .COUT(_21861_),
    .SUM(_21862_));
 sky130_fd_sc_hd__fa_1 _42990_ (.A(_21862_),
    .B(_21817_),
    .CIN(_21860_),
    .COUT(_21863_),
    .SUM(_21864_));
 sky130_fd_sc_hd__fa_1 _42991_ (.A(_21821_),
    .B(_21864_),
    .CIN(_21813_),
    .COUT(_21865_),
    .SUM(_21866_));
 sky130_fd_sc_hd__fa_1 _42992_ (.A(_21866_),
    .B(_21815_),
    .CIN(_21858_),
    .COUT(_21867_),
    .SUM(_21868_));
 sky130_fd_sc_hd__fa_1 _42993_ (.A(_01803_),
    .B(_01804_),
    .CIN(_01805_),
    .COUT(_01806_),
    .SUM(_01807_));
 sky130_fd_sc_hd__fa_1 _42994_ (.A(_01808_),
    .B(_01809_),
    .CIN(_21819_),
    .COUT(_21869_),
    .SUM(_21870_));
 sky130_fd_sc_hd__fa_1 _42995_ (.A(_01810_),
    .B(_01811_),
    .CIN(_01812_),
    .COUT(_21871_),
    .SUM(_21872_));
 sky130_fd_sc_hd__fa_1 _42996_ (.A(_01813_),
    .B(_01814_),
    .CIN(_01815_),
    .COUT(_01816_),
    .SUM(_01817_));
 sky130_fd_sc_hd__fa_1 _42997_ (.A(_01818_),
    .B(_21829_),
    .CIN(_21872_),
    .COUT(_01819_),
    .SUM(_21873_));
 sky130_fd_sc_hd__fa_1 _42998_ (.A(_21873_),
    .B(_21827_),
    .CIN(_21870_),
    .COUT(_21874_),
    .SUM(_21875_));
 sky130_fd_sc_hd__fa_1 _42999_ (.A(_21834_),
    .B(_21875_),
    .CIN(_21823_),
    .COUT(_21876_),
    .SUM(_21877_));
 sky130_fd_sc_hd__fa_1 _43000_ (.A(_21877_),
    .B(_21825_),
    .CIN(_21868_),
    .COUT(_21878_),
    .SUM(_21879_));
 sky130_fd_sc_hd__fa_1 _43001_ (.A(_01820_),
    .B(_21831_),
    .CIN(_01772_),
    .COUT(_01821_),
    .SUM(_01822_));
 sky130_fd_sc_hd__fa_1 _43002_ (.A(_01823_),
    .B(_01824_),
    .CIN(_01825_),
    .COUT(_21880_),
    .SUM(_21881_));
 sky130_fd_sc_hd__fa_1 _43003_ (.A(_21840_),
    .B(_21881_),
    .CIN(_01726_),
    .COUT(_01826_),
    .SUM(_01827_));
 sky130_fd_sc_hd__fa_1 _43004_ (.A(_01828_),
    .B(_01829_),
    .CIN(_21836_),
    .COUT(_01830_),
    .SUM(_21882_));
 sky130_fd_sc_hd__fa_1 _43005_ (.A(_21882_),
    .B(_21838_),
    .CIN(_21879_),
    .COUT(_21883_),
    .SUM(_21884_));
 sky130_fd_sc_hd__fa_1 _43006_ (.A(_01831_),
    .B(_21843_),
    .CIN(_21884_),
    .COUT(_21885_),
    .SUM(_21886_));
 sky130_fd_sc_hd__fa_1 _43007_ (.A(_01832_),
    .B(_21845_),
    .CIN(_21886_),
    .COUT(_01833_),
    .SUM(_01834_));
 sky130_fd_sc_hd__fa_1 _43008_ (.A(_01836_),
    .B(_01837_),
    .CIN(_01838_),
    .COUT(_21887_),
    .SUM(_21888_));
 sky130_fd_sc_hd__fa_1 _43009_ (.A(_01839_),
    .B(_01840_),
    .CIN(_01841_),
    .COUT(_21889_),
    .SUM(_21890_));
 sky130_fd_sc_hd__fa_1 _43010_ (.A(_21890_),
    .B(_21847_),
    .CIN(_21888_),
    .COUT(_21891_),
    .SUM(_21892_));
 sky130_fd_sc_hd__fa_1 _43011_ (.A(_01842_),
    .B(_01843_),
    .CIN(_01844_),
    .COUT(_01845_),
    .SUM(_01846_));
 sky130_fd_sc_hd__fa_1 _43012_ (.A(_21853_),
    .B(_01847_),
    .CIN(_21849_),
    .COUT(_21893_),
    .SUM(_21894_));
 sky130_fd_sc_hd__fa_1 _43013_ (.A(_21894_),
    .B(_21851_),
    .CIN(_21892_),
    .COUT(_21895_),
    .SUM(_21896_));
 sky130_fd_sc_hd__fa_1 _43014_ (.A(_01848_),
    .B(_01849_),
    .CIN(_01850_),
    .COUT(_01851_),
    .SUM(_01852_));
 sky130_fd_sc_hd__fa_1 _43015_ (.A(_01853_),
    .B(_01854_),
    .CIN(_01855_),
    .COUT(_21897_),
    .SUM(_21898_));
 sky130_fd_sc_hd__fa_1 _43016_ (.A(_21898_),
    .B(_21859_),
    .CIN(_01856_),
    .COUT(_21899_),
    .SUM(_21900_));
 sky130_fd_sc_hd__fa_1 _43017_ (.A(_21863_),
    .B(_21900_),
    .CIN(_21855_),
    .COUT(_21901_),
    .SUM(_21902_));
 sky130_fd_sc_hd__fa_1 _43018_ (.A(_21902_),
    .B(_21857_),
    .CIN(_21896_),
    .COUT(_21903_),
    .SUM(_21904_));
 sky130_fd_sc_hd__fa_1 _43019_ (.A(_01857_),
    .B(_01858_),
    .CIN(_01859_),
    .COUT(_01860_),
    .SUM(_01861_));
 sky130_fd_sc_hd__fa_1 _43020_ (.A(_01862_),
    .B(_01863_),
    .CIN(_21861_),
    .COUT(_21905_),
    .SUM(_21906_));
 sky130_fd_sc_hd__fa_1 _43021_ (.A(_01864_),
    .B(_01865_),
    .CIN(_01866_),
    .COUT(_21907_),
    .SUM(_21908_));
 sky130_fd_sc_hd__fa_1 _43022_ (.A(_01867_),
    .B(_01868_),
    .CIN(_01813_),
    .COUT(_01869_),
    .SUM(_01870_));
 sky130_fd_sc_hd__fa_1 _43023_ (.A(_01871_),
    .B(_21871_),
    .CIN(_21908_),
    .COUT(_01872_),
    .SUM(_21909_));
 sky130_fd_sc_hd__fa_1 _43024_ (.A(_21909_),
    .B(_21869_),
    .CIN(_21906_),
    .COUT(_21910_),
    .SUM(_21911_));
 sky130_fd_sc_hd__fa_1 _43025_ (.A(_21874_),
    .B(_21911_),
    .CIN(_21865_),
    .COUT(_21912_),
    .SUM(_21913_));
 sky130_fd_sc_hd__fa_1 _43026_ (.A(_21913_),
    .B(_21867_),
    .CIN(_21904_),
    .COUT(_21914_),
    .SUM(_21915_));
 sky130_fd_sc_hd__fa_1 _43027_ (.A(_01873_),
    .B(_01820_),
    .CIN(_01772_),
    .COUT(_01874_),
    .SUM(_01875_));
 sky130_fd_sc_hd__fa_1 _43028_ (.A(_01876_),
    .B(_01877_),
    .CIN(_01878_),
    .COUT(_21916_),
    .SUM(_21917_));
 sky130_fd_sc_hd__fa_1 _43029_ (.A(_21880_),
    .B(_21917_),
    .CIN(_01726_),
    .COUT(_01879_),
    .SUM(_01880_));
 sky130_fd_sc_hd__fa_1 _43030_ (.A(_01881_),
    .B(_01882_),
    .CIN(_21876_),
    .COUT(_01883_),
    .SUM(_21918_));
 sky130_fd_sc_hd__fa_1 _43031_ (.A(_21918_),
    .B(_21878_),
    .CIN(_21915_),
    .COUT(_21919_),
    .SUM(_21920_));
 sky130_fd_sc_hd__fa_1 _43032_ (.A(_01884_),
    .B(_21883_),
    .CIN(_21920_),
    .COUT(_21921_),
    .SUM(_21922_));
 sky130_fd_sc_hd__fa_1 _43033_ (.A(_01885_),
    .B(_21885_),
    .CIN(_21922_),
    .COUT(_01886_),
    .SUM(_01887_));
 sky130_fd_sc_hd__fa_1 _43034_ (.A(_01889_),
    .B(_01890_),
    .CIN(_01891_),
    .COUT(_21923_),
    .SUM(_21924_));
 sky130_fd_sc_hd__fa_1 _43035_ (.A(_01892_),
    .B(_01893_),
    .CIN(_01894_),
    .COUT(_21925_),
    .SUM(_21926_));
 sky130_fd_sc_hd__fa_1 _43036_ (.A(_21926_),
    .B(_21887_),
    .CIN(_21924_),
    .COUT(_21927_),
    .SUM(_21928_));
 sky130_fd_sc_hd__fa_1 _43037_ (.A(_01895_),
    .B(_01896_),
    .CIN(_01897_),
    .COUT(_01898_),
    .SUM(_01899_));
 sky130_fd_sc_hd__fa_1 _43038_ (.A(_01900_),
    .B(_01901_),
    .CIN(_21889_),
    .COUT(_21929_),
    .SUM(_21930_));
 sky130_fd_sc_hd__fa_1 _43039_ (.A(_21930_),
    .B(_21891_),
    .CIN(_21928_),
    .COUT(_21931_),
    .SUM(_21932_));
 sky130_fd_sc_hd__fa_1 _43040_ (.A(_01902_),
    .B(_01903_),
    .CIN(_01904_),
    .COUT(_01905_),
    .SUM(_01906_));
 sky130_fd_sc_hd__fa_1 _43041_ (.A(_01907_),
    .B(_01908_),
    .CIN(_01909_),
    .COUT(_21933_),
    .SUM(_21934_));
 sky130_fd_sc_hd__fa_1 _43042_ (.A(_21934_),
    .B(_01910_),
    .CIN(_01911_),
    .COUT(_21935_),
    .SUM(_21936_));
 sky130_fd_sc_hd__fa_1 _43043_ (.A(_21899_),
    .B(_21936_),
    .CIN(_21893_),
    .COUT(_21937_),
    .SUM(_21938_));
 sky130_fd_sc_hd__fa_1 _43044_ (.A(_21938_),
    .B(_21895_),
    .CIN(_21932_),
    .COUT(_21939_),
    .SUM(_21940_));
 sky130_fd_sc_hd__fa_1 _43045_ (.A(_01912_),
    .B(_01913_),
    .CIN(_01914_),
    .COUT(_21941_),
    .SUM(_21942_));
 sky130_fd_sc_hd__fa_1 _43046_ (.A(_01915_),
    .B(_21942_),
    .CIN(_21897_),
    .COUT(_21943_),
    .SUM(_21944_));
 sky130_fd_sc_hd__fa_1 _43047_ (.A(_01916_),
    .B(_01917_),
    .CIN(_01918_),
    .COUT(_01919_),
    .SUM(_01920_));
 sky130_fd_sc_hd__fa_1 _43048_ (.A(_01921_),
    .B(_01867_),
    .CIN(_01813_),
    .COUT(_21945_),
    .SUM(_01922_));
 sky130_fd_sc_hd__fa_1 _43049_ (.A(_01923_),
    .B(_21907_),
    .CIN(_01924_),
    .COUT(_01925_),
    .SUM(_21946_));
 sky130_fd_sc_hd__fa_1 _43050_ (.A(_21946_),
    .B(_21905_),
    .CIN(_21944_),
    .COUT(_21947_),
    .SUM(_21948_));
 sky130_fd_sc_hd__fa_1 _43051_ (.A(_21910_),
    .B(_21948_),
    .CIN(_21901_),
    .COUT(_21949_),
    .SUM(_21950_));
 sky130_fd_sc_hd__fa_1 _43052_ (.A(_21950_),
    .B(_21903_),
    .CIN(_21940_),
    .COUT(_21951_),
    .SUM(_21952_));
 sky130_fd_sc_hd__fa_1 _43053_ (.A(_01926_),
    .B(_01820_),
    .CIN(_01772_),
    .COUT(_01927_),
    .SUM(_01928_));
 sky130_fd_sc_hd__fa_1 _43054_ (.A(_01929_),
    .B(_01930_),
    .CIN(_01931_),
    .COUT(_21953_),
    .SUM(_21954_));
 sky130_fd_sc_hd__fa_1 _43055_ (.A(_21916_),
    .B(_21954_),
    .CIN(_01726_),
    .COUT(_01932_),
    .SUM(_01933_));
 sky130_fd_sc_hd__fa_1 _43056_ (.A(_01934_),
    .B(_01935_),
    .CIN(_21912_),
    .COUT(_01936_),
    .SUM(_21955_));
 sky130_fd_sc_hd__fa_1 _43057_ (.A(_21955_),
    .B(_21914_),
    .CIN(_21952_),
    .COUT(_21956_),
    .SUM(_21957_));
 sky130_fd_sc_hd__fa_1 _43058_ (.A(_01937_),
    .B(_21919_),
    .CIN(_21957_),
    .COUT(_21958_),
    .SUM(_21959_));
 sky130_fd_sc_hd__fa_1 _43059_ (.A(_01938_),
    .B(_21921_),
    .CIN(_21959_),
    .COUT(_01939_),
    .SUM(_01940_));
 sky130_fd_sc_hd__fa_1 _43060_ (.A(_01942_),
    .B(_01943_),
    .CIN(_01944_),
    .COUT(_21960_),
    .SUM(_21961_));
 sky130_fd_sc_hd__fa_1 _43061_ (.A(_01945_),
    .B(_01946_),
    .CIN(_01947_),
    .COUT(_21962_),
    .SUM(_21963_));
 sky130_fd_sc_hd__fa_1 _43062_ (.A(_21963_),
    .B(_21923_),
    .CIN(_21961_),
    .COUT(_21964_),
    .SUM(_21965_));
 sky130_fd_sc_hd__fa_1 _43063_ (.A(_01948_),
    .B(_01949_),
    .CIN(_01950_),
    .COUT(_01951_),
    .SUM(_01952_));
 sky130_fd_sc_hd__fa_1 _43064_ (.A(_01953_),
    .B(_01954_),
    .CIN(_21925_),
    .COUT(_21966_),
    .SUM(_21967_));
 sky130_fd_sc_hd__fa_1 _43065_ (.A(_21967_),
    .B(_21927_),
    .CIN(_21965_),
    .COUT(_21968_),
    .SUM(_21969_));
 sky130_fd_sc_hd__fa_1 _43066_ (.A(_01955_),
    .B(_01956_),
    .CIN(_01957_),
    .COUT(_21970_),
    .SUM(_21971_));
 sky130_fd_sc_hd__fa_1 _43067_ (.A(_01959_),
    .B(_01960_),
    .CIN(_01961_),
    .COUT(_21972_),
    .SUM(_21973_));
 sky130_fd_sc_hd__fa_1 _43068_ (.A(_21973_),
    .B(_01962_),
    .CIN(_21971_),
    .COUT(_21974_),
    .SUM(_21975_));
 sky130_fd_sc_hd__fa_1 _43069_ (.A(_21935_),
    .B(_21975_),
    .CIN(_21929_),
    .COUT(_21976_),
    .SUM(_21977_));
 sky130_fd_sc_hd__fa_1 _43070_ (.A(_21977_),
    .B(_21931_),
    .CIN(_21969_),
    .COUT(_21978_),
    .SUM(_21979_));
 sky130_fd_sc_hd__fa_1 _43071_ (.A(_01963_),
    .B(_01964_),
    .CIN(_01965_),
    .COUT(_01966_),
    .SUM(_01967_));
 sky130_fd_sc_hd__fa_1 _43072_ (.A(_21941_),
    .B(_01968_),
    .CIN(_21933_),
    .COUT(_21980_),
    .SUM(_21981_));
 sky130_fd_sc_hd__fa_1 _43073_ (.A(_01969_),
    .B(_01970_),
    .CIN(_01971_),
    .COUT(_21982_),
    .SUM(_01972_));
 sky130_fd_sc_hd__fa_1 _43074_ (.A(_01973_),
    .B(_01974_),
    .CIN(_01923_),
    .COUT(_01975_),
    .SUM(_21983_));
 sky130_fd_sc_hd__fa_1 _43075_ (.A(_21983_),
    .B(_21943_),
    .CIN(_21981_),
    .COUT(_21984_),
    .SUM(_21985_));
 sky130_fd_sc_hd__fa_1 _43076_ (.A(_21947_),
    .B(_21985_),
    .CIN(_21937_),
    .COUT(_21986_),
    .SUM(_21987_));
 sky130_fd_sc_hd__fa_1 _43077_ (.A(_21987_),
    .B(_21939_),
    .CIN(_21979_),
    .COUT(_21988_),
    .SUM(_21989_));
 sky130_fd_sc_hd__fa_1 _43078_ (.A(_21945_),
    .B(_01771_),
    .CIN(_01770_),
    .COUT(_01976_),
    .SUM(_01977_));
 sky130_fd_sc_hd__fa_1 _43079_ (.A(_01978_),
    .B(_01977_),
    .CIN(_01979_),
    .COUT(_21990_),
    .SUM(_21991_));
 sky130_fd_sc_hd__fa_1 _43080_ (.A(_21953_),
    .B(_21991_),
    .CIN(_01726_),
    .COUT(_01980_),
    .SUM(_01981_));
 sky130_fd_sc_hd__fa_1 _43081_ (.A(_01982_),
    .B(_01983_),
    .CIN(_21949_),
    .COUT(_01984_),
    .SUM(_21992_));
 sky130_fd_sc_hd__fa_1 _43082_ (.A(_21992_),
    .B(_21951_),
    .CIN(_21989_),
    .COUT(_21993_),
    .SUM(_21994_));
 sky130_fd_sc_hd__fa_1 _43083_ (.A(_01985_),
    .B(_21956_),
    .CIN(_21994_),
    .COUT(_21995_),
    .SUM(_21996_));
 sky130_fd_sc_hd__fa_1 _43084_ (.A(_01986_),
    .B(_21958_),
    .CIN(_21996_),
    .COUT(_01987_),
    .SUM(_01988_));
 sky130_fd_sc_hd__fa_1 _43085_ (.A(_01990_),
    .B(_01991_),
    .CIN(_01992_),
    .COUT(_21997_),
    .SUM(_21998_));
 sky130_fd_sc_hd__fa_1 _43086_ (.A(_01993_),
    .B(_01994_),
    .CIN(_01995_),
    .COUT(_21999_),
    .SUM(_22000_));
 sky130_fd_sc_hd__fa_1 _43087_ (.A(_22000_),
    .B(_21960_),
    .CIN(_21998_),
    .COUT(_22001_),
    .SUM(_22002_));
 sky130_fd_sc_hd__fa_1 _43088_ (.A(_01996_),
    .B(_01997_),
    .CIN(_01998_),
    .COUT(_01999_),
    .SUM(_02000_));
 sky130_fd_sc_hd__fa_1 _43089_ (.A(_02001_),
    .B(_02002_),
    .CIN(_21962_),
    .COUT(_22003_),
    .SUM(_22004_));
 sky130_fd_sc_hd__fa_1 _43090_ (.A(_22004_),
    .B(_21964_),
    .CIN(_22002_),
    .COUT(_22005_),
    .SUM(_22006_));
 sky130_fd_sc_hd__fa_1 _43091_ (.A(_02003_),
    .B(_02004_),
    .CIN(_02005_),
    .COUT(_22007_),
    .SUM(_22008_));
 sky130_fd_sc_hd__fa_1 _43092_ (.A(_02006_),
    .B(_02007_),
    .CIN(_02008_),
    .COUT(_22009_),
    .SUM(_22010_));
 sky130_fd_sc_hd__fa_1 _43093_ (.A(_22010_),
    .B(_21970_),
    .CIN(_22008_),
    .COUT(_22011_),
    .SUM(_22012_));
 sky130_fd_sc_hd__fa_1 _43094_ (.A(_21974_),
    .B(_22012_),
    .CIN(_21966_),
    .COUT(_22013_),
    .SUM(_22014_));
 sky130_fd_sc_hd__fa_1 _43095_ (.A(_22014_),
    .B(_21968_),
    .CIN(_22006_),
    .COUT(_22015_),
    .SUM(_22016_));
 sky130_fd_sc_hd__fa_1 _43096_ (.A(_02009_),
    .B(_02010_),
    .CIN(_02011_),
    .COUT(_02012_),
    .SUM(_02013_));
 sky130_fd_sc_hd__fa_1 _43097_ (.A(_02014_),
    .B(_02015_),
    .CIN(_21972_),
    .COUT(_22017_),
    .SUM(_22018_));
 sky130_fd_sc_hd__fa_1 _43098_ (.A(_02016_),
    .B(_02017_),
    .CIN(_02018_),
    .COUT(_02019_),
    .SUM(_02020_));
 sky130_fd_sc_hd__fa_1 _43099_ (.A(_21982_),
    .B(_02021_),
    .CIN(_01922_),
    .COUT(_02022_),
    .SUM(_02023_));
 sky130_fd_sc_hd__fa_1 _43100_ (.A(_02024_),
    .B(_21980_),
    .CIN(_22018_),
    .COUT(_22019_),
    .SUM(_22020_));
 sky130_fd_sc_hd__fa_1 _43101_ (.A(_21984_),
    .B(_22020_),
    .CIN(_21976_),
    .COUT(_22021_),
    .SUM(_22022_));
 sky130_fd_sc_hd__fa_1 _43102_ (.A(_22022_),
    .B(_21978_),
    .CIN(_22016_),
    .COUT(_22023_),
    .SUM(_22024_));
 sky130_fd_sc_hd__fa_1 _43103_ (.A(_01976_),
    .B(_02025_),
    .CIN(_01977_),
    .COUT(_02026_),
    .SUM(_22025_));
 sky130_fd_sc_hd__fa_1 _43104_ (.A(_21990_),
    .B(_22025_),
    .CIN(_01726_),
    .COUT(_02027_),
    .SUM(_02028_));
 sky130_fd_sc_hd__fa_1 _43105_ (.A(_02029_),
    .B(_02030_),
    .CIN(_21986_),
    .COUT(_02031_),
    .SUM(_22026_));
 sky130_fd_sc_hd__fa_1 _43106_ (.A(_22026_),
    .B(_21988_),
    .CIN(_22024_),
    .COUT(_22027_),
    .SUM(_22028_));
 sky130_fd_sc_hd__fa_1 _43107_ (.A(_02032_),
    .B(_21993_),
    .CIN(_22028_),
    .COUT(_22029_),
    .SUM(_22030_));
 sky130_fd_sc_hd__fa_1 _43108_ (.A(_02033_),
    .B(_21995_),
    .CIN(_22030_),
    .COUT(_02034_),
    .SUM(_02035_));
 sky130_fd_sc_hd__fa_1 _43109_ (.A(_02037_),
    .B(_02038_),
    .CIN(_02039_),
    .COUT(_22031_),
    .SUM(_22032_));
 sky130_fd_sc_hd__fa_1 _43110_ (.A(_02040_),
    .B(_02041_),
    .CIN(_02042_),
    .COUT(_22033_),
    .SUM(_22034_));
 sky130_fd_sc_hd__fa_1 _43111_ (.A(_22034_),
    .B(_21997_),
    .CIN(_22032_),
    .COUT(_22035_),
    .SUM(_22036_));
 sky130_fd_sc_hd__fa_1 _43112_ (.A(_02043_),
    .B(_02044_),
    .CIN(_02045_),
    .COUT(_02046_),
    .SUM(_02047_));
 sky130_fd_sc_hd__fa_1 _43113_ (.A(_02048_),
    .B(_02049_),
    .CIN(_21999_),
    .COUT(_22037_),
    .SUM(_22038_));
 sky130_fd_sc_hd__fa_1 _43114_ (.A(_22038_),
    .B(_22001_),
    .CIN(_22036_),
    .COUT(_22039_),
    .SUM(_22040_));
 sky130_fd_sc_hd__fa_1 _43115_ (.A(_02050_),
    .B(_02051_),
    .CIN(_02052_),
    .COUT(_22041_),
    .SUM(_22042_));
 sky130_fd_sc_hd__fa_1 _43116_ (.A(_02054_),
    .B(_02055_),
    .CIN(_02056_),
    .COUT(_22043_),
    .SUM(_22044_));
 sky130_fd_sc_hd__fa_1 _43117_ (.A(_22044_),
    .B(_22007_),
    .CIN(_22042_),
    .COUT(_22045_),
    .SUM(_22046_));
 sky130_fd_sc_hd__fa_1 _43118_ (.A(_22011_),
    .B(_22046_),
    .CIN(_22003_),
    .COUT(_22047_),
    .SUM(_22048_));
 sky130_fd_sc_hd__fa_1 _43119_ (.A(_22048_),
    .B(_22005_),
    .CIN(_22040_),
    .COUT(_22049_),
    .SUM(_22050_));
 sky130_fd_sc_hd__fa_1 _43120_ (.A(_02057_),
    .B(_02058_),
    .CIN(_02059_),
    .COUT(_02060_),
    .SUM(_02061_));
 sky130_fd_sc_hd__fa_1 _43121_ (.A(_02062_),
    .B(_02063_),
    .CIN(_22009_),
    .COUT(_22051_),
    .SUM(_22052_));
 sky130_fd_sc_hd__fa_1 _43122_ (.A(_02064_),
    .B(_02016_),
    .CIN(_02018_),
    .COUT(_02065_),
    .SUM(_02066_));
 sky130_fd_sc_hd__fa_1 _43123_ (.A(_02067_),
    .B(_02068_),
    .CIN(_01922_),
    .COUT(_22053_),
    .SUM(_02069_));
 sky130_fd_sc_hd__fa_1 _43124_ (.A(_02070_),
    .B(_22017_),
    .CIN(_22052_),
    .COUT(_22054_),
    .SUM(_22055_));
 sky130_fd_sc_hd__fa_1 _43125_ (.A(_22019_),
    .B(_22055_),
    .CIN(_22013_),
    .COUT(_22056_),
    .SUM(_22057_));
 sky130_fd_sc_hd__fa_1 _43126_ (.A(_22057_),
    .B(_22015_),
    .CIN(_22050_),
    .COUT(_22058_),
    .SUM(_22059_));
 sky130_fd_sc_hd__fa_1 _43127_ (.A(_02071_),
    .B(_02072_),
    .CIN(_02073_),
    .COUT(_02074_),
    .SUM(_22060_));
 sky130_fd_sc_hd__fa_1 _43128_ (.A(_02075_),
    .B(_22060_),
    .CIN(_01727_),
    .COUT(_22061_),
    .SUM(_22062_));
 sky130_fd_sc_hd__fa_1 _43129_ (.A(_02076_),
    .B(_22062_),
    .CIN(_22021_),
    .COUT(_02077_),
    .SUM(_22063_));
 sky130_fd_sc_hd__fa_1 _43130_ (.A(_22063_),
    .B(_22023_),
    .CIN(_22059_),
    .COUT(_22064_),
    .SUM(_22065_));
 sky130_fd_sc_hd__fa_1 _43131_ (.A(_02078_),
    .B(_22027_),
    .CIN(_22065_),
    .COUT(_22066_),
    .SUM(_22067_));
 sky130_fd_sc_hd__fa_1 _43132_ (.A(_02079_),
    .B(_22029_),
    .CIN(_22067_),
    .COUT(_02080_),
    .SUM(_02081_));
 sky130_fd_sc_hd__fa_1 _43133_ (.A(_02083_),
    .B(_02084_),
    .CIN(_02085_),
    .COUT(_22068_),
    .SUM(_22069_));
 sky130_fd_sc_hd__fa_1 _43134_ (.A(_02086_),
    .B(_02087_),
    .CIN(_02088_),
    .COUT(_22070_),
    .SUM(_22071_));
 sky130_fd_sc_hd__fa_1 _43135_ (.A(_22071_),
    .B(_22031_),
    .CIN(_22069_),
    .COUT(_22072_),
    .SUM(_22073_));
 sky130_fd_sc_hd__fa_1 _43136_ (.A(_02089_),
    .B(_02090_),
    .CIN(_02091_),
    .COUT(_02092_),
    .SUM(_02093_));
 sky130_fd_sc_hd__fa_1 _43137_ (.A(_02094_),
    .B(_02095_),
    .CIN(_22033_),
    .COUT(_22074_),
    .SUM(_22075_));
 sky130_fd_sc_hd__fa_1 _43138_ (.A(_22075_),
    .B(_22035_),
    .CIN(_22073_),
    .COUT(_22076_),
    .SUM(_22077_));
 sky130_fd_sc_hd__fa_1 _43139_ (.A(_02096_),
    .B(_02097_),
    .CIN(_02098_),
    .COUT(_22078_),
    .SUM(_22079_));
 sky130_fd_sc_hd__fa_1 _43140_ (.A(_02099_),
    .B(_02100_),
    .CIN(_02101_),
    .COUT(_22080_),
    .SUM(_22081_));
 sky130_fd_sc_hd__fa_1 _43141_ (.A(_22081_),
    .B(_22041_),
    .CIN(_22079_),
    .COUT(_22082_),
    .SUM(_22083_));
 sky130_fd_sc_hd__fa_1 _43142_ (.A(_22045_),
    .B(_22083_),
    .CIN(_22037_),
    .COUT(_22084_),
    .SUM(_22085_));
 sky130_fd_sc_hd__fa_1 _43143_ (.A(_22085_),
    .B(_22039_),
    .CIN(_22077_),
    .COUT(_22086_),
    .SUM(_22087_));
 sky130_fd_sc_hd__fa_1 _43144_ (.A(_02102_),
    .B(_02103_),
    .CIN(_02104_),
    .COUT(_02105_),
    .SUM(_02106_));
 sky130_fd_sc_hd__fa_1 _43145_ (.A(_02107_),
    .B(_02108_),
    .CIN(_22043_),
    .COUT(_22088_),
    .SUM(_22089_));
 sky130_fd_sc_hd__fa_1 _43146_ (.A(_02109_),
    .B(_02068_),
    .CIN(_01922_),
    .COUT(_22090_),
    .SUM(_02110_));
 sky130_fd_sc_hd__fa_1 _43147_ (.A(_02111_),
    .B(_22051_),
    .CIN(_22089_),
    .COUT(_22091_),
    .SUM(_22092_));
 sky130_fd_sc_hd__fa_1 _43148_ (.A(_22054_),
    .B(_22092_),
    .CIN(_22047_),
    .COUT(_22093_),
    .SUM(_22094_));
 sky130_fd_sc_hd__fa_1 _43149_ (.A(_22094_),
    .B(_22049_),
    .CIN(_22087_),
    .COUT(_22095_),
    .SUM(_22096_));
 sky130_fd_sc_hd__fa_1 _43150_ (.A(_22053_),
    .B(_01976_),
    .CIN(_01977_),
    .COUT(_22097_),
    .SUM(_22098_));
 sky130_fd_sc_hd__fa_1 _43151_ (.A(_02112_),
    .B(_22098_),
    .CIN(_01726_),
    .COUT(_02113_),
    .SUM(_02114_));
 sky130_fd_sc_hd__fa_1 _43152_ (.A(_22061_),
    .B(_02115_),
    .CIN(_22056_),
    .COUT(_02116_),
    .SUM(_22099_));
 sky130_fd_sc_hd__fa_1 _43153_ (.A(_22099_),
    .B(_22058_),
    .CIN(_22096_),
    .COUT(_22100_),
    .SUM(_22101_));
 sky130_fd_sc_hd__fa_1 _43154_ (.A(_02117_),
    .B(_22064_),
    .CIN(_22101_),
    .COUT(_22102_),
    .SUM(_22103_));
 sky130_fd_sc_hd__fa_1 _43155_ (.A(_02118_),
    .B(_22066_),
    .CIN(_22103_),
    .COUT(_02119_),
    .SUM(_02120_));
 sky130_fd_sc_hd__fa_1 _43156_ (.A(_02122_),
    .B(_02123_),
    .CIN(_02124_),
    .COUT(_22104_),
    .SUM(_22105_));
 sky130_fd_sc_hd__fa_1 _43157_ (.A(_02125_),
    .B(_02126_),
    .CIN(_02127_),
    .COUT(_22106_),
    .SUM(_22107_));
 sky130_fd_sc_hd__fa_1 _43158_ (.A(_22107_),
    .B(_22068_),
    .CIN(_22105_),
    .COUT(_22108_),
    .SUM(_22109_));
 sky130_fd_sc_hd__fa_1 _43159_ (.A(_02128_),
    .B(_02129_),
    .CIN(_02130_),
    .COUT(_22110_),
    .SUM(_22111_));
 sky130_fd_sc_hd__fa_1 _43160_ (.A(_02131_),
    .B(_22111_),
    .CIN(_22070_),
    .COUT(_22112_),
    .SUM(_22113_));
 sky130_fd_sc_hd__fa_1 _43161_ (.A(_22113_),
    .B(_22072_),
    .CIN(_22109_),
    .COUT(_22114_),
    .SUM(_22115_));
 sky130_fd_sc_hd__fa_1 _43162_ (.A(_02132_),
    .B(_02133_),
    .CIN(_02134_),
    .COUT(_22116_),
    .SUM(_22117_));
 sky130_fd_sc_hd__fa_1 _43163_ (.A(_02135_),
    .B(_02136_),
    .CIN(_02137_),
    .COUT(_22118_),
    .SUM(_22119_));
 sky130_fd_sc_hd__fa_1 _43164_ (.A(_22119_),
    .B(_22078_),
    .CIN(_22117_),
    .COUT(_22120_),
    .SUM(_22121_));
 sky130_fd_sc_hd__fa_1 _43165_ (.A(_22082_),
    .B(_22121_),
    .CIN(_22074_),
    .COUT(_22122_),
    .SUM(_22123_));
 sky130_fd_sc_hd__fa_1 _43166_ (.A(_22123_),
    .B(_22076_),
    .CIN(_22115_),
    .COUT(_22124_),
    .SUM(_22125_));
 sky130_fd_sc_hd__fa_1 _43167_ (.A(_02138_),
    .B(_02139_),
    .CIN(_02140_),
    .COUT(_22126_),
    .SUM(_22127_));
 sky130_fd_sc_hd__fa_1 _43168_ (.A(_02141_),
    .B(_22127_),
    .CIN(_22080_),
    .COUT(_22128_),
    .SUM(_22129_));
 sky130_fd_sc_hd__fa_1 _43169_ (.A(_22088_),
    .B(_22129_),
    .CIN(_02111_),
    .COUT(_22130_),
    .SUM(_22131_));
 sky130_fd_sc_hd__fa_1 _43170_ (.A(_22091_),
    .B(_22131_),
    .CIN(_22084_),
    .COUT(_22132_),
    .SUM(_22133_));
 sky130_fd_sc_hd__fa_1 _43171_ (.A(_22133_),
    .B(_22086_),
    .CIN(_22125_),
    .COUT(_22134_),
    .SUM(_22135_));
 sky130_fd_sc_hd__fa_1 _43172_ (.A(_22090_),
    .B(_01976_),
    .CIN(_01977_),
    .COUT(_22136_),
    .SUM(_22137_));
 sky130_fd_sc_hd__fa_1 _43173_ (.A(_22097_),
    .B(_22137_),
    .CIN(_01726_),
    .COUT(_02142_),
    .SUM(_02143_));
 sky130_fd_sc_hd__fa_1 _43174_ (.A(_02144_),
    .B(_02145_),
    .CIN(_22093_),
    .COUT(_02146_),
    .SUM(_22138_));
 sky130_fd_sc_hd__fa_1 _43175_ (.A(_22138_),
    .B(_22095_),
    .CIN(_22135_),
    .COUT(_22139_),
    .SUM(_22140_));
 sky130_fd_sc_hd__fa_1 _43176_ (.A(_02147_),
    .B(_22100_),
    .CIN(_22140_),
    .COUT(_22141_),
    .SUM(_22142_));
 sky130_fd_sc_hd__fa_1 _43177_ (.A(_02148_),
    .B(_22102_),
    .CIN(_22142_),
    .COUT(_02149_),
    .SUM(_02150_));
 sky130_fd_sc_hd__fa_1 _43178_ (.A(_02152_),
    .B(_02153_),
    .CIN(_02154_),
    .COUT(_22143_),
    .SUM(_22144_));
 sky130_fd_sc_hd__fa_1 _43179_ (.A(_02155_),
    .B(_02156_),
    .CIN(_02157_),
    .COUT(_22145_),
    .SUM(_22146_));
 sky130_fd_sc_hd__fa_1 _43180_ (.A(_22146_),
    .B(_22104_),
    .CIN(_22144_),
    .COUT(_22147_),
    .SUM(_22148_));
 sky130_fd_sc_hd__fa_1 _43181_ (.A(_02158_),
    .B(_02159_),
    .CIN(_02160_),
    .COUT(_02161_),
    .SUM(_02162_));
 sky130_fd_sc_hd__fa_1 _43182_ (.A(_22110_),
    .B(_02163_),
    .CIN(_22106_),
    .COUT(_22149_),
    .SUM(_22150_));
 sky130_fd_sc_hd__fa_1 _43183_ (.A(_22150_),
    .B(_22108_),
    .CIN(_22148_),
    .COUT(_22151_),
    .SUM(_22152_));
 sky130_fd_sc_hd__fa_1 _43184_ (.A(_02164_),
    .B(_02165_),
    .CIN(_02166_),
    .COUT(_22153_),
    .SUM(_22154_));
 sky130_fd_sc_hd__fa_1 _43185_ (.A(_02167_),
    .B(_02168_),
    .CIN(_02169_),
    .COUT(_22155_),
    .SUM(_22156_));
 sky130_fd_sc_hd__fa_1 _43186_ (.A(_22156_),
    .B(_22116_),
    .CIN(_22154_),
    .COUT(_22157_),
    .SUM(_22158_));
 sky130_fd_sc_hd__fa_1 _43187_ (.A(_22120_),
    .B(_22158_),
    .CIN(_22112_),
    .COUT(_22159_),
    .SUM(_22160_));
 sky130_fd_sc_hd__fa_1 _43188_ (.A(_22160_),
    .B(_22114_),
    .CIN(_22152_),
    .COUT(_22161_),
    .SUM(_22162_));
 sky130_fd_sc_hd__fa_1 _43189_ (.A(_02170_),
    .B(_02171_),
    .CIN(_02102_),
    .COUT(_02172_),
    .SUM(_02173_));
 sky130_fd_sc_hd__fa_1 _43190_ (.A(_22126_),
    .B(_02174_),
    .CIN(_22118_),
    .COUT(_22163_),
    .SUM(_22164_));
 sky130_fd_sc_hd__fa_1 _43191_ (.A(_22128_),
    .B(_22164_),
    .CIN(_02111_),
    .COUT(_22165_),
    .SUM(_22166_));
 sky130_fd_sc_hd__fa_1 _43192_ (.A(_22130_),
    .B(_22166_),
    .CIN(_22122_),
    .COUT(_22167_),
    .SUM(_22168_));
 sky130_fd_sc_hd__fa_1 _43193_ (.A(_22168_),
    .B(_22124_),
    .CIN(_22162_),
    .COUT(_22169_),
    .SUM(_22170_));
 sky130_fd_sc_hd__fa_1 _43194_ (.A(_22136_),
    .B(_22137_),
    .CIN(_01726_),
    .COUT(_02175_),
    .SUM(_02176_));
 sky130_fd_sc_hd__fa_1 _43195_ (.A(_02177_),
    .B(net789),
    .CIN(_22132_),
    .COUT(_02179_),
    .SUM(_22171_));
 sky130_fd_sc_hd__fa_1 _43196_ (.A(_22171_),
    .B(_22134_),
    .CIN(_22170_),
    .COUT(_22172_),
    .SUM(_22173_));
 sky130_fd_sc_hd__fa_1 _43197_ (.A(_02180_),
    .B(_22139_),
    .CIN(_22173_),
    .COUT(_22174_),
    .SUM(_22175_));
 sky130_fd_sc_hd__fa_1 _43198_ (.A(_02181_),
    .B(_22141_),
    .CIN(_22175_),
    .COUT(_02182_),
    .SUM(_02183_));
 sky130_fd_sc_hd__fa_1 _43199_ (.A(_02185_),
    .B(_02186_),
    .CIN(_02187_),
    .COUT(_22176_),
    .SUM(_22177_));
 sky130_fd_sc_hd__fa_1 _43200_ (.A(_02188_),
    .B(_02189_),
    .CIN(_02190_),
    .COUT(_02191_),
    .SUM(_02192_));
 sky130_fd_sc_hd__fa_1 _43201_ (.A(_02193_),
    .B(_22143_),
    .CIN(_22177_),
    .COUT(_22178_),
    .SUM(_22179_));
 sky130_fd_sc_hd__fa_1 _43202_ (.A(_02194_),
    .B(_02195_),
    .CIN(_02196_),
    .COUT(_22180_),
    .SUM(_22181_));
 sky130_fd_sc_hd__fa_1 _43203_ (.A(_02197_),
    .B(_22181_),
    .CIN(_22145_),
    .COUT(_22182_),
    .SUM(_22183_));
 sky130_fd_sc_hd__fa_1 _43204_ (.A(_22183_),
    .B(_22147_),
    .CIN(_22179_),
    .COUT(_22184_),
    .SUM(_22185_));
 sky130_fd_sc_hd__fa_1 _43205_ (.A(_02198_),
    .B(_02199_),
    .CIN(_02200_),
    .COUT(_22186_),
    .SUM(_22187_));
 sky130_fd_sc_hd__fa_1 _43206_ (.A(_02201_),
    .B(_02202_),
    .CIN(_02203_),
    .COUT(_22188_),
    .SUM(_22189_));
 sky130_fd_sc_hd__fa_1 _43207_ (.A(_22189_),
    .B(_22153_),
    .CIN(_22187_),
    .COUT(_22190_),
    .SUM(_22191_));
 sky130_fd_sc_hd__fa_1 _43208_ (.A(_22157_),
    .B(_22191_),
    .CIN(_22149_),
    .COUT(_22192_),
    .SUM(_22193_));
 sky130_fd_sc_hd__fa_1 _43209_ (.A(_22193_),
    .B(_22151_),
    .CIN(_22185_),
    .COUT(_22194_),
    .SUM(_22195_));
 sky130_fd_sc_hd__fa_1 _43210_ (.A(_02204_),
    .B(_22155_),
    .CIN(_02174_),
    .COUT(_22196_),
    .SUM(_22197_));
 sky130_fd_sc_hd__fa_1 _43211_ (.A(_22163_),
    .B(_22197_),
    .CIN(_02111_),
    .COUT(_22198_),
    .SUM(_22199_));
 sky130_fd_sc_hd__fa_1 _43212_ (.A(_22165_),
    .B(_22199_),
    .CIN(_22159_),
    .COUT(_22200_),
    .SUM(_22201_));
 sky130_fd_sc_hd__fa_1 _43213_ (.A(_22201_),
    .B(_22161_),
    .CIN(_22195_),
    .COUT(_22202_),
    .SUM(_22203_));
 sky130_fd_sc_hd__fa_1 _43214_ (.A(net788),
    .B(_22167_),
    .CIN(_02178_),
    .COUT(_02206_),
    .SUM(_22204_));
 sky130_fd_sc_hd__fa_1 _43215_ (.A(_22204_),
    .B(_22169_),
    .CIN(_22203_),
    .COUT(_22205_),
    .SUM(_22206_));
 sky130_fd_sc_hd__fa_1 _43216_ (.A(_02207_),
    .B(_22172_),
    .CIN(_22206_),
    .COUT(_22207_),
    .SUM(_22208_));
 sky130_fd_sc_hd__fa_1 _43217_ (.A(_02208_),
    .B(_22174_),
    .CIN(_22208_),
    .COUT(_02209_),
    .SUM(_02210_));
 sky130_fd_sc_hd__fa_1 _43218_ (.A(_02212_),
    .B(_02213_),
    .CIN(_02214_),
    .COUT(_22209_),
    .SUM(_22210_));
 sky130_fd_sc_hd__fa_1 _43219_ (.A(_02215_),
    .B(_02216_),
    .CIN(_02217_),
    .COUT(_02218_),
    .SUM(_02219_));
 sky130_fd_sc_hd__fa_1 _43220_ (.A(_02220_),
    .B(_22176_),
    .CIN(_22210_),
    .COUT(_22211_),
    .SUM(_22212_));
 sky130_fd_sc_hd__fa_1 _43221_ (.A(_02221_),
    .B(_02222_),
    .CIN(_02223_),
    .COUT(_02224_),
    .SUM(_02225_));
 sky130_fd_sc_hd__fa_1 _43222_ (.A(_22180_),
    .B(_02226_),
    .CIN(_02227_),
    .COUT(_22213_),
    .SUM(_22214_));
 sky130_fd_sc_hd__fa_1 _43223_ (.A(_22214_),
    .B(_22178_),
    .CIN(_22212_),
    .COUT(_22215_),
    .SUM(_22216_));
 sky130_fd_sc_hd__fa_1 _43224_ (.A(_02228_),
    .B(_02229_),
    .CIN(_02230_),
    .COUT(_02231_),
    .SUM(_02232_));
 sky130_fd_sc_hd__fa_1 _43225_ (.A(_02233_),
    .B(_02234_),
    .CIN(_02201_),
    .COUT(_02235_),
    .SUM(_22217_));
 sky130_fd_sc_hd__fa_1 _43226_ (.A(_22217_),
    .B(_22186_),
    .CIN(_02238_),
    .COUT(_22218_),
    .SUM(_22219_));
 sky130_fd_sc_hd__fa_1 _43227_ (.A(_22190_),
    .B(_22219_),
    .CIN(_22182_),
    .COUT(_22220_),
    .SUM(_22221_));
 sky130_fd_sc_hd__fa_1 _43228_ (.A(_22221_),
    .B(_22184_),
    .CIN(_22216_),
    .COUT(_22222_),
    .SUM(_22223_));
 sky130_fd_sc_hd__fa_1 _43229_ (.A(_22188_),
    .B(_02204_),
    .CIN(_02174_),
    .COUT(_02239_),
    .SUM(_22224_));
 sky130_fd_sc_hd__fa_1 _43230_ (.A(_22196_),
    .B(_22224_),
    .CIN(_02111_),
    .COUT(_22225_),
    .SUM(_22226_));
 sky130_fd_sc_hd__fa_1 _43231_ (.A(_22198_),
    .B(_22226_),
    .CIN(_22192_),
    .COUT(_22227_),
    .SUM(_22228_));
 sky130_fd_sc_hd__fa_1 _43232_ (.A(_22228_),
    .B(_22194_),
    .CIN(_22223_),
    .COUT(_22229_),
    .SUM(_22230_));
 sky130_fd_sc_hd__fa_1 _43233_ (.A(_22200_),
    .B(net788),
    .CIN(_02178_),
    .COUT(_02240_),
    .SUM(_22231_));
 sky130_fd_sc_hd__fa_1 _43234_ (.A(_22231_),
    .B(_22202_),
    .CIN(_22230_),
    .COUT(_22232_),
    .SUM(_22233_));
 sky130_fd_sc_hd__fa_1 _43235_ (.A(_02241_),
    .B(_22205_),
    .CIN(_22233_),
    .COUT(_22234_),
    .SUM(_22235_));
 sky130_fd_sc_hd__fa_1 _43236_ (.A(_02242_),
    .B(_22207_),
    .CIN(_22235_),
    .COUT(_02243_),
    .SUM(_02244_));
 sky130_fd_sc_hd__fa_1 _43237_ (.A(_02246_),
    .B(_02247_),
    .CIN(_02248_),
    .COUT(_22236_),
    .SUM(_22237_));
 sky130_fd_sc_hd__fa_1 _43238_ (.A(_02249_),
    .B(_02250_),
    .CIN(_02251_),
    .COUT(_02252_),
    .SUM(_02253_));
 sky130_fd_sc_hd__fa_1 _43239_ (.A(_02254_),
    .B(_22209_),
    .CIN(_22237_),
    .COUT(_22238_),
    .SUM(_22239_));
 sky130_fd_sc_hd__fa_1 _43240_ (.A(_02255_),
    .B(_02256_),
    .CIN(_02257_),
    .COUT(_02258_),
    .SUM(_02259_));
 sky130_fd_sc_hd__fa_1 _43241_ (.A(_02260_),
    .B(_02261_),
    .CIN(_02262_),
    .COUT(_22240_),
    .SUM(_22241_));
 sky130_fd_sc_hd__fa_1 _43242_ (.A(_22241_),
    .B(_22211_),
    .CIN(_22239_),
    .COUT(_22242_),
    .SUM(_22243_));
 sky130_fd_sc_hd__fa_1 _43243_ (.A(_02263_),
    .B(_02264_),
    .CIN(_02265_),
    .COUT(_02266_),
    .SUM(_02267_));
 sky130_fd_sc_hd__fa_1 _43244_ (.A(_02268_),
    .B(_02236_),
    .CIN(_02237_),
    .COUT(_22244_),
    .SUM(_02269_));
 sky130_fd_sc_hd__fa_1 _43245_ (.A(_02270_),
    .B(_02271_),
    .CIN(_02272_),
    .COUT(_22245_),
    .SUM(_22246_));
 sky130_fd_sc_hd__fa_1 _43246_ (.A(_22218_),
    .B(_22246_),
    .CIN(_22213_),
    .COUT(_22247_),
    .SUM(_22248_));
 sky130_fd_sc_hd__fa_1 _43247_ (.A(_22248_),
    .B(_22215_),
    .CIN(_22243_),
    .COUT(_22249_),
    .SUM(_22250_));
 sky130_fd_sc_hd__fa_1 _43248_ (.A(_02273_),
    .B(_02172_),
    .CIN(_02173_),
    .COUT(_02274_),
    .SUM(_22251_));
 sky130_fd_sc_hd__fa_1 _43249_ (.A(_02275_),
    .B(_22251_),
    .CIN(_02110_),
    .COUT(_02276_),
    .SUM(_02277_));
 sky130_fd_sc_hd__fa_1 _43250_ (.A(_22225_),
    .B(_02278_),
    .CIN(_22220_),
    .COUT(_22252_),
    .SUM(_22253_));
 sky130_fd_sc_hd__fa_1 _43251_ (.A(_22253_),
    .B(_22222_),
    .CIN(_22250_),
    .COUT(_22254_),
    .SUM(_22255_));
 sky130_fd_sc_hd__fa_1 _43252_ (.A(_22227_),
    .B(_02205_),
    .CIN(_02178_),
    .COUT(_02279_),
    .SUM(_22256_));
 sky130_fd_sc_hd__fa_1 _43253_ (.A(_22256_),
    .B(_22229_),
    .CIN(_22255_),
    .COUT(_22257_),
    .SUM(_22258_));
 sky130_fd_sc_hd__fa_1 _43254_ (.A(_02280_),
    .B(_22232_),
    .CIN(_22258_),
    .COUT(_22259_),
    .SUM(_22260_));
 sky130_fd_sc_hd__fa_1 _43255_ (.A(_02281_),
    .B(_22234_),
    .CIN(_22260_),
    .COUT(_02282_),
    .SUM(_02283_));
 sky130_fd_sc_hd__fa_1 _43256_ (.A(_02285_),
    .B(_02286_),
    .CIN(_02287_),
    .COUT(_22261_),
    .SUM(_22262_));
 sky130_fd_sc_hd__fa_1 _43257_ (.A(_02288_),
    .B(_02289_),
    .CIN(_02290_),
    .COUT(_02291_),
    .SUM(_02292_));
 sky130_fd_sc_hd__fa_1 _43258_ (.A(_02293_),
    .B(_22236_),
    .CIN(_22262_),
    .COUT(_22263_),
    .SUM(_22264_));
 sky130_fd_sc_hd__fa_1 _43259_ (.A(_02294_),
    .B(_02295_),
    .CIN(_02296_),
    .COUT(_02297_),
    .SUM(_02298_));
 sky130_fd_sc_hd__fa_1 _43260_ (.A(_02299_),
    .B(_02300_),
    .CIN(_02301_),
    .COUT(_22265_),
    .SUM(_22266_));
 sky130_fd_sc_hd__fa_1 _43261_ (.A(_22266_),
    .B(_22238_),
    .CIN(_22264_),
    .COUT(_22267_),
    .SUM(_22268_));
 sky130_fd_sc_hd__fa_1 _43262_ (.A(_02302_),
    .B(_02303_),
    .CIN(_02304_),
    .COUT(_02305_),
    .SUM(_02306_));
 sky130_fd_sc_hd__fa_1 _43263_ (.A(_02307_),
    .B(_02308_),
    .CIN(_02270_),
    .COUT(_22269_),
    .SUM(_22270_));
 sky130_fd_sc_hd__fa_1 _43264_ (.A(_22245_),
    .B(_22270_),
    .CIN(_22240_),
    .COUT(_22271_),
    .SUM(_22272_));
 sky130_fd_sc_hd__fa_1 _43265_ (.A(_22272_),
    .B(_22242_),
    .CIN(_22268_),
    .COUT(_22273_),
    .SUM(_22274_));
 sky130_fd_sc_hd__fa_1 _43266_ (.A(_22244_),
    .B(_02172_),
    .CIN(_02173_),
    .COUT(_22275_),
    .SUM(_02309_));
 sky130_fd_sc_hd__fa_1 _43267_ (.A(_02310_),
    .B(_02311_),
    .CIN(_02111_),
    .COUT(_22276_),
    .SUM(_22277_));
 sky130_fd_sc_hd__fa_1 _43268_ (.A(_02312_),
    .B(_22277_),
    .CIN(_22247_),
    .COUT(_22278_),
    .SUM(_22279_));
 sky130_fd_sc_hd__fa_1 _43269_ (.A(_22279_),
    .B(_22249_),
    .CIN(_22274_),
    .COUT(_22280_),
    .SUM(_22281_));
 sky130_fd_sc_hd__fa_1 _43270_ (.A(_22252_),
    .B(_02205_),
    .CIN(_02178_),
    .COUT(_02313_),
    .SUM(_22282_));
 sky130_fd_sc_hd__fa_1 _43271_ (.A(_22282_),
    .B(_22254_),
    .CIN(_22281_),
    .COUT(_22283_),
    .SUM(_22284_));
 sky130_fd_sc_hd__fa_1 _43272_ (.A(_02314_),
    .B(_22257_),
    .CIN(_22284_),
    .COUT(_22285_),
    .SUM(_22286_));
 sky130_fd_sc_hd__fa_1 _43273_ (.A(_02315_),
    .B(_22259_),
    .CIN(_22286_),
    .COUT(_02316_),
    .SUM(_02317_));
 sky130_fd_sc_hd__fa_1 _43274_ (.A(_02319_),
    .B(_02320_),
    .CIN(_02321_),
    .COUT(_22287_),
    .SUM(_22288_));
 sky130_fd_sc_hd__fa_1 _43275_ (.A(_02322_),
    .B(_02323_),
    .CIN(_02324_),
    .COUT(_22289_),
    .SUM(_22290_));
 sky130_fd_sc_hd__fa_1 _43276_ (.A(_22290_),
    .B(_22261_),
    .CIN(_22288_),
    .COUT(_22291_),
    .SUM(_22292_));
 sky130_fd_sc_hd__fa_1 _43277_ (.A(_02325_),
    .B(_02326_),
    .CIN(_02327_),
    .COUT(_02328_),
    .SUM(_02329_));
 sky130_fd_sc_hd__fa_1 _43278_ (.A(_02330_),
    .B(_02331_),
    .CIN(_02332_),
    .COUT(_22293_),
    .SUM(_22294_));
 sky130_fd_sc_hd__fa_1 _43279_ (.A(_22294_),
    .B(_22263_),
    .CIN(_22292_),
    .COUT(_22295_),
    .SUM(_22296_));
 sky130_fd_sc_hd__fa_1 _43280_ (.A(_02333_),
    .B(_02334_),
    .CIN(_02335_),
    .COUT(_22297_),
    .SUM(_22298_));
 sky130_fd_sc_hd__fa_1 _43281_ (.A(_02336_),
    .B(_22298_),
    .CIN(_02270_),
    .COUT(_22299_),
    .SUM(_22300_));
 sky130_fd_sc_hd__fa_1 _43282_ (.A(_22269_),
    .B(_22300_),
    .CIN(_22265_),
    .COUT(_22301_),
    .SUM(_22302_));
 sky130_fd_sc_hd__fa_1 _43283_ (.A(_22302_),
    .B(_22267_),
    .CIN(_22296_),
    .COUT(_22303_),
    .SUM(_22304_));
 sky130_fd_sc_hd__fa_1 _43284_ (.A(_22275_),
    .B(_02309_),
    .CIN(_02110_),
    .COUT(_02337_),
    .SUM(_02338_));
 sky130_fd_sc_hd__fa_1 _43285_ (.A(_22276_),
    .B(_02339_),
    .CIN(_22271_),
    .COUT(_22305_),
    .SUM(_22306_));
 sky130_fd_sc_hd__fa_1 _43286_ (.A(_22306_),
    .B(_22273_),
    .CIN(_22304_),
    .COUT(_22307_),
    .SUM(_22308_));
 sky130_fd_sc_hd__fa_1 _43287_ (.A(_22278_),
    .B(_02205_),
    .CIN(net789),
    .COUT(_02340_),
    .SUM(_22309_));
 sky130_fd_sc_hd__fa_1 _43288_ (.A(_22309_),
    .B(_22280_),
    .CIN(_22308_),
    .COUT(_22310_),
    .SUM(_22311_));
 sky130_fd_sc_hd__fa_1 _43289_ (.A(_02341_),
    .B(_22283_),
    .CIN(_22311_),
    .COUT(_22312_),
    .SUM(_22313_));
 sky130_fd_sc_hd__fa_1 _43290_ (.A(_02342_),
    .B(_22285_),
    .CIN(_22313_),
    .COUT(_02343_),
    .SUM(_02344_));
 sky130_fd_sc_hd__fa_1 _43291_ (.A(_02346_),
    .B(_02347_),
    .CIN(_02348_),
    .COUT(_02349_),
    .SUM(_02350_));
 sky130_fd_sc_hd__fa_1 _43292_ (.A(_02351_),
    .B(_02352_),
    .CIN(_02353_),
    .COUT(_02354_),
    .SUM(_02355_));
 sky130_fd_sc_hd__fa_1 _43293_ (.A(_02356_),
    .B(_22287_),
    .CIN(_02357_),
    .COUT(_22314_),
    .SUM(_22315_));
 sky130_fd_sc_hd__fa_1 _43294_ (.A(_02358_),
    .B(_02359_),
    .CIN(_02360_),
    .COUT(_02361_),
    .SUM(_02362_));
 sky130_fd_sc_hd__fa_1 _43295_ (.A(_02363_),
    .B(_02364_),
    .CIN(_22289_),
    .COUT(_22316_),
    .SUM(_22317_));
 sky130_fd_sc_hd__fa_1 _43296_ (.A(_22317_),
    .B(_22291_),
    .CIN(_22315_),
    .COUT(_22318_),
    .SUM(_22319_));
 sky130_fd_sc_hd__fa_1 _43297_ (.A(_02365_),
    .B(_02366_),
    .CIN(_02302_),
    .COUT(_22320_),
    .SUM(_02367_));
 sky130_fd_sc_hd__fa_1 _43298_ (.A(_22297_),
    .B(_02368_),
    .CIN(_02270_),
    .COUT(_22321_),
    .SUM(_22322_));
 sky130_fd_sc_hd__fa_1 _43299_ (.A(_22299_),
    .B(_22322_),
    .CIN(_22293_),
    .COUT(_22323_),
    .SUM(_22324_));
 sky130_fd_sc_hd__fa_1 _43300_ (.A(_22324_),
    .B(_22295_),
    .CIN(_22319_),
    .COUT(_22325_),
    .SUM(_22326_));
 sky130_fd_sc_hd__fa_1 _43301_ (.A(_02369_),
    .B(_22301_),
    .CIN(_02339_),
    .COUT(_22327_),
    .SUM(_22328_));
 sky130_fd_sc_hd__fa_1 _43302_ (.A(_22328_),
    .B(_22303_),
    .CIN(_22326_),
    .COUT(_22329_),
    .SUM(_22330_));
 sky130_fd_sc_hd__fa_1 _43303_ (.A(_22305_),
    .B(net788),
    .CIN(net789),
    .COUT(_02370_),
    .SUM(_22331_));
 sky130_fd_sc_hd__fa_1 _43304_ (.A(_22331_),
    .B(_22307_),
    .CIN(_22330_),
    .COUT(_22332_),
    .SUM(_22333_));
 sky130_fd_sc_hd__fa_1 _43305_ (.A(_02371_),
    .B(_22310_),
    .CIN(_22333_),
    .COUT(_22334_),
    .SUM(_22335_));
 sky130_fd_sc_hd__fa_1 _43306_ (.A(_02372_),
    .B(_22312_),
    .CIN(_22335_),
    .COUT(_02373_),
    .SUM(_02374_));
 sky130_fd_sc_hd__fa_1 _43307_ (.A(_02376_),
    .B(_02377_),
    .CIN(_02378_),
    .COUT(_02379_),
    .SUM(_02380_));
 sky130_fd_sc_hd__fa_1 _43308_ (.A(_02381_),
    .B(_02382_),
    .CIN(_02383_),
    .COUT(_02384_),
    .SUM(_02385_));
 sky130_fd_sc_hd__fa_1 _43309_ (.A(_02386_),
    .B(_02387_),
    .CIN(_02388_),
    .COUT(_22336_),
    .SUM(_22337_));
 sky130_fd_sc_hd__fa_1 _43310_ (.A(_02389_),
    .B(_02390_),
    .CIN(_02391_),
    .COUT(_02392_),
    .SUM(_02393_));
 sky130_fd_sc_hd__fa_1 _43311_ (.A(_02394_),
    .B(_02395_),
    .CIN(_02396_),
    .COUT(_22338_),
    .SUM(_22339_));
 sky130_fd_sc_hd__fa_1 _43312_ (.A(_22339_),
    .B(_22314_),
    .CIN(_22337_),
    .COUT(_22340_),
    .SUM(_22341_));
 sky130_fd_sc_hd__fa_1 _43313_ (.A(_22320_),
    .B(_02367_),
    .CIN(_02269_),
    .COUT(_02397_),
    .SUM(_02398_));
 sky130_fd_sc_hd__fa_1 _43314_ (.A(_22321_),
    .B(_02399_),
    .CIN(_22316_),
    .COUT(_22342_),
    .SUM(_22343_));
 sky130_fd_sc_hd__fa_1 _43315_ (.A(_22343_),
    .B(_22318_),
    .CIN(_22341_),
    .COUT(_22344_),
    .SUM(_22345_));
 sky130_fd_sc_hd__fa_1 _43316_ (.A(_22323_),
    .B(_02369_),
    .CIN(_02339_),
    .COUT(_22346_),
    .SUM(_22347_));
 sky130_fd_sc_hd__fa_1 _43317_ (.A(_22347_),
    .B(_22325_),
    .CIN(_22345_),
    .COUT(_22348_),
    .SUM(_22349_));
 sky130_fd_sc_hd__fa_1 _43318_ (.A(_22327_),
    .B(net788),
    .CIN(net789),
    .COUT(_02400_),
    .SUM(_22350_));
 sky130_fd_sc_hd__fa_1 _43319_ (.A(_22350_),
    .B(_22329_),
    .CIN(_22349_),
    .COUT(_22351_),
    .SUM(_22352_));
 sky130_fd_sc_hd__fa_1 _43320_ (.A(_02401_),
    .B(_22332_),
    .CIN(_22352_),
    .COUT(_22353_),
    .SUM(_22354_));
 sky130_fd_sc_hd__fa_1 _43321_ (.A(_02402_),
    .B(_22334_),
    .CIN(_22354_),
    .COUT(_02403_),
    .SUM(_02404_));
 sky130_fd_sc_hd__fa_1 _43322_ (.A(_02406_),
    .B(_02407_),
    .CIN(_02408_),
    .COUT(_02409_),
    .SUM(_02410_));
 sky130_fd_sc_hd__fa_1 _43323_ (.A(_02411_),
    .B(_02412_),
    .CIN(_02413_),
    .COUT(_02414_),
    .SUM(_02415_));
 sky130_fd_sc_hd__fa_1 _43324_ (.A(_02416_),
    .B(_02417_),
    .CIN(_02418_),
    .COUT(_22355_),
    .SUM(_22356_));
 sky130_fd_sc_hd__fa_1 _43325_ (.A(_02419_),
    .B(_02420_),
    .CIN(_02421_),
    .COUT(_22357_),
    .SUM(_22358_));
 sky130_fd_sc_hd__fa_1 _43326_ (.A(_02422_),
    .B(_22358_),
    .CIN(_02423_),
    .COUT(_22359_),
    .SUM(_22360_));
 sky130_fd_sc_hd__fa_1 _43327_ (.A(_22360_),
    .B(_22336_),
    .CIN(_22356_),
    .COUT(_22361_),
    .SUM(_22362_));
 sky130_fd_sc_hd__fa_1 _43328_ (.A(_02424_),
    .B(_22338_),
    .CIN(_02399_),
    .COUT(_22363_),
    .SUM(_22364_));
 sky130_fd_sc_hd__fa_1 _43329_ (.A(_22364_),
    .B(_22340_),
    .CIN(_22362_),
    .COUT(_22365_),
    .SUM(_22366_));
 sky130_fd_sc_hd__fa_1 _43330_ (.A(_22342_),
    .B(_02369_),
    .CIN(_02339_),
    .COUT(_22367_),
    .SUM(_22368_));
 sky130_fd_sc_hd__fa_1 _43331_ (.A(_22368_),
    .B(_22344_),
    .CIN(_22366_),
    .COUT(_22369_),
    .SUM(_22370_));
 sky130_fd_sc_hd__fa_1 _43332_ (.A(_22346_),
    .B(net788),
    .CIN(net789),
    .COUT(_02425_),
    .SUM(_22371_));
 sky130_fd_sc_hd__fa_1 _43333_ (.A(_22371_),
    .B(_22348_),
    .CIN(_22370_),
    .COUT(_22372_),
    .SUM(_22373_));
 sky130_fd_sc_hd__fa_1 _43334_ (.A(_02426_),
    .B(_22351_),
    .CIN(_22373_),
    .COUT(_22374_),
    .SUM(_22375_));
 sky130_fd_sc_hd__fa_1 _43335_ (.A(_02427_),
    .B(_22353_),
    .CIN(_22375_),
    .COUT(_02428_),
    .SUM(_02429_));
 sky130_fd_sc_hd__fa_1 _43336_ (.A(_02431_),
    .B(_02432_),
    .CIN(_02433_),
    .COUT(_02434_),
    .SUM(_02435_));
 sky130_fd_sc_hd__fa_1 _43337_ (.A(_02436_),
    .B(_02437_),
    .CIN(_02438_),
    .COUT(_02439_),
    .SUM(_02440_));
 sky130_fd_sc_hd__fa_1 _43338_ (.A(_02441_),
    .B(_02442_),
    .CIN(_02443_),
    .COUT(_22376_),
    .SUM(_22377_));
 sky130_fd_sc_hd__fa_1 _43339_ (.A(_02444_),
    .B(_02445_),
    .CIN(_02389_),
    .COUT(_02446_),
    .SUM(_02447_));
 sky130_fd_sc_hd__fa_1 _43340_ (.A(_22357_),
    .B(_02448_),
    .CIN(_02449_),
    .COUT(_22378_),
    .SUM(_22379_));
 sky130_fd_sc_hd__fa_1 _43341_ (.A(_22379_),
    .B(_22355_),
    .CIN(_22377_),
    .COUT(_22380_),
    .SUM(_22381_));
 sky130_fd_sc_hd__fa_1 _43342_ (.A(_22359_),
    .B(_02424_),
    .CIN(_02399_),
    .COUT(_22382_),
    .SUM(_22383_));
 sky130_fd_sc_hd__fa_1 _43343_ (.A(_22383_),
    .B(_22361_),
    .CIN(_22381_),
    .COUT(_22384_),
    .SUM(_22385_));
 sky130_fd_sc_hd__fa_1 _43344_ (.A(_22363_),
    .B(_02369_),
    .CIN(_02339_),
    .COUT(_22386_),
    .SUM(_22387_));
 sky130_fd_sc_hd__fa_1 _43345_ (.A(_22387_),
    .B(_22365_),
    .CIN(_22385_),
    .COUT(_22388_),
    .SUM(_22389_));
 sky130_fd_sc_hd__fa_1 _43346_ (.A(_22367_),
    .B(net788),
    .CIN(net789),
    .COUT(_02450_),
    .SUM(_22390_));
 sky130_fd_sc_hd__fa_1 _43347_ (.A(_22390_),
    .B(_22369_),
    .CIN(_22389_),
    .COUT(_22391_),
    .SUM(_22392_));
 sky130_fd_sc_hd__fa_1 _43348_ (.A(_02451_),
    .B(_22372_),
    .CIN(_22392_),
    .COUT(_22393_),
    .SUM(_22394_));
 sky130_fd_sc_hd__fa_1 _43349_ (.A(_02452_),
    .B(_22374_),
    .CIN(_22394_),
    .COUT(_02453_),
    .SUM(_02454_));
 sky130_fd_sc_hd__fa_1 _43350_ (.A(_02456_),
    .B(_02457_),
    .CIN(_02458_),
    .COUT(_02459_),
    .SUM(_02460_));
 sky130_fd_sc_hd__fa_1 _43351_ (.A(_02461_),
    .B(_02462_),
    .CIN(_02463_),
    .COUT(_02464_),
    .SUM(_02465_));
 sky130_fd_sc_hd__fa_1 _43352_ (.A(_02466_),
    .B(_02467_),
    .CIN(_02468_),
    .COUT(_22395_),
    .SUM(_22396_));
 sky130_fd_sc_hd__fa_1 _43353_ (.A(_02469_),
    .B(_02470_),
    .CIN(_02448_),
    .COUT(_22397_),
    .SUM(_22398_));
 sky130_fd_sc_hd__fa_1 _43354_ (.A(_22398_),
    .B(_22376_),
    .CIN(_22396_),
    .COUT(_22399_),
    .SUM(_22400_));
 sky130_fd_sc_hd__fa_1 _43355_ (.A(_22378_),
    .B(_02424_),
    .CIN(_02399_),
    .COUT(_22401_),
    .SUM(_22402_));
 sky130_fd_sc_hd__fa_1 _43356_ (.A(_22402_),
    .B(_22380_),
    .CIN(_22400_),
    .COUT(_22403_),
    .SUM(_22404_));
 sky130_fd_sc_hd__fa_1 _43357_ (.A(_22382_),
    .B(_02369_),
    .CIN(_02339_),
    .COUT(_22405_),
    .SUM(_22406_));
 sky130_fd_sc_hd__fa_1 _43358_ (.A(_22406_),
    .B(_22384_),
    .CIN(_22404_),
    .COUT(_22407_),
    .SUM(_22408_));
 sky130_fd_sc_hd__fa_1 _43359_ (.A(_22386_),
    .B(net788),
    .CIN(net789),
    .COUT(_02471_),
    .SUM(_22409_));
 sky130_fd_sc_hd__fa_1 _43360_ (.A(_22409_),
    .B(_22388_),
    .CIN(_22408_),
    .COUT(_22410_),
    .SUM(_22411_));
 sky130_fd_sc_hd__fa_1 _43361_ (.A(_02472_),
    .B(_22391_),
    .CIN(_22411_),
    .COUT(_22412_),
    .SUM(_22413_));
 sky130_fd_sc_hd__fa_1 _43362_ (.A(_02473_),
    .B(_22393_),
    .CIN(_22413_),
    .COUT(_02474_),
    .SUM(_02475_));
 sky130_fd_sc_hd__fa_1 _43363_ (.A(_02477_),
    .B(_02478_),
    .CIN(_02479_),
    .COUT(_02480_),
    .SUM(_22414_));
 sky130_fd_sc_hd__fa_1 _43364_ (.A(_02481_),
    .B(_02482_),
    .CIN(_02483_),
    .COUT(_22415_),
    .SUM(_22416_));
 sky130_fd_sc_hd__fa_1 _43365_ (.A(_22416_),
    .B(_02484_),
    .CIN(_22414_),
    .COUT(_22417_),
    .SUM(_22418_));
 sky130_fd_sc_hd__fa_1 _43366_ (.A(_02485_),
    .B(_02469_),
    .CIN(_02448_),
    .COUT(_22419_),
    .SUM(_22420_));
 sky130_fd_sc_hd__fa_1 _43367_ (.A(_22420_),
    .B(_22395_),
    .CIN(_22418_),
    .COUT(_22421_),
    .SUM(_22422_));
 sky130_fd_sc_hd__fa_1 _43368_ (.A(_22397_),
    .B(_02424_),
    .CIN(_02399_),
    .COUT(_22423_),
    .SUM(_22424_));
 sky130_fd_sc_hd__fa_1 _43369_ (.A(_22424_),
    .B(_22399_),
    .CIN(_22422_),
    .COUT(_22425_),
    .SUM(_22426_));
 sky130_fd_sc_hd__fa_1 _43370_ (.A(_22401_),
    .B(_02369_),
    .CIN(_02339_),
    .COUT(_22427_),
    .SUM(_22428_));
 sky130_fd_sc_hd__fa_1 _43371_ (.A(_22428_),
    .B(_22403_),
    .CIN(_22426_),
    .COUT(_22429_),
    .SUM(_22430_));
 sky130_fd_sc_hd__fa_1 _43372_ (.A(_22405_),
    .B(net788),
    .CIN(net789),
    .COUT(_02486_),
    .SUM(_22431_));
 sky130_fd_sc_hd__fa_1 _43373_ (.A(_22431_),
    .B(_22407_),
    .CIN(_22430_),
    .COUT(_22432_),
    .SUM(_22433_));
 sky130_fd_sc_hd__fa_1 _43374_ (.A(_02487_),
    .B(_22410_),
    .CIN(_22433_),
    .COUT(_22434_),
    .SUM(_22435_));
 sky130_fd_sc_hd__fa_1 _43375_ (.A(_02488_),
    .B(_22412_),
    .CIN(_22435_),
    .COUT(_02489_),
    .SUM(_02490_));
 sky130_fd_sc_hd__fa_1 _43376_ (.A(_02492_),
    .B(_02493_),
    .CIN(_02494_),
    .COUT(_02495_),
    .SUM(_22436_));
 sky130_fd_sc_hd__fa_1 _43377_ (.A(_02496_),
    .B(_02497_),
    .CIN(_02461_),
    .COUT(_02498_),
    .SUM(_02499_));
 sky130_fd_sc_hd__fa_1 _43378_ (.A(_02499_),
    .B(_02500_),
    .CIN(_22436_),
    .COUT(_22437_),
    .SUM(_02501_));
 sky130_fd_sc_hd__fa_1 _43379_ (.A(_22415_),
    .B(_02469_),
    .CIN(_02448_),
    .COUT(_02503_),
    .SUM(_22438_));
 sky130_fd_sc_hd__fa_1 _43380_ (.A(_22438_),
    .B(_22417_),
    .CIN(_02504_),
    .COUT(_22439_),
    .SUM(_22440_));
 sky130_fd_sc_hd__fa_1 _43381_ (.A(_22419_),
    .B(_02424_),
    .CIN(_02399_),
    .COUT(_22441_),
    .SUM(_22442_));
 sky130_fd_sc_hd__fa_1 _43382_ (.A(_22442_),
    .B(_22421_),
    .CIN(_22440_),
    .COUT(_22443_),
    .SUM(_22444_));
 sky130_fd_sc_hd__fa_1 _43383_ (.A(_22423_),
    .B(_02369_),
    .CIN(_02339_),
    .COUT(_22445_),
    .SUM(_22446_));
 sky130_fd_sc_hd__fa_1 _43384_ (.A(_22446_),
    .B(_22425_),
    .CIN(_22444_),
    .COUT(_22447_),
    .SUM(_22448_));
 sky130_fd_sc_hd__fa_1 _43385_ (.A(_22427_),
    .B(net788),
    .CIN(net789),
    .COUT(_02505_),
    .SUM(_22449_));
 sky130_fd_sc_hd__fa_1 _43386_ (.A(_22449_),
    .B(_22429_),
    .CIN(_22448_),
    .COUT(_22450_),
    .SUM(_22451_));
 sky130_fd_sc_hd__fa_1 _43387_ (.A(_02506_),
    .B(_22432_),
    .CIN(_22451_),
    .COUT(_22452_),
    .SUM(_22453_));
 sky130_fd_sc_hd__fa_1 _43388_ (.A(_02507_),
    .B(_22434_),
    .CIN(_22453_),
    .COUT(_02508_),
    .SUM(_02509_));
 sky130_fd_sc_hd__fa_1 _43389_ (.A(_02511_),
    .B(_02512_),
    .CIN(_02513_),
    .COUT(_02514_),
    .SUM(_22454_));
 sky130_fd_sc_hd__fa_1 _43390_ (.A(_02515_),
    .B(_22454_),
    .CIN(_02502_),
    .COUT(_02516_),
    .SUM(_02517_));
 sky130_fd_sc_hd__fa_1 _43391_ (.A(_02518_),
    .B(_02469_),
    .CIN(_02448_),
    .COUT(_02519_),
    .SUM(_02520_));
 sky130_fd_sc_hd__fa_1 _43392_ (.A(_02521_),
    .B(_22437_),
    .CIN(_02522_),
    .COUT(_02523_),
    .SUM(_02524_));
 sky130_fd_sc_hd__fa_1 _43393_ (.A(_02525_),
    .B(_02397_),
    .CIN(_02398_),
    .COUT(_02526_),
    .SUM(_02527_));
 sky130_fd_sc_hd__fa_1 _43394_ (.A(_02528_),
    .B(_22439_),
    .CIN(_02529_),
    .COUT(_02530_),
    .SUM(_22455_));
 sky130_fd_sc_hd__fa_1 _43395_ (.A(_22441_),
    .B(_02369_),
    .CIN(_02339_),
    .COUT(_02531_),
    .SUM(_22456_));
 sky130_fd_sc_hd__fa_1 _43396_ (.A(_22456_),
    .B(_22443_),
    .CIN(_22455_),
    .COUT(_02532_),
    .SUM(_22457_));
 sky130_fd_sc_hd__fa_1 _43397_ (.A(_22445_),
    .B(net788),
    .CIN(net789),
    .COUT(_02533_),
    .SUM(_22458_));
 sky130_fd_sc_hd__fa_1 _43398_ (.A(_22458_),
    .B(_22447_),
    .CIN(_22457_),
    .COUT(_02534_),
    .SUM(_22459_));
 sky130_fd_sc_hd__fa_1 _43399_ (.A(_02535_),
    .B(_22450_),
    .CIN(_22459_),
    .COUT(_02536_),
    .SUM(_22460_));
 sky130_fd_sc_hd__fa_1 _43400_ (.A(_02537_),
    .B(_22452_),
    .CIN(_22460_),
    .COUT(_02538_),
    .SUM(_02539_));
 sky130_fd_sc_hd__fa_1 _43401_ (.A(\inst$top.soc.cpu.divider.remainder[0] ),
    .B(_02541_),
    .CIN(_02542_),
    .COUT(_02543_),
    .SUM(_02544_));
 sky130_fd_sc_hd__fa_1 _43402_ (.A(net884),
    .B(\inst$top.soc.cpu.sink__payload$6[3] ),
    .CIN(_02545_),
    .COUT(_02546_),
    .SUM(\inst$top.soc.cpu.d_branch_target[3] ));
 sky130_fd_sc_hd__fa_1 _43403_ (.A(_02547_),
    .B(_22461_),
    .CIN(_22462_),
    .COUT(_02548_),
    .SUM(\inst$top.soc.cpu.multiplier.x_prod[6] ));
 sky130_fd_sc_hd__ha_1 _43404_ (.A(_02549_),
    .B(_21755_),
    .COUT(_01787_),
    .SUM(_02550_));
 sky130_fd_sc_hd__ha_1 _43405_ (.A(_02551_),
    .B(_02552_),
    .COUT(_02553_),
    .SUM(_02554_));
 sky130_fd_sc_hd__ha_1 _43406_ (.A(net819),
    .B(_21800_),
    .COUT(_01835_),
    .SUM(_02556_));
 sky130_fd_sc_hd__ha_1 _43407_ (.A(_02557_),
    .B(_02558_),
    .COUT(_02559_),
    .SUM(_02560_));
 sky130_fd_sc_hd__ha_1 _43408_ (.A(_02561_),
    .B(net819),
    .COUT(_01888_),
    .SUM(_02562_));
 sky130_fd_sc_hd__ha_1 _43409_ (.A(_02563_),
    .B(_02564_),
    .COUT(_02565_),
    .SUM(_02566_));
 sky130_fd_sc_hd__ha_1 _43410_ (.A(_02567_),
    .B(net819),
    .COUT(_01941_),
    .SUM(_02568_));
 sky130_fd_sc_hd__ha_1 _43411_ (.A(_02569_),
    .B(_02570_),
    .COUT(_02571_),
    .SUM(_02572_));
 sky130_fd_sc_hd__ha_1 _43412_ (.A(_02573_),
    .B(net819),
    .COUT(_01989_),
    .SUM(_02574_));
 sky130_fd_sc_hd__ha_1 _43413_ (.A(_02575_),
    .B(_02576_),
    .COUT(_02577_),
    .SUM(_02578_));
 sky130_fd_sc_hd__ha_1 _43414_ (.A(_02579_),
    .B(net819),
    .COUT(_02036_),
    .SUM(_02580_));
 sky130_fd_sc_hd__ha_1 _43415_ (.A(_02581_),
    .B(_02582_),
    .COUT(_02583_),
    .SUM(_02584_));
 sky130_fd_sc_hd__ha_1 _43416_ (.A(_02585_),
    .B(net819),
    .COUT(_02082_),
    .SUM(_02586_));
 sky130_fd_sc_hd__ha_1 _43417_ (.A(_02587_),
    .B(_02588_),
    .COUT(_02589_),
    .SUM(_02590_));
 sky130_fd_sc_hd__ha_1 _43418_ (.A(_02591_),
    .B(net820),
    .COUT(_02121_),
    .SUM(_02592_));
 sky130_fd_sc_hd__ha_1 _43419_ (.A(_02593_),
    .B(_02594_),
    .COUT(_02595_),
    .SUM(_02596_));
 sky130_fd_sc_hd__ha_1 _43420_ (.A(_02597_),
    .B(net819),
    .COUT(_02151_),
    .SUM(_02598_));
 sky130_fd_sc_hd__ha_1 _43421_ (.A(_02599_),
    .B(_02600_),
    .COUT(_02601_),
    .SUM(_02602_));
 sky130_fd_sc_hd__ha_1 _43422_ (.A(_02604_),
    .B(net819),
    .COUT(_02184_),
    .SUM(_02605_));
 sky130_fd_sc_hd__ha_1 _43423_ (.A(_02606_),
    .B(_02607_),
    .COUT(_02608_),
    .SUM(_02609_));
 sky130_fd_sc_hd__ha_1 _43424_ (.A(_02610_),
    .B(net819),
    .COUT(_02211_),
    .SUM(_02611_));
 sky130_fd_sc_hd__ha_1 _43425_ (.A(_02612_),
    .B(_02613_),
    .COUT(_02614_),
    .SUM(_02615_));
 sky130_fd_sc_hd__ha_1 _43426_ (.A(_02617_),
    .B(net819),
    .COUT(_02245_),
    .SUM(_02618_));
 sky130_fd_sc_hd__ha_1 _43427_ (.A(_02619_),
    .B(_02620_),
    .COUT(_02621_),
    .SUM(_02622_));
 sky130_fd_sc_hd__ha_1 _43428_ (.A(_02623_),
    .B(net818),
    .COUT(_02284_),
    .SUM(_02624_));
 sky130_fd_sc_hd__ha_1 _43429_ (.A(_02625_),
    .B(_02626_),
    .COUT(_02627_),
    .SUM(_02628_));
 sky130_fd_sc_hd__ha_1 _43430_ (.A(_02629_),
    .B(net818),
    .COUT(_02318_),
    .SUM(_02630_));
 sky130_fd_sc_hd__ha_1 _43431_ (.A(_02631_),
    .B(_02632_),
    .COUT(_02633_),
    .SUM(_02634_));
 sky130_fd_sc_hd__ha_1 _43432_ (.A(_02635_),
    .B(net820),
    .COUT(_02345_),
    .SUM(_02636_));
 sky130_fd_sc_hd__ha_1 _43433_ (.A(_02637_),
    .B(_02638_),
    .COUT(_02639_),
    .SUM(_02640_));
 sky130_fd_sc_hd__ha_1 _43434_ (.A(_02642_),
    .B(net820),
    .COUT(_02375_),
    .SUM(_02643_));
 sky130_fd_sc_hd__ha_1 _43435_ (.A(_02644_),
    .B(_02645_),
    .COUT(_02646_),
    .SUM(_02647_));
 sky130_fd_sc_hd__ha_1 _43436_ (.A(_02648_),
    .B(net820),
    .COUT(_02405_),
    .SUM(_02649_));
 sky130_fd_sc_hd__ha_1 _43437_ (.A(_02650_),
    .B(_02651_),
    .COUT(_02652_),
    .SUM(_02653_));
 sky130_fd_sc_hd__ha_1 _43438_ (.A(_02654_),
    .B(net818),
    .COUT(_02430_),
    .SUM(_02655_));
 sky130_fd_sc_hd__ha_1 _43439_ (.A(_02656_),
    .B(_02657_),
    .COUT(_02658_),
    .SUM(_02659_));
 sky130_fd_sc_hd__ha_1 _43440_ (.A(_02660_),
    .B(net818),
    .COUT(_02455_),
    .SUM(_02661_));
 sky130_fd_sc_hd__ha_1 _43441_ (.A(_02662_),
    .B(_02663_),
    .COUT(_02664_),
    .SUM(_02665_));
 sky130_fd_sc_hd__ha_1 _43442_ (.A(_02666_),
    .B(net818),
    .COUT(_02476_),
    .SUM(_02667_));
 sky130_fd_sc_hd__ha_1 _43443_ (.A(_02668_),
    .B(_02669_),
    .COUT(_02670_),
    .SUM(_02671_));
 sky130_fd_sc_hd__ha_1 _43444_ (.A(_02672_),
    .B(net818),
    .COUT(_02491_),
    .SUM(_02673_));
 sky130_fd_sc_hd__ha_1 _43445_ (.A(_02674_),
    .B(_02675_),
    .COUT(_02676_),
    .SUM(_02677_));
 sky130_fd_sc_hd__ha_1 _43446_ (.A(_02679_),
    .B(net818),
    .COUT(_02510_),
    .SUM(_02680_));
 sky130_fd_sc_hd__ha_1 _43447_ (.A(_02681_),
    .B(_02682_),
    .COUT(_02683_),
    .SUM(_02684_));
 sky130_fd_sc_hd__ha_1 _43448_ (.A(_02685_),
    .B(net818),
    .COUT(_02540_),
    .SUM(_02686_));
 sky130_fd_sc_hd__ha_1 _43449_ (.A(_02687_),
    .B(_02688_),
    .COUT(_02689_),
    .SUM(_02690_));
 sky130_fd_sc_hd__ha_1 _43450_ (.A(_02692_),
    .B(net818),
    .COUT(_02693_),
    .SUM(_02694_));
 sky130_fd_sc_hd__ha_1 _43451_ (.A(_02695_),
    .B(_02696_),
    .COUT(_02697_),
    .SUM(_02698_));
 sky130_fd_sc_hd__ha_1 _43452_ (.A(net1682),
    .B(net1697),
    .COUT(_02700_),
    .SUM(_02701_));
 sky130_fd_sc_hd__ha_1 _43453_ (.A(_02702_),
    .B(_02703_),
    .COUT(_02704_),
    .SUM(_02705_));
 sky130_fd_sc_hd__ha_1 _43454_ (.A(_02706_),
    .B(_02707_),
    .COUT(_02708_),
    .SUM(_02709_));
 sky130_fd_sc_hd__ha_1 _43455_ (.A(_02710_),
    .B(_02711_),
    .COUT(_02712_),
    .SUM(_02713_));
 sky130_fd_sc_hd__ha_1 _43456_ (.A(_02714_),
    .B(_02715_),
    .COUT(_02716_),
    .SUM(_02717_));
 sky130_fd_sc_hd__ha_1 _43457_ (.A(_02714_),
    .B(_02715_),
    .COUT(_02718_),
    .SUM(_22463_));
 sky130_fd_sc_hd__ha_1 _43458_ (.A(_02719_),
    .B(_02720_),
    .COUT(_02721_),
    .SUM(_02722_));
 sky130_fd_sc_hd__ha_1 _43459_ (.A(_02723_),
    .B(_02724_),
    .COUT(_02725_),
    .SUM(_02726_));
 sky130_fd_sc_hd__ha_1 _43460_ (.A(_02727_),
    .B(_02728_),
    .COUT(_02729_),
    .SUM(_02730_));
 sky130_fd_sc_hd__ha_1 _43461_ (.A(\inst$top.soc.spiflash.ctrl.o_data_count[0] ),
    .B(\inst$top.soc.spiflash.ctrl.o_data_count[1] ),
    .COUT(_02731_),
    .SUM(_22464_));
 sky130_fd_sc_hd__ha_1 _43462_ (.A(_02732_),
    .B(_02733_),
    .COUT(_02734_),
    .SUM(_02735_));
 sky130_fd_sc_hd__ha_1 _43463_ (.A(_02732_),
    .B(\inst$top.soc.spiflash.ctrl.i_data_count[1] ),
    .COUT(_02736_),
    .SUM(_22465_));
 sky130_fd_sc_hd__ha_1 _43464_ (.A(\inst$top.soc.spiflash.ctrl.i_data_count[0] ),
    .B(_02733_),
    .COUT(_02737_),
    .SUM(_22466_));
 sky130_fd_sc_hd__ha_1 _43465_ (.A(\inst$top.soc.spiflash.ctrl.i_data_count[0] ),
    .B(\inst$top.soc.spiflash.ctrl.i_data_count[1] ),
    .COUT(_02738_),
    .SUM(_22467_));
 sky130_fd_sc_hd__ha_1 _43466_ (.A(_02739_),
    .B(_02740_),
    .COUT(_02741_),
    .SUM(_02742_));
 sky130_fd_sc_hd__ha_1 _43467_ (.A(\inst$top.soc.spiflash.phy.io_clocker.timer[0] ),
    .B(_02740_),
    .COUT(_02743_),
    .SUM(_22468_));
 sky130_fd_sc_hd__ha_1 _43468_ (.A(_02744_),
    .B(_02745_),
    .COUT(_02746_),
    .SUM(_02747_));
 sky130_fd_sc_hd__ha_1 _43469_ (.A(net2579),
    .B(net2578),
    .COUT(_02748_),
    .SUM(_22469_));
 sky130_fd_sc_hd__ha_1 _43470_ (.A(\inst$top.soc.spiflash.phy.deframer.cycle[0] ),
    .B(\inst$top.soc.spiflash.phy.deframer.cycle[1] ),
    .COUT(_02749_),
    .SUM(_02750_));
 sky130_fd_sc_hd__ha_1 _43471_ (.A(\inst$top.soc.cpu.divider.remainder[30] ),
    .B(_02751_),
    .COUT(_02752_),
    .SUM(_02753_));
 sky130_fd_sc_hd__ha_1 _43472_ (.A(\inst$top.soc.cpu.divider.remainder[29] ),
    .B(_02754_),
    .COUT(_02755_),
    .SUM(_02756_));
 sky130_fd_sc_hd__ha_1 _43473_ (.A(\inst$top.soc.cpu.divider.remainder[28] ),
    .B(_02757_),
    .COUT(_02758_),
    .SUM(_02759_));
 sky130_fd_sc_hd__ha_1 _43474_ (.A(\inst$top.soc.cpu.divider.remainder[27] ),
    .B(_02760_),
    .COUT(_02761_),
    .SUM(_02762_));
 sky130_fd_sc_hd__ha_1 _43475_ (.A(\inst$top.soc.cpu.divider.remainder[26] ),
    .B(_02763_),
    .COUT(_02764_),
    .SUM(_02765_));
 sky130_fd_sc_hd__ha_1 _43476_ (.A(\inst$top.soc.cpu.divider.remainder[25] ),
    .B(_02766_),
    .COUT(_02767_),
    .SUM(_02768_));
 sky130_fd_sc_hd__ha_1 _43477_ (.A(\inst$top.soc.cpu.divider.remainder[24] ),
    .B(_02769_),
    .COUT(_02770_),
    .SUM(_02771_));
 sky130_fd_sc_hd__ha_1 _43478_ (.A(\inst$top.soc.cpu.divider.remainder[23] ),
    .B(_02772_),
    .COUT(_02773_),
    .SUM(_02774_));
 sky130_fd_sc_hd__ha_1 _43479_ (.A(\inst$top.soc.cpu.divider.remainder[22] ),
    .B(_02775_),
    .COUT(_02776_),
    .SUM(_02777_));
 sky130_fd_sc_hd__ha_1 _43480_ (.A(\inst$top.soc.cpu.divider.remainder[21] ),
    .B(_02778_),
    .COUT(_02779_),
    .SUM(_02780_));
 sky130_fd_sc_hd__ha_1 _43481_ (.A(\inst$top.soc.cpu.divider.remainder[20] ),
    .B(_02781_),
    .COUT(_02782_),
    .SUM(_02783_));
 sky130_fd_sc_hd__ha_1 _43482_ (.A(\inst$top.soc.cpu.divider.remainder[19] ),
    .B(_02784_),
    .COUT(_02785_),
    .SUM(_02786_));
 sky130_fd_sc_hd__ha_1 _43483_ (.A(\inst$top.soc.cpu.divider.remainder[18] ),
    .B(_02787_),
    .COUT(_02788_),
    .SUM(_02789_));
 sky130_fd_sc_hd__ha_1 _43484_ (.A(\inst$top.soc.cpu.divider.remainder[17] ),
    .B(_02790_),
    .COUT(_02791_),
    .SUM(_02792_));
 sky130_fd_sc_hd__ha_1 _43485_ (.A(\inst$top.soc.cpu.divider.remainder[16] ),
    .B(_02793_),
    .COUT(_02794_),
    .SUM(_02795_));
 sky130_fd_sc_hd__ha_1 _43486_ (.A(\inst$top.soc.cpu.divider.remainder[15] ),
    .B(_02796_),
    .COUT(_02797_),
    .SUM(_02798_));
 sky130_fd_sc_hd__ha_1 _43487_ (.A(\inst$top.soc.cpu.divider.remainder[14] ),
    .B(_02799_),
    .COUT(_02800_),
    .SUM(_02801_));
 sky130_fd_sc_hd__ha_1 _43488_ (.A(\inst$top.soc.cpu.divider.remainder[13] ),
    .B(_02802_),
    .COUT(_02803_),
    .SUM(_02804_));
 sky130_fd_sc_hd__ha_1 _43489_ (.A(\inst$top.soc.cpu.divider.remainder[12] ),
    .B(_02805_),
    .COUT(_02806_),
    .SUM(_02807_));
 sky130_fd_sc_hd__ha_1 _43490_ (.A(\inst$top.soc.cpu.divider.remainder[11] ),
    .B(_02808_),
    .COUT(_02809_),
    .SUM(_02810_));
 sky130_fd_sc_hd__ha_1 _43491_ (.A(\inst$top.soc.cpu.divider.remainder[10] ),
    .B(_02811_),
    .COUT(_02812_),
    .SUM(_02813_));
 sky130_fd_sc_hd__ha_1 _43492_ (.A(\inst$top.soc.cpu.divider.remainder[9] ),
    .B(_02814_),
    .COUT(_02815_),
    .SUM(_02816_));
 sky130_fd_sc_hd__ha_1 _43493_ (.A(\inst$top.soc.cpu.divider.remainder[8] ),
    .B(_02817_),
    .COUT(_02818_),
    .SUM(_02819_));
 sky130_fd_sc_hd__ha_1 _43494_ (.A(\inst$top.soc.cpu.divider.remainder[7] ),
    .B(_02820_),
    .COUT(_02821_),
    .SUM(_02822_));
 sky130_fd_sc_hd__ha_1 _43495_ (.A(\inst$top.soc.cpu.divider.remainder[6] ),
    .B(_02823_),
    .COUT(_02824_),
    .SUM(_02825_));
 sky130_fd_sc_hd__ha_1 _43496_ (.A(\inst$top.soc.cpu.divider.remainder[5] ),
    .B(_02826_),
    .COUT(_02827_),
    .SUM(_02828_));
 sky130_fd_sc_hd__ha_1 _43497_ (.A(\inst$top.soc.cpu.divider.remainder[4] ),
    .B(_02829_),
    .COUT(_02830_),
    .SUM(_02831_));
 sky130_fd_sc_hd__ha_1 _43498_ (.A(\inst$top.soc.cpu.divider.remainder[3] ),
    .B(_02832_),
    .COUT(_02833_),
    .SUM(_02834_));
 sky130_fd_sc_hd__ha_1 _43499_ (.A(\inst$top.soc.cpu.divider.remainder[2] ),
    .B(_02835_),
    .COUT(_02836_),
    .SUM(_02837_));
 sky130_fd_sc_hd__ha_1 _43500_ (.A(\inst$top.soc.cpu.divider.remainder[1] ),
    .B(_02838_),
    .COUT(_02839_),
    .SUM(_02840_));
 sky130_fd_sc_hd__ha_1 _43501_ (.A(\inst$top.soc.cpu.divider.remainder[0] ),
    .B(_02541_),
    .COUT(_02841_),
    .SUM(_02842_));
 sky130_fd_sc_hd__ha_1 _43502_ (.A(net1691),
    .B(net1706),
    .COUT(_02844_),
    .SUM(_02845_));
 sky130_fd_sc_hd__ha_1 _43503_ (.A(_02846_),
    .B(_02847_),
    .COUT(_02848_),
    .SUM(_02849_));
 sky130_fd_sc_hd__ha_1 _43504_ (.A(_02850_),
    .B(\inst$top.soc.cpu.divider.divisor[0] ),
    .COUT(_02851_),
    .SUM(_02852_));
 sky130_fd_sc_hd__ha_1 _43505_ (.A(_02853_),
    .B(_02854_),
    .COUT(_02855_),
    .SUM(_02856_));
 sky130_fd_sc_hd__ha_1 _43506_ (.A(_02857_),
    .B(_02858_),
    .COUT(_02859_),
    .SUM(_02860_));
 sky130_fd_sc_hd__ha_1 _43507_ (.A(_02861_),
    .B(\inst$top.soc.cpu.d.sink__payload$6.branch_predict_taken ),
    .COUT(_02862_),
    .SUM(_02863_));
 sky130_fd_sc_hd__ha_1 _43508_ (.A(\inst$top.soc.cpu.d.sink__payload$6.branch_taken ),
    .B(_02864_),
    .COUT(_02865_),
    .SUM(_22470_));
 sky130_fd_sc_hd__ha_1 _43509_ (.A(\inst$top.soc.cpu.sink__payload[2] ),
    .B(\inst$top.soc.cpu.sink__payload[3] ),
    .COUT(_02866_),
    .SUM(_02867_));
 sky130_fd_sc_hd__ha_1 _43510_ (.A(_02868_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__2._storage[1] ),
    .COUT(_02869_),
    .SUM(_02870_));
 sky130_fd_sc_hd__ha_1 _43511_ (.A(_02871_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__0._storage[1] ),
    .COUT(_02872_),
    .SUM(_02873_));
 sky130_fd_sc_hd__ha_1 _43512_ (.A(_02874_),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__3._storage[1] ),
    .COUT(_02875_),
    .SUM(_02876_));
 sky130_fd_sc_hd__ha_1 _43513_ (.A(_02877_),
    .B(_02878_),
    .COUT(_02879_),
    .SUM(_02880_));
 sky130_fd_sc_hd__ha_1 _43514_ (.A(_02877_),
    .B(\inst$top.soc.uart_0._phy.rx.lower.fsm_state[1] ),
    .COUT(_02881_),
    .SUM(_22471_));
 sky130_fd_sc_hd__ha_1 _43515_ (.A(\inst$top.soc.uart_0._phy.rx.lower.fsm_state[0] ),
    .B(_02878_),
    .COUT(_02882_),
    .SUM(_22472_));
 sky130_fd_sc_hd__ha_1 _43516_ (.A(\inst$top.soc.uart_0._phy.rx.lower.fsm_state[0] ),
    .B(\inst$top.soc.uart_0._phy.rx.lower.fsm_state[1] ),
    .COUT(_02883_),
    .SUM(_22473_));
 sky130_fd_sc_hd__ha_1 _43517_ (.A(_02884_),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__1._storage[1] ),
    .COUT(_02885_),
    .SUM(_02886_));
 sky130_fd_sc_hd__ha_1 _43518_ (.A(_02887_),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__0._storage[1] ),
    .COUT(_02888_),
    .SUM(_02889_));
 sky130_fd_sc_hd__ha_1 _43519_ (.A(_02890_),
    .B(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__2._storage[1] ),
    .COUT(_02891_),
    .SUM(_02892_));
 sky130_fd_sc_hd__ha_1 _43520_ (.A(_02893_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__1._storage[1] ),
    .COUT(_02894_),
    .SUM(_02895_));
 sky130_fd_sc_hd__ha_1 _43521_ (.A(_02896_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__3._storage[1] ),
    .COUT(_02897_),
    .SUM(_02898_));
 sky130_fd_sc_hd__ha_1 _43522_ (.A(_02899_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__7._storage[1] ),
    .COUT(_02900_),
    .SUM(_02901_));
 sky130_fd_sc_hd__ha_1 _43523_ (.A(_02902_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__6._storage[1] ),
    .COUT(_02903_),
    .SUM(_02904_));
 sky130_fd_sc_hd__ha_1 _43524_ (.A(_02905_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__5._storage[1] ),
    .COUT(_02906_),
    .SUM(_02907_));
 sky130_fd_sc_hd__ha_1 _43525_ (.A(_02908_),
    .B(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__4._storage[1] ),
    .COUT(_02909_),
    .SUM(_02910_));
 sky130_fd_sc_hd__ha_1 _43526_ (.A(_06044_),
    .B(\inst$top.soc.cpu.sink__payload$6[2] ),
    .COUT(_02545_),
    .SUM(\inst$top.soc.cpu.d_branch_target[2] ));
 sky130_fd_sc_hd__ha_1 _43527_ (.A(_02912_),
    .B(_02913_),
    .COUT(_22474_),
    .SUM(\inst$top.soc.cpu.multiplier.x_prod[1] ));
 sky130_fd_sc_hd__ha_1 _43528_ (.A(_02914_),
    .B(_22474_),
    .COUT(_22475_),
    .SUM(\inst$top.soc.cpu.multiplier.x_prod[2] ));
 sky130_fd_sc_hd__ha_1 _43529_ (.A(_22476_),
    .B(_22475_),
    .COUT(_22477_),
    .SUM(\inst$top.soc.cpu.multiplier.x_prod[3] ));
 sky130_fd_sc_hd__ha_1 _43530_ (.A(_22477_),
    .B(_22478_),
    .COUT(_22479_),
    .SUM(\inst$top.soc.cpu.multiplier.x_prod[4] ));
 sky130_fd_sc_hd__ha_1 _43531_ (.A(_22479_),
    .B(_22480_),
    .COUT(_02547_),
    .SUM(\inst$top.soc.cpu.multiplier.x_prod[5] ));
 sky130_fd_sc_hd__ha_1 _43532_ (.A(net1734),
    .B(net1453),
    .COUT(_02641_),
    .SUM(_02918_));
 sky130_fd_sc_hd__ha_1 _43533_ (.A(net1739),
    .B(net1482),
    .COUT(_02921_),
    .SUM(_02922_));
 sky130_fd_sc_hd__ha_1 _43534_ (.A(net1480),
    .B(net1482),
    .COUT(_02691_),
    .SUM(_22481_));
 sky130_fd_sc_hd__ha_1 _43535_ (.A(net1480),
    .B(net1222),
    .COUT(_02925_),
    .SUM(_22482_));
 sky130_fd_sc_hd__ha_1 _43536_ (.A(net1473),
    .B(net1476),
    .COUT(_02678_),
    .SUM(_02928_));
 sky130_fd_sc_hd__ha_1 _43537_ (.A(net1219),
    .B(net1475),
    .COUT(_02930_),
    .SUM(_22483_));
 sky130_fd_sc_hd__ha_1 _43538_ (.A(net1465),
    .B(net1467),
    .COUT(_02438_),
    .SUM(_02933_));
 sky130_fd_sc_hd__ha_1 _43539_ (.A(net1218),
    .B(net1469),
    .COUT(_02935_),
    .SUM(_22484_));
 sky130_fd_sc_hd__ha_1 _43540_ (.A(net1457),
    .B(net1460),
    .COUT(_02383_),
    .SUM(_02938_));
 sky130_fd_sc_hd__ha_1 _43541_ (.A(net1217),
    .B(net1460),
    .COUT(_02940_),
    .SUM(_22485_));
 sky130_fd_sc_hd__ha_1 _43542_ (.A(net1264),
    .B(net1453),
    .COUT(_02942_),
    .SUM(_02943_));
 sky130_fd_sc_hd__ha_1 _43543_ (.A(net1265),
    .B(net1253),
    .COUT(_02946_),
    .SUM(_02947_));
 sky130_fd_sc_hd__ha_1 _43544_ (.A(net1730),
    .B(net1253),
    .COUT(_02257_),
    .SUM(_22486_));
 sky130_fd_sc_hd__ha_1 _43545_ (.A(net1268),
    .B(net1256),
    .COUT(_02951_),
    .SUM(_02952_));
 sky130_fd_sc_hd__ha_1 _43546_ (.A(net1726),
    .B(net1257),
    .COUT(_02616_),
    .SUM(_22487_));
 sky130_fd_sc_hd__ha_1 _43547_ (.A(net1450),
    .B(net1272),
    .COUT(_02956_),
    .SUM(_02957_));
 sky130_fd_sc_hd__ha_1 _43548_ (.A(net1216),
    .B(net1272),
    .COUT(_02603_),
    .SUM(_22488_));
 sky130_fd_sc_hd__ha_2 _43549_ (.A(net1447),
    .B(net1273),
    .COUT(_02053_),
    .SUM(_02961_));
 sky130_fd_sc_hd__ha_1 _43550_ (.A(net1213),
    .B(net1276),
    .COUT(_02963_),
    .SUM(_22489_));
 sky130_fd_sc_hd__ha_1 _43551_ (.A(net1442),
    .B(net1258),
    .COUT(_01958_),
    .SUM(_02966_));
 sky130_fd_sc_hd__ha_1 _43552_ (.A(net1211),
    .B(net1260),
    .COUT(_02968_),
    .SUM(_22490_));
 sky130_fd_sc_hd__ha_1 _43553_ (.A(net1438),
    .B(net1281),
    .COUT(_02971_),
    .SUM(_02972_));
 sky130_fd_sc_hd__ha_1 _43554_ (.A(net1209),
    .B(net1278),
    .COUT(_01850_),
    .SUM(_22491_));
 sky130_fd_sc_hd__ha_1 _43555_ (.A(net1134),
    .B(net1283),
    .COUT(_02555_),
    .SUM(_02976_));
 sky130_fd_sc_hd__ha_1 _43556_ (.A(_20003_),
    .B(net1285),
    .COUT(_02978_),
    .SUM(_22492_));
 sky130_fd_sc_hd__ha_1 _43557_ (.A(net1434),
    .B(net1288),
    .COUT(_02981_),
    .SUM(_02982_));
 sky130_fd_sc_hd__ha_1 _43558_ (.A(_02983_),
    .B(net1290),
    .COUT(_02984_),
    .SUM(_22493_));
 sky130_fd_sc_hd__ha_1 _43559_ (.A(net1722),
    .B(net1295),
    .COUT(_02987_),
    .SUM(_02988_));
 sky130_fd_sc_hd__ha_1 _43560_ (.A(net1431),
    .B(net1292),
    .COUT(_01539_),
    .SUM(_22494_));
 sky130_fd_sc_hd__ha_1 _43561_ (.A(net1719),
    .B(net1299),
    .COUT(_02992_),
    .SUM(_02993_));
 sky130_fd_sc_hd__ha_1 _43562_ (.A(net1428),
    .B(net1296),
    .COUT(_01428_),
    .SUM(_22495_));
 sky130_fd_sc_hd__ha_1 _43563_ (.A(net1715),
    .B(net1302),
    .COUT(_02997_),
    .SUM(_02998_));
 sky130_fd_sc_hd__ha_1 _43564_ (.A(net1427),
    .B(net1300),
    .COUT(_03000_),
    .SUM(_22496_));
 sky130_fd_sc_hd__ha_1 _43565_ (.A(net1712),
    .B(net1307),
    .COUT(_03003_),
    .SUM(_03004_));
 sky130_fd_sc_hd__ha_1 _43566_ (.A(net1425),
    .B(net1307),
    .COUT(_03006_),
    .SUM(_22497_));
 sky130_fd_sc_hd__ha_1 _43567_ (.A(net1423),
    .B(net1311),
    .COUT(_03009_),
    .SUM(_03010_));
 sky130_fd_sc_hd__ha_1 _43568_ (.A(_03011_),
    .B(net1312),
    .COUT(_03012_),
    .SUM(_22498_));
 sky130_fd_sc_hd__ha_1 _43569_ (.A(net1419),
    .B(net1316),
    .COUT(_03015_),
    .SUM(_03016_));
 sky130_fd_sc_hd__ha_1 _43570_ (.A(_03017_),
    .B(net1317),
    .COUT(_03018_),
    .SUM(_22499_));
 sky130_fd_sc_hd__ha_1 _43571_ (.A(net1318),
    .B(net1322),
    .COUT(_03021_),
    .SUM(_03022_));
 sky130_fd_sc_hd__ha_1 _43572_ (.A(net1414),
    .B(net1321),
    .COUT(_00826_),
    .SUM(_22500_));
 sky130_fd_sc_hd__ha_1 _43573_ (.A(net1323),
    .B(net1327),
    .COUT(_03026_),
    .SUM(_03027_));
 sky130_fd_sc_hd__ha_1 _43574_ (.A(net1410),
    .B(net1326),
    .COUT(_03029_),
    .SUM(_22501_));
 sky130_fd_sc_hd__ha_1 _43575_ (.A(net1407),
    .B(net1331),
    .COUT(_03032_),
    .SUM(_03033_));
 sky130_fd_sc_hd__ha_1 _43576_ (.A(net1206),
    .B(net1330),
    .COUT(_03035_),
    .SUM(_22502_));
 sky130_fd_sc_hd__ha_1 _43577_ (.A(net1709),
    .B(net1336),
    .COUT(_03038_),
    .SUM(_03039_));
 sky130_fd_sc_hd__ha_1 _43578_ (.A(net1403),
    .B(net1335),
    .COUT(_00531_),
    .SUM(_22503_));
 sky130_fd_sc_hd__ha_1 _43579_ (.A(net1399),
    .B(net1341),
    .COUT(_03043_),
    .SUM(_03044_));
 sky130_fd_sc_hd__ha_1 _43580_ (.A(_03045_),
    .B(net1341),
    .COUT(_00465_),
    .SUM(_22504_));
 sky130_fd_sc_hd__ha_1 _43581_ (.A(net3043),
    .B(net1345),
    .COUT(_03048_),
    .SUM(_03049_));
 sky130_fd_sc_hd__ha_1 _43582_ (.A(net1398),
    .B(net1346),
    .COUT(_00391_),
    .SUM(_22505_));
 sky130_fd_sc_hd__ha_1 _43583_ (.A(net1166),
    .B(net1350),
    .COUT(_03053_),
    .SUM(_03054_));
 sky130_fd_sc_hd__ha_1 _43584_ (.A(net1397),
    .B(net1350),
    .COUT(_03056_),
    .SUM(_22506_));
 sky130_fd_sc_hd__ha_1 _43585_ (.A(net1172),
    .B(net1355),
    .COUT(_03059_),
    .SUM(_03060_));
 sky130_fd_sc_hd__ha_1 _43586_ (.A(net1396),
    .B(net1355),
    .COUT(_00273_),
    .SUM(_22507_));
 sky130_fd_sc_hd__ha_1 _43587_ (.A(net1197),
    .B(net1357),
    .COUT(_03064_),
    .SUM(_03065_));
 sky130_fd_sc_hd__ha_1 _43588_ (.A(net1077),
    .B(net1356),
    .COUT(_00230_),
    .SUM(_22508_));
 sky130_fd_sc_hd__ha_1 _43589_ (.A(net1174),
    .B(net1361),
    .COUT(_03069_),
    .SUM(_03070_));
 sky130_fd_sc_hd__ha_1 _43590_ (.A(net1394),
    .B(net1361),
    .COUT(_03072_),
    .SUM(_22509_));
 sky130_fd_sc_hd__ha_1 _43591_ (.A(net1182),
    .B(net1153),
    .COUT(_03075_),
    .SUM(_03076_));
 sky130_fd_sc_hd__ha_1 _43592_ (.A(net1389),
    .B(net1153),
    .COUT(_03078_),
    .SUM(_22510_));
 sky130_fd_sc_hd__ha_1 _43593_ (.A(net1698),
    .B(net1262),
    .COUT(_03079_),
    .SUM(_03080_));
 sky130_fd_sc_hd__ha_1 _43594_ (.A(net1385),
    .B(net1262),
    .COUT(_03081_),
    .SUM(_22511_));
 sky130_fd_sc_hd__ha_1 _43595_ (.A(net1251),
    .B(_03082_),
    .COUT(\inst$top.soc.cpu.multiplier.x_prod[0] ),
    .SUM(_03083_));
 sky130_fd_sc_hd__ha_1 _43596_ (.A(net1251),
    .B(net1692),
    .COUT(_00169_),
    .SUM(_22512_));
 sky130_fd_sc_hd__ha_1 _43597_ (.A(_03084_),
    .B(_03085_),
    .COUT(_03086_),
    .SUM(_03087_));
 sky130_fd_sc_hd__ha_1 _43598_ (.A(_03088_),
    .B(_03089_),
    .COUT(_03090_),
    .SUM(_22513_));
 sky130_fd_sc_hd__ha_1 _43599_ (.A(_03091_),
    .B(_03092_),
    .COUT(_03093_),
    .SUM(_03094_));
 sky130_fd_sc_hd__ha_1 _43600_ (.A(_03095_),
    .B(_03096_),
    .COUT(_03097_),
    .SUM(_22514_));
 sky130_fd_sc_hd__ha_1 _43601_ (.A(_03098_),
    .B(_03099_),
    .COUT(_03100_),
    .SUM(_03101_));
 sky130_fd_sc_hd__ha_1 _43602_ (.A(_03102_),
    .B(_03103_),
    .COUT(_03104_),
    .SUM(_22515_));
 sky130_fd_sc_hd__ha_1 _43603_ (.A(_03105_),
    .B(_03106_),
    .COUT(_03107_),
    .SUM(_03108_));
 sky130_fd_sc_hd__ha_1 _43604_ (.A(_03109_),
    .B(_03110_),
    .COUT(_03111_),
    .SUM(_22516_));
 sky130_fd_sc_hd__ha_1 _43605_ (.A(\inst$top.soc.cpu.sink__payload$12[2] ),
    .B(\inst$top.soc.cpu.sink__payload$12[3] ),
    .COUT(_03112_),
    .SUM(_03113_));
 sky130_fd_sc_hd__ha_1 _43606_ (.A(_03114_),
    .B(_03115_),
    .COUT(_03116_),
    .SUM(_03117_));
 sky130_fd_sc_hd__ha_1 _43607_ (.A(_03118_),
    .B(_03119_),
    .COUT(_03120_),
    .SUM(_22517_));
 sky130_fd_sc_hd__ha_1 _43608_ (.A(_03121_),
    .B(_03122_),
    .COUT(_03123_),
    .SUM(_03124_));
 sky130_fd_sc_hd__ha_1 _43609_ (.A(_03125_),
    .B(_03126_),
    .COUT(_03127_),
    .SUM(_22518_));
 sky130_fd_sc_hd__ha_1 _43610_ (.A(_03128_),
    .B(_03129_),
    .COUT(_03130_),
    .SUM(_03131_));
 sky130_fd_sc_hd__ha_1 _43611_ (.A(_03132_),
    .B(_03133_),
    .COUT(_03134_),
    .SUM(_22519_));
 sky130_fd_sc_hd__ha_1 _43612_ (.A(_03135_),
    .B(_03136_),
    .COUT(_03137_),
    .SUM(_03138_));
 sky130_fd_sc_hd__ha_1 _43613_ (.A(_03139_),
    .B(_03140_),
    .COUT(_03141_),
    .SUM(_22520_));
 sky130_fd_sc_hd__ha_1 _43614_ (.A(_03142_),
    .B(_03143_),
    .COUT(_03144_),
    .SUM(_03145_));
 sky130_fd_sc_hd__ha_1 _43615_ (.A(_03146_),
    .B(_03147_),
    .COUT(_03148_),
    .SUM(_22521_));
 sky130_fd_sc_hd__ha_1 _43616_ (.A(_03149_),
    .B(_03150_),
    .COUT(_03151_),
    .SUM(_03152_));
 sky130_fd_sc_hd__ha_1 _43617_ (.A(_03153_),
    .B(_03154_),
    .COUT(_03155_),
    .SUM(_22522_));
 sky130_fd_sc_hd__ha_1 _43618_ (.A(_03156_),
    .B(_03157_),
    .COUT(_03158_),
    .SUM(_03159_));
 sky130_fd_sc_hd__ha_1 _43619_ (.A(_03160_),
    .B(_03161_),
    .COUT(_03162_),
    .SUM(_22523_));
 sky130_fd_sc_hd__ha_1 _43620_ (.A(_03163_),
    .B(_03164_),
    .COUT(_03165_),
    .SUM(_03166_));
 sky130_fd_sc_hd__ha_1 _43621_ (.A(_03167_),
    .B(_03168_),
    .COUT(_03169_),
    .SUM(_22524_));
 sky130_fd_sc_hd__ha_1 _43622_ (.A(_03170_),
    .B(_03171_),
    .COUT(_03172_),
    .SUM(_03173_));
 sky130_fd_sc_hd__ha_1 _43623_ (.A(_03174_),
    .B(_03175_),
    .COUT(_03176_),
    .SUM(_22525_));
 sky130_fd_sc_hd__ha_1 _43624_ (.A(_03177_),
    .B(_03178_),
    .COUT(_03179_),
    .SUM(_03180_));
 sky130_fd_sc_hd__ha_1 _43625_ (.A(_03181_),
    .B(_03182_),
    .COUT(_03183_),
    .SUM(_22526_));
 sky130_fd_sc_hd__ha_1 _43626_ (.A(_03184_),
    .B(_03185_),
    .COUT(_03186_),
    .SUM(_03187_));
 sky130_fd_sc_hd__ha_1 _43627_ (.A(_03188_),
    .B(_03189_),
    .COUT(_03190_),
    .SUM(_22527_));
 sky130_fd_sc_hd__ha_1 _43628_ (.A(_03191_),
    .B(_03192_),
    .COUT(_03193_),
    .SUM(_03194_));
 sky130_fd_sc_hd__ha_1 _43629_ (.A(_03195_),
    .B(_03196_),
    .COUT(_03197_),
    .SUM(_22528_));
 sky130_fd_sc_hd__ha_1 _43630_ (.A(_03198_),
    .B(_03199_),
    .COUT(_03200_),
    .SUM(_03201_));
 sky130_fd_sc_hd__ha_1 _43631_ (.A(_03202_),
    .B(_03203_),
    .COUT(_03204_),
    .SUM(_22529_));
 sky130_fd_sc_hd__ha_1 _43632_ (.A(_03205_),
    .B(_03206_),
    .COUT(_03207_),
    .SUM(_03208_));
 sky130_fd_sc_hd__ha_1 _43633_ (.A(_03209_),
    .B(_03210_),
    .COUT(_03211_),
    .SUM(_22530_));
 sky130_fd_sc_hd__ha_1 _43634_ (.A(_03212_),
    .B(_03213_),
    .COUT(_03214_),
    .SUM(_03215_));
 sky130_fd_sc_hd__ha_1 _43635_ (.A(_03216_),
    .B(_03217_),
    .COUT(_03218_),
    .SUM(_22531_));
 sky130_fd_sc_hd__ha_1 _43636_ (.A(_03219_),
    .B(_03220_),
    .COUT(_03221_),
    .SUM(_03222_));
 sky130_fd_sc_hd__ha_1 _43637_ (.A(_03223_),
    .B(_03224_),
    .COUT(_03225_),
    .SUM(_22532_));
 sky130_fd_sc_hd__ha_1 _43638_ (.A(_03226_),
    .B(_03227_),
    .COUT(_03228_),
    .SUM(_03229_));
 sky130_fd_sc_hd__ha_1 _43639_ (.A(_03230_),
    .B(_03231_),
    .COUT(_03232_),
    .SUM(_22533_));
 sky130_fd_sc_hd__ha_1 _43640_ (.A(_03233_),
    .B(_03234_),
    .COUT(_03235_),
    .SUM(_03236_));
 sky130_fd_sc_hd__ha_1 _43641_ (.A(_03237_),
    .B(_03238_),
    .COUT(_03239_),
    .SUM(_22534_));
 sky130_fd_sc_hd__ha_1 _43642_ (.A(_03240_),
    .B(_03241_),
    .COUT(_03242_),
    .SUM(_03243_));
 sky130_fd_sc_hd__ha_1 _43643_ (.A(_03244_),
    .B(_03245_),
    .COUT(_03246_),
    .SUM(_22535_));
 sky130_fd_sc_hd__ha_1 _43644_ (.A(_03247_),
    .B(_03248_),
    .COUT(_03249_),
    .SUM(_03250_));
 sky130_fd_sc_hd__ha_1 _43645_ (.A(_03251_),
    .B(_03252_),
    .COUT(_03253_),
    .SUM(_22536_));
 sky130_fd_sc_hd__ha_1 _43646_ (.A(_03254_),
    .B(_03255_),
    .COUT(_03256_),
    .SUM(_03257_));
 sky130_fd_sc_hd__ha_1 _43647_ (.A(_03258_),
    .B(_03259_),
    .COUT(_03260_),
    .SUM(_22537_));
 sky130_fd_sc_hd__ha_1 _43648_ (.A(_03261_),
    .B(_03262_),
    .COUT(_03263_),
    .SUM(_03264_));
 sky130_fd_sc_hd__ha_1 _43649_ (.A(_03265_),
    .B(_03266_),
    .COUT(_03267_),
    .SUM(_22538_));
 sky130_fd_sc_hd__ha_1 _43650_ (.A(_03268_),
    .B(_03269_),
    .COUT(_03270_),
    .SUM(_03271_));
 sky130_fd_sc_hd__ha_1 _43651_ (.A(_03272_),
    .B(_03273_),
    .COUT(_03274_),
    .SUM(_22539_));
 sky130_fd_sc_hd__ha_1 _43652_ (.A(_03275_),
    .B(_03276_),
    .COUT(_03277_),
    .SUM(_03278_));
 sky130_fd_sc_hd__ha_1 _43653_ (.A(_03279_),
    .B(_03280_),
    .COUT(_03281_),
    .SUM(_22540_));
 sky130_fd_sc_hd__ha_1 _43654_ (.A(_03282_),
    .B(_03283_),
    .COUT(_03284_),
    .SUM(_03285_));
 sky130_fd_sc_hd__ha_1 _43655_ (.A(_03286_),
    .B(_03287_),
    .COUT(_03288_),
    .SUM(_22541_));
 sky130_fd_sc_hd__ha_1 _43656_ (.A(_03289_),
    .B(_03290_),
    .COUT(_03291_),
    .SUM(_03292_));
 sky130_fd_sc_hd__ha_1 _43657_ (.A(_03293_),
    .B(_03294_),
    .COUT(_03295_),
    .SUM(_22542_));
 sky130_fd_sc_hd__ha_1 _43658_ (.A(_03296_),
    .B(_03297_),
    .COUT(_03298_),
    .SUM(_03299_));
 sky130_fd_sc_hd__ha_1 _43659_ (.A(_03300_),
    .B(_03301_),
    .COUT(_03302_),
    .SUM(_22543_));
 sky130_fd_sc_hd__ha_1 _43660_ (.A(_03303_),
    .B(_03304_),
    .COUT(_03305_),
    .SUM(_03306_));
 sky130_fd_sc_hd__ha_1 _43661_ (.A(_03307_),
    .B(_03308_),
    .COUT(_03309_),
    .SUM(_22544_));
 sky130_fd_sc_hd__ha_1 _43662_ (.A(net884),
    .B(\inst$top.soc.cpu.sink__payload$6[3] ),
    .COUT(_03310_),
    .SUM(_02911_));
 sky130_fd_sc_hd__ha_1 _43663_ (.A(\inst$top.soc.cpu.csrf.d_addr[4] ),
    .B(\inst$top.soc.cpu.sink__payload$6[4] ),
    .COUT(_03311_),
    .SUM(_03312_));
 sky130_fd_sc_hd__ha_1 _43664_ (.A(\inst$top.soc.cpu.csrf.d_addr[5] ),
    .B(\inst$top.soc.cpu.sink__payload$6[5] ),
    .COUT(_03313_),
    .SUM(_03314_));
 sky130_fd_sc_hd__ha_1 _43665_ (.A(\inst$top.soc.cpu.csrf.d_addr[6] ),
    .B(\inst$top.soc.cpu.sink__payload$6[6] ),
    .COUT(_03315_),
    .SUM(_03316_));
 sky130_fd_sc_hd__ha_1 _43666_ (.A(\inst$top.soc.cpu.csrf.d_addr[7] ),
    .B(\inst$top.soc.cpu.sink__payload$6[7] ),
    .COUT(_03317_),
    .SUM(_03318_));
 sky130_fd_sc_hd__ha_1 _43667_ (.A(\inst$top.soc.cpu.csrf.d_addr[8] ),
    .B(\inst$top.soc.cpu.sink__payload$6[8] ),
    .COUT(_03319_),
    .SUM(_03320_));
 sky130_fd_sc_hd__ha_1 _43668_ (.A(\inst$top.soc.cpu.csrf.d_addr[9] ),
    .B(\inst$top.soc.cpu.sink__payload$6[9] ),
    .COUT(_03321_),
    .SUM(_03322_));
 sky130_fd_sc_hd__ha_1 _43669_ (.A(\inst$top.soc.cpu.csrf.d_addr[10] ),
    .B(\inst$top.soc.cpu.sink__payload$6[10] ),
    .COUT(_03323_),
    .SUM(_03324_));
 sky130_fd_sc_hd__ha_1 _43670_ (.A(\inst$top.soc.cpu.csrf.d_addr[11] ),
    .B(\inst$top.soc.cpu.sink__payload$6[11] ),
    .COUT(_03325_),
    .SUM(_03326_));
 sky130_fd_sc_hd__ha_1 _43671_ (.A(\inst$top.soc.cpu.d_offset[12] ),
    .B(\inst$top.soc.cpu.sink__payload$6[12] ),
    .COUT(_03327_),
    .SUM(_03328_));
 sky130_fd_sc_hd__ha_1 _43672_ (.A(\inst$top.soc.cpu.d_offset[13] ),
    .B(\inst$top.soc.cpu.sink__payload$6[13] ),
    .COUT(_03329_),
    .SUM(_03330_));
 sky130_fd_sc_hd__ha_1 _43673_ (.A(\inst$top.soc.cpu.d_offset[14] ),
    .B(\inst$top.soc.cpu.sink__payload$6[14] ),
    .COUT(_03331_),
    .SUM(_03332_));
 sky130_fd_sc_hd__ha_1 _43674_ (.A(\inst$top.soc.cpu.d_offset[15] ),
    .B(\inst$top.soc.cpu.sink__payload$6[15] ),
    .COUT(_03333_),
    .SUM(_03334_));
 sky130_fd_sc_hd__ha_1 _43675_ (.A(\inst$top.soc.cpu.d_offset[16] ),
    .B(\inst$top.soc.cpu.sink__payload$6[16] ),
    .COUT(_03335_),
    .SUM(_03336_));
 sky130_fd_sc_hd__ha_1 _43676_ (.A(\inst$top.soc.cpu.d_offset[17] ),
    .B(\inst$top.soc.cpu.sink__payload$6[17] ),
    .COUT(_03337_),
    .SUM(_03338_));
 sky130_fd_sc_hd__ha_1 _43677_ (.A(\inst$top.soc.cpu.d_offset[18] ),
    .B(\inst$top.soc.cpu.sink__payload$6[18] ),
    .COUT(_03339_),
    .SUM(_03340_));
 sky130_fd_sc_hd__ha_1 _43678_ (.A(\inst$top.soc.cpu.d_offset[19] ),
    .B(\inst$top.soc.cpu.sink__payload$6[19] ),
    .COUT(_03341_),
    .SUM(_03342_));
 sky130_fd_sc_hd__ha_1 _43679_ (.A(\inst$top.soc.cpu.d_offset[20] ),
    .B(\inst$top.soc.cpu.sink__payload$6[20] ),
    .COUT(_03343_),
    .SUM(_03344_));
 sky130_fd_sc_hd__ha_1 _43680_ (.A(\inst$top.soc.cpu.d_offset[21] ),
    .B(\inst$top.soc.cpu.sink__payload$6[21] ),
    .COUT(_03345_),
    .SUM(_03346_));
 sky130_fd_sc_hd__ha_1 _43681_ (.A(\inst$top.soc.cpu.d_offset[22] ),
    .B(\inst$top.soc.cpu.sink__payload$6[22] ),
    .COUT(_03347_),
    .SUM(_03348_));
 sky130_fd_sc_hd__ha_1 _43682_ (.A(\inst$top.soc.cpu.d_offset[23] ),
    .B(\inst$top.soc.cpu.sink__payload$6[23] ),
    .COUT(_03349_),
    .SUM(_03350_));
 sky130_fd_sc_hd__ha_1 _43683_ (.A(\inst$top.soc.cpu.d_offset[24] ),
    .B(\inst$top.soc.cpu.sink__payload$6[24] ),
    .COUT(_03351_),
    .SUM(_03352_));
 sky130_fd_sc_hd__ha_1 _43684_ (.A(\inst$top.soc.cpu.d_offset[25] ),
    .B(\inst$top.soc.cpu.sink__payload$6[25] ),
    .COUT(_03353_),
    .SUM(_03354_));
 sky130_fd_sc_hd__ha_1 _43685_ (.A(\inst$top.soc.cpu.d_offset[26] ),
    .B(\inst$top.soc.cpu.sink__payload$6[26] ),
    .COUT(_03355_),
    .SUM(_03356_));
 sky130_fd_sc_hd__ha_1 _43686_ (.A(\inst$top.soc.cpu.d_offset[27] ),
    .B(\inst$top.soc.cpu.sink__payload$6[27] ),
    .COUT(_03357_),
    .SUM(_03358_));
 sky130_fd_sc_hd__ha_1 _43687_ (.A(\inst$top.soc.cpu.d_offset[28] ),
    .B(\inst$top.soc.cpu.sink__payload$6[28] ),
    .COUT(_03359_),
    .SUM(_03360_));
 sky130_fd_sc_hd__ha_1 _43688_ (.A(\inst$top.soc.cpu.d_offset[29] ),
    .B(\inst$top.soc.cpu.sink__payload$6[29] ),
    .COUT(_03361_),
    .SUM(_03362_));
 sky130_fd_sc_hd__ha_1 _43689_ (.A(\inst$top.soc.cpu.d_offset[30] ),
    .B(\inst$top.soc.cpu.sink__payload$6[30] ),
    .COUT(_03363_),
    .SUM(_03364_));
 sky130_fd_sc_hd__ha_1 _43690_ (.A(_03366_),
    .B(_03367_),
    .COUT(_22545_),
    .SUM(_22546_));
 sky130_fd_sc_hd__ha_1 _43691_ (.A(_03368_),
    .B(_03369_),
    .COUT(_03365_),
    .SUM(_22547_));
 sky130_fd_sc_hd__ha_1 _43692_ (.A(_03371_),
    .B(_22546_),
    .COUT(_22548_),
    .SUM(_22549_));
 sky130_fd_sc_hd__ha_1 _43693_ (.A(_22547_),
    .B(_03372_),
    .COUT(_03370_),
    .SUM(_03373_));
 sky130_fd_sc_hd__ha_1 _43694_ (.A(_22550_),
    .B(_22549_),
    .COUT(_22551_),
    .SUM(_22462_));
 sky130_fd_sc_hd__ha_1 _43695_ (.A(_03375_),
    .B(_03376_),
    .COUT(_22550_),
    .SUM(_22552_));
 sky130_fd_sc_hd__ha_1 _43696_ (.A(_03377_),
    .B(_03378_),
    .COUT(_03374_),
    .SUM(_22553_));
 sky130_fd_sc_hd__ha_1 _43697_ (.A(_22461_),
    .B(_22462_),
    .COUT(_03379_),
    .SUM(_02915_));
 sky130_fd_sc_hd__ha_1 _43698_ (.A(_22554_),
    .B(_22552_),
    .COUT(_22461_),
    .SUM(_22480_));
 sky130_fd_sc_hd__ha_1 _43699_ (.A(_03380_),
    .B(_22555_),
    .COUT(_22554_),
    .SUM(_22478_));
 sky130_fd_sc_hd__ha_1 _43700_ (.A(_22553_),
    .B(_03381_),
    .COUT(_22555_),
    .SUM(_22476_));
 sky130_fd_sc_hd__ha_1 _43701_ (.A(_03382_),
    .B(_03383_),
    .COUT(_22556_),
    .SUM(_22557_));
 sky130_fd_sc_hd__ha_1 _43702_ (.A(_03384_),
    .B(_22557_),
    .COUT(_22558_),
    .SUM(_22559_));
 sky130_fd_sc_hd__ha_1 _43703_ (.A(_22545_),
    .B(_22559_),
    .COUT(_22560_),
    .SUM(_22561_));
 sky130_fd_sc_hd__ha_1 _43704_ (.A(_03385_),
    .B(_22561_),
    .COUT(_22562_),
    .SUM(_22563_));
 sky130_fd_sc_hd__ha_1 _43705_ (.A(_22548_),
    .B(_22563_),
    .COUT(_22564_),
    .SUM(_22565_));
 sky130_fd_sc_hd__ha_1 _43706_ (.A(_22551_),
    .B(_22565_),
    .COUT(_03386_),
    .SUM(_03387_));
 sky130_fd_sc_hd__ha_1 _43707_ (.A(_22556_),
    .B(_20840_),
    .COUT(_22566_),
    .SUM(_22567_));
 sky130_fd_sc_hd__ha_1 _43708_ (.A(_03388_),
    .B(_22567_),
    .COUT(_22568_),
    .SUM(_22569_));
 sky130_fd_sc_hd__ha_1 _43709_ (.A(_22558_),
    .B(_22569_),
    .COUT(_22570_),
    .SUM(_22571_));
 sky130_fd_sc_hd__ha_1 _43710_ (.A(_03389_),
    .B(_22560_),
    .COUT(_03390_),
    .SUM(_22572_));
 sky130_fd_sc_hd__ha_1 _43711_ (.A(_22572_),
    .B(_22571_),
    .COUT(_03391_),
    .SUM(_22573_));
 sky130_fd_sc_hd__ha_1 _43712_ (.A(_22562_),
    .B(_22573_),
    .COUT(_22574_),
    .SUM(_22575_));
 sky130_fd_sc_hd__ha_1 _43713_ (.A(_22564_),
    .B(_22575_),
    .COUT(_03392_),
    .SUM(_03393_));
 sky130_fd_sc_hd__ha_1 _43714_ (.A(_20839_),
    .B(_20844_),
    .COUT(_22576_),
    .SUM(_22577_));
 sky130_fd_sc_hd__ha_1 _43715_ (.A(_22566_),
    .B(_22577_),
    .COUT(_20851_),
    .SUM(_22578_));
 sky130_fd_sc_hd__ha_1 _43716_ (.A(_03394_),
    .B(_22578_),
    .COUT(_22579_),
    .SUM(_22580_));
 sky130_fd_sc_hd__ha_1 _43717_ (.A(_22568_),
    .B(_22580_),
    .COUT(_22581_),
    .SUM(_22582_));
 sky130_fd_sc_hd__ha_1 _43718_ (.A(_22582_),
    .B(_03395_),
    .COUT(_20856_),
    .SUM(_22583_));
 sky130_fd_sc_hd__ha_1 _43719_ (.A(_03396_),
    .B(_22570_),
    .COUT(_03397_),
    .SUM(_22584_));
 sky130_fd_sc_hd__ha_1 _43720_ (.A(_22584_),
    .B(_22583_),
    .COUT(_03398_),
    .SUM(_03399_));
 sky130_fd_sc_hd__ha_1 _43721_ (.A(_22574_),
    .B(_03400_),
    .COUT(_03401_),
    .SUM(_03402_));
 sky130_fd_sc_hd__ha_1 _43722_ (.A(_03403_),
    .B(_03404_),
    .COUT(_20861_),
    .SUM(_22585_));
 sky130_fd_sc_hd__ha_1 _43723_ (.A(_20843_),
    .B(_20848_),
    .COUT(_22586_),
    .SUM(_22587_));
 sky130_fd_sc_hd__ha_1 _43724_ (.A(_22576_),
    .B(_22587_),
    .COUT(_20866_),
    .SUM(_20852_));
 sky130_fd_sc_hd__ha_1 _43725_ (.A(_22579_),
    .B(_20854_),
    .COUT(_22588_),
    .SUM(_22589_));
 sky130_fd_sc_hd__ha_1 _43726_ (.A(_22589_),
    .B(_22585_),
    .COUT(_20871_),
    .SUM(_20857_));
 sky130_fd_sc_hd__ha_1 _43727_ (.A(_03405_),
    .B(_22581_),
    .COUT(_20875_),
    .SUM(_20855_));
 sky130_fd_sc_hd__ha_1 _43728_ (.A(_03406_),
    .B(_03407_),
    .COUT(_03408_),
    .SUM(_03409_));
 sky130_fd_sc_hd__ha_1 _43729_ (.A(_22586_),
    .B(_20863_),
    .COUT(_20883_),
    .SUM(_20867_));
 sky130_fd_sc_hd__ha_1 _43730_ (.A(_20853_),
    .B(_20869_),
    .COUT(_22590_),
    .SUM(_22591_));
 sky130_fd_sc_hd__ha_1 _43731_ (.A(_22591_),
    .B(_03410_),
    .COUT(_20888_),
    .SUM(_20872_));
 sky130_fd_sc_hd__ha_1 _43732_ (.A(_03411_),
    .B(_22588_),
    .COUT(_20892_),
    .SUM(_20870_));
 sky130_fd_sc_hd__ha_1 _43733_ (.A(_03412_),
    .B(_20877_),
    .COUT(_03413_),
    .SUM(_03414_));
 sky130_fd_sc_hd__ha_1 _43734_ (.A(_03415_),
    .B(_03416_),
    .COUT(_20896_),
    .SUM(_22592_));
 sky130_fd_sc_hd__ha_1 _43735_ (.A(_20862_),
    .B(_03417_),
    .COUT(_20900_),
    .SUM(_20884_));
 sky130_fd_sc_hd__ha_1 _43736_ (.A(_20868_),
    .B(_20886_),
    .COUT(_22593_),
    .SUM(_22594_));
 sky130_fd_sc_hd__ha_1 _43737_ (.A(_22594_),
    .B(_22592_),
    .COUT(_20904_),
    .SUM(_20889_));
 sky130_fd_sc_hd__ha_1 _43738_ (.A(_03418_),
    .B(_22590_),
    .COUT(_20908_),
    .SUM(_20887_));
 sky130_fd_sc_hd__ha_1 _43739_ (.A(_20876_),
    .B(_20894_),
    .COUT(_03419_),
    .SUM(_03420_));
 sky130_fd_sc_hd__ha_1 _43740_ (.A(_03421_),
    .B(_03422_),
    .COUT(_03423_),
    .SUM(_22595_));
 sky130_fd_sc_hd__ha_1 _43741_ (.A(_03424_),
    .B(_22595_),
    .COUT(_20915_),
    .SUM(_22596_));
 sky130_fd_sc_hd__ha_1 _43742_ (.A(_20885_),
    .B(_20902_),
    .COUT(_22597_),
    .SUM(_22598_));
 sky130_fd_sc_hd__ha_1 _43743_ (.A(_22598_),
    .B(_22596_),
    .COUT(_20920_),
    .SUM(_20905_));
 sky130_fd_sc_hd__ha_1 _43744_ (.A(_03425_),
    .B(_22593_),
    .COUT(_20924_),
    .SUM(_20903_));
 sky130_fd_sc_hd__ha_1 _43745_ (.A(_20893_),
    .B(_20910_),
    .COUT(_03426_),
    .SUM(_03427_));
 sky130_fd_sc_hd__ha_1 _43746_ (.A(_20901_),
    .B(_03428_),
    .COUT(_22599_),
    .SUM(_22600_));
 sky130_fd_sc_hd__ha_1 _43747_ (.A(_22600_),
    .B(_03429_),
    .COUT(_03430_),
    .SUM(_20921_));
 sky130_fd_sc_hd__ha_1 _43748_ (.A(_03431_),
    .B(_22597_),
    .COUT(_20942_),
    .SUM(_20919_));
 sky130_fd_sc_hd__ha_1 _43749_ (.A(_20909_),
    .B(_20926_),
    .COUT(_03432_),
    .SUM(_03433_));
 sky130_fd_sc_hd__ha_1 _43750_ (.A(_03434_),
    .B(_03435_),
    .COUT(_22601_),
    .SUM(_22602_));
 sky130_fd_sc_hd__ha_1 _43751_ (.A(_03436_),
    .B(_03437_),
    .COUT(_22603_),
    .SUM(_22604_));
 sky130_fd_sc_hd__ha_1 _43752_ (.A(_22604_),
    .B(_22602_),
    .COUT(_03438_),
    .SUM(_03439_));
 sky130_fd_sc_hd__ha_1 _43753_ (.A(_03440_),
    .B(_22599_),
    .COUT(_00485_),
    .SUM(_03441_));
 sky130_fd_sc_hd__ha_1 _43754_ (.A(_20925_),
    .B(_20944_),
    .COUT(_03442_),
    .SUM(_03443_));
 sky130_fd_sc_hd__ha_1 _43755_ (.A(_03444_),
    .B(_03445_),
    .COUT(_22605_),
    .SUM(_22606_));
 sky130_fd_sc_hd__ha_1 _43756_ (.A(_03446_),
    .B(_22606_),
    .COUT(_22607_),
    .SUM(_22608_));
 sky130_fd_sc_hd__ha_1 _43757_ (.A(_22601_),
    .B(_22608_),
    .COUT(_03447_),
    .SUM(_22609_));
 sky130_fd_sc_hd__ha_1 _43758_ (.A(_03448_),
    .B(_03449_),
    .COUT(_22610_),
    .SUM(_22611_));
 sky130_fd_sc_hd__ha_1 _43759_ (.A(_22611_),
    .B(_22609_),
    .COUT(_20983_),
    .SUM(_03450_));
 sky130_fd_sc_hd__ha_1 _43760_ (.A(_03451_),
    .B(_22603_),
    .COUT(_00522_),
    .SUM(_03452_));
 sky130_fd_sc_hd__ha_1 _43761_ (.A(_20943_),
    .B(_03453_),
    .COUT(_03454_),
    .SUM(_03455_));
 sky130_fd_sc_hd__ha_1 _43762_ (.A(_22605_),
    .B(_20965_),
    .COUT(_20990_),
    .SUM(_22612_));
 sky130_fd_sc_hd__ha_1 _43763_ (.A(_03456_),
    .B(_22612_),
    .COUT(_22613_),
    .SUM(_22614_));
 sky130_fd_sc_hd__ha_1 _43764_ (.A(_22607_),
    .B(_22614_),
    .COUT(_03457_),
    .SUM(_22615_));
 sky130_fd_sc_hd__ha_1 _43765_ (.A(_03458_),
    .B(_22615_),
    .COUT(_03459_),
    .SUM(_20984_));
 sky130_fd_sc_hd__ha_1 _43766_ (.A(_03460_),
    .B(_22610_),
    .COUT(_00565_),
    .SUM(_20982_));
 sky130_fd_sc_hd__ha_1 _43767_ (.A(_03461_),
    .B(_03462_),
    .COUT(_03463_),
    .SUM(_03464_));
 sky130_fd_sc_hd__ha_1 _43768_ (.A(_20964_),
    .B(_20986_),
    .COUT(_21012_),
    .SUM(_20991_));
 sky130_fd_sc_hd__ha_1 _43769_ (.A(_22613_),
    .B(_20993_),
    .COUT(_03465_),
    .SUM(_22616_));
 sky130_fd_sc_hd__ha_1 _43770_ (.A(_22616_),
    .B(_03466_),
    .COUT(_21027_),
    .SUM(_22617_));
 sky130_fd_sc_hd__ha_1 _43771_ (.A(_03467_),
    .B(_22617_),
    .COUT(_03468_),
    .SUM(_03469_));
 sky130_fd_sc_hd__ha_1 _43772_ (.A(_03470_),
    .B(_03471_),
    .COUT(_00610_),
    .SUM(_03472_));
 sky130_fd_sc_hd__ha_1 _43773_ (.A(_03473_),
    .B(_03474_),
    .COUT(_03475_),
    .SUM(_03476_));
 sky130_fd_sc_hd__ha_1 _43774_ (.A(_03477_),
    .B(_03478_),
    .COUT(_21033_),
    .SUM(_22618_));
 sky130_fd_sc_hd__ha_1 _43775_ (.A(_20985_),
    .B(_03479_),
    .COUT(_21040_),
    .SUM(_21013_));
 sky130_fd_sc_hd__ha_1 _43776_ (.A(_20992_),
    .B(_21015_),
    .COUT(_03480_),
    .SUM(_22619_));
 sky130_fd_sc_hd__ha_1 _43777_ (.A(_22619_),
    .B(_22618_),
    .COUT(_21054_),
    .SUM(_21028_));
 sky130_fd_sc_hd__ha_1 _43778_ (.A(_03481_),
    .B(_03482_),
    .COUT(_00660_),
    .SUM(_03483_));
 sky130_fd_sc_hd__ha_1 _43779_ (.A(_03484_),
    .B(_03485_),
    .COUT(_03486_),
    .SUM(_03487_));
 sky130_fd_sc_hd__ha_1 _43780_ (.A(_21014_),
    .B(_21042_),
    .COUT(_03488_),
    .SUM(_22620_));
 sky130_fd_sc_hd__ha_1 _43781_ (.A(_22620_),
    .B(_03489_),
    .COUT(_21079_),
    .SUM(_21055_));
 sky130_fd_sc_hd__ha_1 _43782_ (.A(_03490_),
    .B(_03491_),
    .COUT(_00708_),
    .SUM(_03492_));
 sky130_fd_sc_hd__ha_1 _43783_ (.A(_03493_),
    .B(_03494_),
    .COUT(_03495_),
    .SUM(_03496_));
 sky130_fd_sc_hd__ha_1 _43784_ (.A(_03497_),
    .B(_03498_),
    .COUT(_22621_),
    .SUM(_22622_));
 sky130_fd_sc_hd__ha_1 _43785_ (.A(_21041_),
    .B(_03499_),
    .COUT(_03500_),
    .SUM(_22623_));
 sky130_fd_sc_hd__ha_1 _43786_ (.A(_22623_),
    .B(_22622_),
    .COUT(_03501_),
    .SUM(_21080_));
 sky130_fd_sc_hd__ha_1 _43787_ (.A(_03502_),
    .B(_03503_),
    .COUT(_00756_),
    .SUM(_03504_));
 sky130_fd_sc_hd__ha_1 _43788_ (.A(_03505_),
    .B(_03506_),
    .COUT(_03507_),
    .SUM(_03508_));
 sky130_fd_sc_hd__ha_1 _43789_ (.A(_03509_),
    .B(_03510_),
    .COUT(_03511_),
    .SUM(_22624_));
 sky130_fd_sc_hd__ha_1 _43790_ (.A(_03512_),
    .B(_22624_),
    .COUT(_22625_),
    .SUM(_22626_));
 sky130_fd_sc_hd__ha_1 _43791_ (.A(_22621_),
    .B(_22626_),
    .COUT(_03513_),
    .SUM(_22627_));
 sky130_fd_sc_hd__ha_1 _43792_ (.A(_03514_),
    .B(_21092_),
    .COUT(_21131_),
    .SUM(_22628_));
 sky130_fd_sc_hd__ha_1 _43793_ (.A(_22628_),
    .B(_22627_),
    .COUT(_21134_),
    .SUM(_03515_));
 sky130_fd_sc_hd__ha_1 _43794_ (.A(_03516_),
    .B(_03517_),
    .COUT(_00811_),
    .SUM(_03518_));
 sky130_fd_sc_hd__ha_1 _43795_ (.A(_03519_),
    .B(_03520_),
    .COUT(_03521_),
    .SUM(_03522_));
 sky130_fd_sc_hd__ha_1 _43796_ (.A(_22625_),
    .B(_03523_),
    .COUT(_03524_),
    .SUM(_22629_));
 sky130_fd_sc_hd__ha_1 _43797_ (.A(_03525_),
    .B(_22629_),
    .COUT(_03526_),
    .SUM(_21135_));
 sky130_fd_sc_hd__ha_1 _43798_ (.A(_03527_),
    .B(_03528_),
    .COUT(_00868_),
    .SUM(_03529_));
 sky130_fd_sc_hd__ha_1 _43799_ (.A(_03530_),
    .B(_03531_),
    .COUT(_03532_),
    .SUM(_03533_));
 sky130_fd_sc_hd__ha_1 _43800_ (.A(_03534_),
    .B(_03535_),
    .COUT(_03536_),
    .SUM(_22630_));
 sky130_fd_sc_hd__ha_1 _43801_ (.A(_22630_),
    .B(_03537_),
    .COUT(_21182_),
    .SUM(_22631_));
 sky130_fd_sc_hd__ha_1 _43802_ (.A(_03538_),
    .B(_22631_),
    .COUT(_03539_),
    .SUM(_03540_));
 sky130_fd_sc_hd__ha_1 _43803_ (.A(_03541_),
    .B(_21132_),
    .COUT(_00924_),
    .SUM(_03542_));
 sky130_fd_sc_hd__ha_1 _43804_ (.A(_03543_),
    .B(_03544_),
    .COUT(_03545_),
    .SUM(_03546_));
 sky130_fd_sc_hd__ha_1 _43805_ (.A(_03547_),
    .B(_03548_),
    .COUT(_22632_),
    .SUM(_22633_));
 sky130_fd_sc_hd__ha_1 _43806_ (.A(_03549_),
    .B(_03550_),
    .COUT(_03551_),
    .SUM(_22634_));
 sky130_fd_sc_hd__ha_1 _43807_ (.A(_22634_),
    .B(_22633_),
    .COUT(_03552_),
    .SUM(_21183_));
 sky130_fd_sc_hd__ha_1 _43808_ (.A(_03553_),
    .B(_21161_),
    .COUT(_00978_),
    .SUM(_03554_));
 sky130_fd_sc_hd__ha_1 _43809_ (.A(_03555_),
    .B(_03556_),
    .COUT(_03557_),
    .SUM(_03558_));
 sky130_fd_sc_hd__ha_1 _43810_ (.A(_22632_),
    .B(_21199_),
    .COUT(_03559_),
    .SUM(_22635_));
 sky130_fd_sc_hd__ha_1 _43811_ (.A(_03560_),
    .B(_03561_),
    .COUT(_03562_),
    .SUM(_22636_));
 sky130_fd_sc_hd__ha_1 _43812_ (.A(_22636_),
    .B(_22635_),
    .COUT(_03563_),
    .SUM(_03564_));
 sky130_fd_sc_hd__ha_1 _43813_ (.A(_03565_),
    .B(_21193_),
    .COUT(_01037_),
    .SUM(_03566_));
 sky130_fd_sc_hd__ha_1 _43814_ (.A(_03567_),
    .B(_03568_),
    .COUT(_03569_),
    .SUM(_03570_));
 sky130_fd_sc_hd__ha_1 _43815_ (.A(_21198_),
    .B(_03571_),
    .COUT(_03572_),
    .SUM(_22637_));
 sky130_fd_sc_hd__ha_1 _43816_ (.A(_22637_),
    .B(_03573_),
    .COUT(_21276_),
    .SUM(_22638_));
 sky130_fd_sc_hd__ha_1 _43817_ (.A(_03574_),
    .B(_22638_),
    .COUT(_03575_),
    .SUM(_03576_));
 sky130_fd_sc_hd__ha_1 _43818_ (.A(_03577_),
    .B(_21229_),
    .COUT(_01098_),
    .SUM(_03578_));
 sky130_fd_sc_hd__ha_1 _43819_ (.A(_03579_),
    .B(_03580_),
    .COUT(_03581_),
    .SUM(_03582_));
 sky130_fd_sc_hd__ha_1 _43820_ (.A(_03583_),
    .B(_03584_),
    .COUT(_03585_),
    .SUM(_22639_));
 sky130_fd_sc_hd__ha_1 _43821_ (.A(_03586_),
    .B(_03587_),
    .COUT(_03588_),
    .SUM(_22640_));
 sky130_fd_sc_hd__ha_1 _43822_ (.A(_22640_),
    .B(_22639_),
    .COUT(_03589_),
    .SUM(_21277_));
 sky130_fd_sc_hd__ha_1 _43823_ (.A(_03590_),
    .B(_21263_),
    .COUT(_01164_),
    .SUM(_03591_));
 sky130_fd_sc_hd__ha_1 _43824_ (.A(_03592_),
    .B(_03593_),
    .COUT(_03594_),
    .SUM(_03595_));
 sky130_fd_sc_hd__ha_1 _43825_ (.A(_03596_),
    .B(_03597_),
    .COUT(_21355_),
    .SUM(_03598_));
 sky130_fd_sc_hd__ha_1 _43826_ (.A(_03599_),
    .B(_21300_),
    .COUT(_01226_),
    .SUM(_03600_));
 sky130_fd_sc_hd__ha_1 _43827_ (.A(_03601_),
    .B(_03602_),
    .COUT(_03603_),
    .SUM(_03604_));
 sky130_fd_sc_hd__ha_1 _43828_ (.A(_03605_),
    .B(_03606_),
    .COUT(_03607_),
    .SUM(_22641_));
 sky130_fd_sc_hd__ha_1 _43829_ (.A(_03608_),
    .B(_22641_),
    .COUT(_03609_),
    .SUM(_21356_));
 sky130_fd_sc_hd__ha_1 _43830_ (.A(_03610_),
    .B(_21339_),
    .COUT(_01285_),
    .SUM(_03611_));
 sky130_fd_sc_hd__ha_1 _43831_ (.A(_03612_),
    .B(_03613_),
    .COUT(_03614_),
    .SUM(_03615_));
 sky130_fd_sc_hd__ha_1 _43832_ (.A(_03616_),
    .B(_03617_),
    .COUT(_03618_),
    .SUM(_22642_));
 sky130_fd_sc_hd__ha_1 _43833_ (.A(_03619_),
    .B(_22642_),
    .COUT(_03620_),
    .SUM(_03621_));
 sky130_fd_sc_hd__ha_1 _43834_ (.A(_03622_),
    .B(_21381_),
    .COUT(_01350_),
    .SUM(_03623_));
 sky130_fd_sc_hd__ha_1 _43835_ (.A(_03624_),
    .B(_03625_),
    .COUT(_03626_),
    .SUM(_03627_));
 sky130_fd_sc_hd__ha_1 _43836_ (.A(_03628_),
    .B(_03629_),
    .COUT(_03630_),
    .SUM(_03631_));
 sky130_fd_sc_hd__ha_1 _43837_ (.A(_03632_),
    .B(_03633_),
    .COUT(_03634_),
    .SUM(_03635_));
 sky130_fd_sc_hd__ha_1 _43838_ (.A(_03636_),
    .B(_21471_),
    .COUT(_01468_),
    .SUM(_03637_));
 sky130_fd_sc_hd__ha_1 _43839_ (.A(_03638_),
    .B(_03639_),
    .COUT(_03640_),
    .SUM(_03641_));
 sky130_fd_sc_hd__ha_1 _43840_ (.A(_03642_),
    .B(_21520_),
    .COUT(_01524_),
    .SUM(_03643_));
 sky130_fd_sc_hd__ha_1 _43841_ (.A(_03644_),
    .B(_03645_),
    .COUT(_03646_),
    .SUM(_03647_));
 sky130_fd_sc_hd__ha_1 _43842_ (.A(_03648_),
    .B(_21569_),
    .COUT(_01582_),
    .SUM(_03649_));
 sky130_fd_sc_hd__ha_1 _43843_ (.A(_03650_),
    .B(_03651_),
    .COUT(_03652_),
    .SUM(_03653_));
 sky130_fd_sc_hd__ha_1 _43844_ (.A(_03654_),
    .B(_21616_),
    .COUT(_01636_),
    .SUM(_03655_));
 sky130_fd_sc_hd__ha_1 _43845_ (.A(_03656_),
    .B(_03657_),
    .COUT(_03658_),
    .SUM(_03659_));
 sky130_fd_sc_hd__ha_1 _43846_ (.A(_03660_),
    .B(_21661_),
    .COUT(_01688_),
    .SUM(_03661_));
 sky130_fd_sc_hd__ha_1 _43847_ (.A(_03662_),
    .B(_03663_),
    .COUT(_03664_),
    .SUM(_03665_));
 sky130_fd_sc_hd__ha_1 _43848_ (.A(_03666_),
    .B(_21710_),
    .COUT(_01738_),
    .SUM(_03667_));
 sky130_fd_sc_hd__ha_1 _43849_ (.A(_03668_),
    .B(_03669_),
    .COUT(_03670_),
    .SUM(_03671_));
 sky130_fd_sc_hd__dfxtp_1 _43850_ (.CLK(clknet_leaf_130_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[0] ),
    .Q(_00096_));
 sky130_fd_sc_hd__dfxtp_1 _43851_ (.CLK(clknet_leaf_128_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[1] ),
    .Q(_00107_));
 sky130_fd_sc_hd__dfxtp_1 _43852_ (.CLK(clknet_leaf_128_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[2] ),
    .Q(_00118_));
 sky130_fd_sc_hd__dfxtp_1 _43853_ (.CLK(clknet_leaf_129_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[3] ),
    .Q(_00121_));
 sky130_fd_sc_hd__dfxtp_1 _43854_ (.CLK(clknet_leaf_130_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[4] ),
    .Q(_00122_));
 sky130_fd_sc_hd__dfxtp_1 _43855_ (.CLK(clknet_leaf_130_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[5] ),
    .Q(_00123_));
 sky130_fd_sc_hd__dfxtp_1 _43856_ (.CLK(clknet_leaf_129_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[6] ),
    .Q(_00124_));
 sky130_fd_sc_hd__dfxtp_1 _43857_ (.CLK(clknet_leaf_127_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[7] ),
    .Q(_00125_));
 sky130_fd_sc_hd__dfxtp_1 _43858_ (.CLK(clknet_leaf_131_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[8] ),
    .Q(_00126_));
 sky130_fd_sc_hd__dfxtp_1 _43859_ (.CLK(clknet_leaf_127_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[9] ),
    .Q(_00127_));
 sky130_fd_sc_hd__dfxtp_1 _43860_ (.CLK(clknet_leaf_129_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[10] ),
    .Q(_00097_));
 sky130_fd_sc_hd__dfxtp_1 _43861_ (.CLK(clknet_leaf_131_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[11] ),
    .Q(_00098_));
 sky130_fd_sc_hd__dfxtp_1 _43862_ (.CLK(clknet_leaf_128_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[12] ),
    .Q(_00099_));
 sky130_fd_sc_hd__dfxtp_1 _43863_ (.CLK(clknet_leaf_128_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[13] ),
    .Q(_00100_));
 sky130_fd_sc_hd__dfxtp_1 _43864_ (.CLK(clknet_leaf_131_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[14] ),
    .Q(_00101_));
 sky130_fd_sc_hd__dfxtp_1 _43865_ (.CLK(clknet_leaf_129_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[15] ),
    .Q(_00102_));
 sky130_fd_sc_hd__dfxtp_1 _43866_ (.CLK(clknet_leaf_132_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[16] ),
    .Q(_00103_));
 sky130_fd_sc_hd__dfxtp_1 _43867_ (.CLK(clknet_leaf_132_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[17] ),
    .Q(_00104_));
 sky130_fd_sc_hd__dfxtp_1 _43868_ (.CLK(clknet_leaf_127_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[18] ),
    .Q(_00105_));
 sky130_fd_sc_hd__dfxtp_1 _43869_ (.CLK(clknet_leaf_132_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[19] ),
    .Q(_00106_));
 sky130_fd_sc_hd__dfxtp_1 _43870_ (.CLK(clknet_leaf_127_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[20] ),
    .Q(_00108_));
 sky130_fd_sc_hd__dfxtp_1 _43871_ (.CLK(clknet_leaf_132_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[21] ),
    .Q(_00109_));
 sky130_fd_sc_hd__dfxtp_1 _43872_ (.CLK(clknet_leaf_132_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[22] ),
    .Q(_00110_));
 sky130_fd_sc_hd__dfxtp_1 _43873_ (.CLK(clknet_6_32__leaf_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[23] ),
    .Q(_00111_));
 sky130_fd_sc_hd__dfxtp_1 _43874_ (.CLK(clknet_leaf_129_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[24] ),
    .Q(_00112_));
 sky130_fd_sc_hd__dfxtp_1 _43875_ (.CLK(clknet_leaf_128_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[25] ),
    .Q(_00113_));
 sky130_fd_sc_hd__dfxtp_1 _43876_ (.CLK(clknet_leaf_129_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[26] ),
    .Q(_00114_));
 sky130_fd_sc_hd__dfxtp_1 _43877_ (.CLK(clknet_leaf_128_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[27] ),
    .Q(_00115_));
 sky130_fd_sc_hd__dfxtp_1 _43878_ (.CLK(clknet_leaf_129_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[28] ),
    .Q(_00116_));
 sky130_fd_sc_hd__dfxtp_1 _43879_ (.CLK(clknet_leaf_131_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[29] ),
    .Q(_00117_));
 sky130_fd_sc_hd__dfxtp_1 _43880_ (.CLK(clknet_leaf_129_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[30] ),
    .Q(_00119_));
 sky130_fd_sc_hd__dfxtp_1 _43881_ (.CLK(clknet_leaf_129_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__data[31] ),
    .Q(_00120_));
 sky130_fd_sc_hd__dfxtp_1 _43882_ (.CLK(clknet_leaf_127_clk_in_regs),
    .D(\inst$top.soc.sram.read_port__en ),
    .Q(_00128_));
 sky130_fd_sc_hd__conb_1 _44017__442 (.HI(gpio_dm0[0]));
 sky130_fd_sc_hd__dfxtp_2 \inst$top.rst_n_sync.rst$_DFF_P_  (.CLK(clknet_6_17__leaf_clk_in_regs),
    .D(\inst$top.rst_n_sync.stage0 ),
    .Q(\inst$top.rst_n_sync.rst ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.rst_n_sync.stage0$_DFF_P_  (.CLK(clknet_6_5__leaf_clk_in_regs),
    .D(\inst$top.i$88 ),
    .Q(\inst$top.rst_n_sync.stage0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.a.source__valid$_SDFFE_PP0P_  (.CLK(clknet_leaf_776_clk_in_regs),
    .D(_03672_),
    .Q(\inst$top.soc.cpu.a.source__valid ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.csrf.bank_300_m_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_659_clk_in_regs),
    .D(_03673_),
    .Q(\inst$top.soc.cpu.csrf.bank_300_m_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.csrf.bank_300_w_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_716_clk_in_regs),
    .D(_03674_),
    .Q(\inst$top.soc.cpu.csrf.bank_300_w_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.csrf.bank_300_x_select$_SDFFE_PP0P_  (.CLK(clknet_leaf_593_clk_in_regs),
    .D(_03675_),
    .Q(\inst$top.soc.cpu.csrf.bank_300_x_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.d.source__valid$_SDFFE_PP0P_  (.CLK(clknet_leaf_758_clk_in_regs),
    .D(_03676_),
    .Q(\inst$top.soc.cpu.d.source__valid ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_551_clk_in_regs),
    .D(_03677_),
    .Q(\inst$top.soc.cpu.divider.divisor[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_700_clk_in_regs),
    .D(_03678_),
    .Q(\inst$top.soc.cpu.divider.divisor[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_696_clk_in_regs),
    .D(_03679_),
    .Q(\inst$top.soc.cpu.divider.divisor[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_702_clk_in_regs),
    .D(_03680_),
    .Q(\inst$top.soc.cpu.divider.divisor[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_702_clk_in_regs),
    .D(_03681_),
    .Q(\inst$top.soc.cpu.divider.divisor[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_702_clk_in_regs),
    .D(_03682_),
    .Q(\inst$top.soc.cpu.divider.divisor[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_550_clk_in_regs),
    .D(_03683_),
    .Q(\inst$top.soc.cpu.divider.divisor[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_703_clk_in_regs),
    .D(_03684_),
    .Q(\inst$top.soc.cpu.divider.divisor[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_712_clk_in_regs),
    .D(_03685_),
    .Q(\inst$top.soc.cpu.divider.divisor[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_712_clk_in_regs),
    .D(_03686_),
    .Q(\inst$top.soc.cpu.divider.divisor[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_711_clk_in_regs),
    .D(_03687_),
    .Q(\inst$top.soc.cpu.divider.divisor[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_551_clk_in_regs),
    .D(_03688_),
    .Q(\inst$top.soc.cpu.divider.divisor[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_711_clk_in_regs),
    .D(_03689_),
    .Q(\inst$top.soc.cpu.divider.divisor[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_708_clk_in_regs),
    .D(_03690_),
    .Q(\inst$top.soc.cpu.divider.divisor[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_708_clk_in_regs),
    .D(_03691_),
    .Q(\inst$top.soc.cpu.divider.divisor[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_549_clk_in_regs),
    .D(_03692_),
    .Q(\inst$top.soc.cpu.divider.divisor[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_547_clk_in_regs),
    .D(_03693_),
    .Q(\inst$top.soc.cpu.divider.divisor[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_547_clk_in_regs),
    .D(_03694_),
    .Q(\inst$top.soc.cpu.divider.divisor[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_709_clk_in_regs),
    .D(_03695_),
    .Q(\inst$top.soc.cpu.divider.divisor[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[27]$_SDFFE_PP0P_  (.CLK(clknet_6_18__leaf_clk_in_regs),
    .D(_03696_),
    .Q(\inst$top.soc.cpu.divider.divisor[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[28]$_SDFFE_PP0P_  (.CLK(clknet_6_21__leaf_clk_in_regs),
    .D(_03697_),
    .Q(\inst$top.soc.cpu.divider.divisor[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_546_clk_in_regs),
    .D(_03698_),
    .Q(\inst$top.soc.cpu.divider.divisor[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[2]$_SDFFE_PP0P_  (.CLK(clknet_6_20__leaf_clk_in_regs),
    .D(_03699_),
    .Q(\inst$top.soc.cpu.divider.divisor[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_547_clk_in_regs),
    .D(_03700_),
    .Q(\inst$top.soc.cpu.divider.divisor[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_549_clk_in_regs),
    .D(_03701_),
    .Q(\inst$top.soc.cpu.divider.divisor[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_671_clk_in_regs),
    .D(_03702_),
    .Q(\inst$top.soc.cpu.divider.divisor[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_550_clk_in_regs),
    .D(_03703_),
    .Q(\inst$top.soc.cpu.divider.divisor[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_550_clk_in_regs),
    .D(_03704_),
    .Q(\inst$top.soc.cpu.divider.divisor[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_696_clk_in_regs),
    .D(_03705_),
    .Q(\inst$top.soc.cpu.divider.divisor[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_701_clk_in_regs),
    .D(_03706_),
    .Q(\inst$top.soc.cpu.divider.divisor[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_701_clk_in_regs),
    .D(_03707_),
    .Q(\inst$top.soc.cpu.divider.divisor[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.divisor[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_701_clk_in_regs),
    .D(_03708_),
    .Q(\inst$top.soc.cpu.divider.divisor[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.fsm_state$_SDFF_PP0_  (.CLK(clknet_leaf_675_clk_in_regs),
    .D(_03709_),
    .Q(\inst$top.soc.cpu.divider.fsm_state ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.m_modulus$_SDFFE_PP0P_  (.CLK(clknet_6_19__leaf_clk_in_regs),
    .D(_03710_),
    .Q(\inst$top.soc.cpu.divider.m_modulus ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.m_negative$_SDFFE_PP0P_  (.CLK(clknet_leaf_566_clk_in_regs),
    .D(_03711_),
    .Q(\inst$top.soc.cpu.divider.m_negative ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[0]$_SDFFE_PP0P_  (.CLK(clknet_6_18__leaf_clk_in_regs),
    .D(_03712_),
    .Q(\inst$top.soc.cpu.divider.quotient[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_698_clk_in_regs),
    .D(_03713_),
    .Q(\inst$top.soc.cpu.divider.quotient[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_691_clk_in_regs),
    .D(_03714_),
    .Q(\inst$top.soc.cpu.divider.quotient[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_682_clk_in_regs),
    .D(_03715_),
    .Q(\inst$top.soc.cpu.divider.quotient[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_682_clk_in_regs),
    .D(_03716_),
    .Q(\inst$top.soc.cpu.divider.quotient[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[14]$_SDFFE_PP0P_  (.CLK(clknet_6_16__leaf_clk_in_regs),
    .D(_03717_),
    .Q(\inst$top.soc.cpu.divider.quotient[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_675_clk_in_regs),
    .D(_03718_),
    .Q(\inst$top.soc.cpu.divider.quotient[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_681_clk_in_regs),
    .D(_03719_),
    .Q(\inst$top.soc.cpu.divider.quotient[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_681_clk_in_regs),
    .D(_03720_),
    .Q(\inst$top.soc.cpu.divider.quotient[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_680_clk_in_regs),
    .D(_03721_),
    .Q(\inst$top.soc.cpu.divider.quotient[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_684_clk_in_regs),
    .D(_03722_),
    .Q(\inst$top.soc.cpu.divider.quotient[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_689_clk_in_regs),
    .D(_03723_),
    .Q(\inst$top.soc.cpu.divider.quotient[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_690_clk_in_regs),
    .D(_03724_),
    .Q(\inst$top.soc.cpu.divider.quotient[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_690_clk_in_regs),
    .D(_03725_),
    .Q(\inst$top.soc.cpu.divider.quotient[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_684_clk_in_regs),
    .D(_03726_),
    .Q(\inst$top.soc.cpu.divider.quotient[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_686_clk_in_regs),
    .D(_03727_),
    .Q(\inst$top.soc.cpu.divider.quotient[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_684_clk_in_regs),
    .D(_03728_),
    .Q(\inst$top.soc.cpu.divider.quotient[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_687_clk_in_regs),
    .D(_03729_),
    .Q(\inst$top.soc.cpu.divider.quotient[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_679_clk_in_regs),
    .D(_03730_),
    .Q(\inst$top.soc.cpu.divider.quotient[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_687_clk_in_regs),
    .D(_03731_),
    .Q(\inst$top.soc.cpu.divider.quotient[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_687_clk_in_regs),
    .D(_03732_),
    .Q(\inst$top.soc.cpu.divider.quotient[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_688_clk_in_regs),
    .D(_03733_),
    .Q(\inst$top.soc.cpu.divider.quotient[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_689_clk_in_regs),
    .D(_03734_),
    .Q(\inst$top.soc.cpu.divider.quotient[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_688_clk_in_regs),
    .D(_03735_),
    .Q(\inst$top.soc.cpu.divider.quotient[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_692_clk_in_regs),
    .D(_03736_),
    .Q(\inst$top.soc.cpu.divider.quotient[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_694_clk_in_regs),
    .D(_03737_),
    .Q(\inst$top.soc.cpu.divider.quotient[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_691_clk_in_regs),
    .D(_03738_),
    .Q(\inst$top.soc.cpu.divider.quotient[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_690_clk_in_regs),
    .D(_03739_),
    .Q(\inst$top.soc.cpu.divider.quotient[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_697_clk_in_regs),
    .D(_03740_),
    .Q(\inst$top.soc.cpu.divider.quotient[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_690_clk_in_regs),
    .D(_03741_),
    .Q(\inst$top.soc.cpu.divider.quotient[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_683_clk_in_regs),
    .D(_03742_),
    .Q(\inst$top.soc.cpu.divider.quotient[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.quotient[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_683_clk_in_regs),
    .D(_03743_),
    .Q(\inst$top.soc.cpu.divider.quotient[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_695_clk_in_regs),
    .D(_03744_),
    .Q(\inst$top.soc.cpu.divider.remainder[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_697_clk_in_regs),
    .D(_03745_),
    .Q(\inst$top.soc.cpu.divider.remainder[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[11]$_SDFFE_PP0P_  (.CLK(clknet_6_17__leaf_clk_in_regs),
    .D(_03746_),
    .Q(\inst$top.soc.cpu.divider.remainder[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_673_clk_in_regs),
    .D(_03747_),
    .Q(\inst$top.soc.cpu.divider.remainder[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_700_clk_in_regs),
    .D(_03748_),
    .Q(\inst$top.soc.cpu.divider.remainder[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_696_clk_in_regs),
    .D(_03749_),
    .Q(\inst$top.soc.cpu.divider.remainder[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_705_clk_in_regs),
    .D(_03750_),
    .Q(\inst$top.soc.cpu.divider.remainder[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_703_clk_in_regs),
    .D(_03751_),
    .Q(\inst$top.soc.cpu.divider.remainder[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_704_clk_in_regs),
    .D(_03752_),
    .Q(\inst$top.soc.cpu.divider.remainder[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_695_clk_in_regs),
    .D(_03753_),
    .Q(\inst$top.soc.cpu.divider.remainder[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_704_clk_in_regs),
    .D(_03754_),
    .Q(\inst$top.soc.cpu.divider.remainder[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_695_clk_in_regs),
    .D(_03755_),
    .Q(\inst$top.soc.cpu.divider.remainder[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_704_clk_in_regs),
    .D(_03756_),
    .Q(\inst$top.soc.cpu.divider.remainder[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_705_clk_in_regs),
    .D(_03757_),
    .Q(\inst$top.soc.cpu.divider.remainder[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_706_clk_in_regs),
    .D(_03758_),
    .Q(\inst$top.soc.cpu.divider.remainder[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_706_clk_in_regs),
    .D(_03759_),
    .Q(\inst$top.soc.cpu.divider.remainder[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_706_clk_in_regs),
    .D(_03760_),
    .Q(\inst$top.soc.cpu.divider.remainder[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_550_clk_in_regs),
    .D(_03761_),
    .Q(\inst$top.soc.cpu.divider.remainder[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_549_clk_in_regs),
    .D(_03762_),
    .Q(\inst$top.soc.cpu.divider.remainder[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_709_clk_in_regs),
    .D(_03763_),
    .Q(\inst$top.soc.cpu.divider.remainder[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_707_clk_in_regs),
    .D(_03764_),
    .Q(\inst$top.soc.cpu.divider.remainder[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_546_clk_in_regs),
    .D(_03765_),
    .Q(\inst$top.soc.cpu.divider.remainder[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_694_clk_in_regs),
    .D(_03766_),
    .Q(\inst$top.soc.cpu.divider.remainder[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_549_clk_in_regs),
    .D(_03767_),
    .Q(\inst$top.soc.cpu.divider.remainder[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_707_clk_in_regs),
    .D(_03768_),
    .Q(\inst$top.soc.cpu.divider.remainder[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_694_clk_in_regs),
    .D(_03769_),
    .Q(\inst$top.soc.cpu.divider.remainder[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_692_clk_in_regs),
    .D(_03770_),
    .Q(\inst$top.soc.cpu.divider.remainder[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_697_clk_in_regs),
    .D(_03771_),
    .Q(\inst$top.soc.cpu.divider.remainder[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_697_clk_in_regs),
    .D(_03772_),
    .Q(\inst$top.soc.cpu.divider.remainder[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_698_clk_in_regs),
    .D(_03773_),
    .Q(\inst$top.soc.cpu.divider.remainder[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_673_clk_in_regs),
    .D(_03774_),
    .Q(\inst$top.soc.cpu.divider.remainder[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.remainder[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_673_clk_in_regs),
    .D(_03775_),
    .Q(\inst$top.soc.cpu.divider.remainder[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.timer[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_672_clk_in_regs),
    .D(_03776_),
    .Q(\inst$top.soc.cpu.divider.timer[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.timer[1]$_SDFFE_PP0P_  (.CLK(clknet_6_16__leaf_clk_in_regs),
    .D(_03777_),
    .Q(\inst$top.soc.cpu.divider.timer[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.timer[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_672_clk_in_regs),
    .D(_03778_),
    .Q(\inst$top.soc.cpu.divider.timer[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.timer[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_671_clk_in_regs),
    .D(_03779_),
    .Q(\inst$top.soc.cpu.divider.timer[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.timer[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_671_clk_in_regs),
    .D(_03780_),
    .Q(\inst$top.soc.cpu.divider.timer[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.divider.timer[5]$_SDFFE_PP1P_  (.CLK(clknet_leaf_673_clk_in_regs),
    .D(_03781_),
    .Q(\inst$top.soc.cpu.divider.timer[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_663_clk_in_regs),
    .D(_03782_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_603_clk_in_regs),
    .D(_03783_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_652_clk_in_regs),
    .D(_03784_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_612_clk_in_regs),
    .D(_03785_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_620_clk_in_regs),
    .D(_03786_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_606_clk_in_regs),
    .D(_03787_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_606_clk_in_regs),
    .D(_03788_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_657_clk_in_regs),
    .D(_03789_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_641_clk_in_regs),
    .D(_03790_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_642_clk_in_regs),
    .D(_03791_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_642_clk_in_regs),
    .D(_03792_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_662_clk_in_regs),
    .D(_03793_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_643_clk_in_regs),
    .D(_03794_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_649_clk_in_regs),
    .D(_03795_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_685_clk_in_regs),
    .D(_03796_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_685_clk_in_regs),
    .D(_03797_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_618_clk_in_regs),
    .D(_03798_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_661_clk_in_regs),
    .D(_03799_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_685_clk_in_regs),
    .D(_03800_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_637_clk_in_regs),
    .D(_03801_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_629_clk_in_regs),
    .D(_03802_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_619_clk_in_regs),
    .D(_03803_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_737_clk_in_regs),
    .D(_03804_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_616_clk_in_regs),
    .D(_03805_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_723_clk_in_regs),
    .D(_03806_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_656_clk_in_regs),
    .D(_03807_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_721_clk_in_regs),
    .D(_03808_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_739_clk_in_regs),
    .D(_03809_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_738_clk_in_regs),
    .D(_03810_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_722_clk_in_regs),
    .D(_03811_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_610_clk_in_regs),
    .D(_03812_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_610_clk_in_regs),
    .D(_03813_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.$field.x_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause_m_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_724_clk_in_regs),
    .D(_03814_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause_m_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause_w_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_723_clk_in_regs),
    .D(_03815_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause_w_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mcause_x_select$_SDFFE_PP0P_  (.CLK(clknet_leaf_730_clk_in_regs),
    .D(_03816_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause_x_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_735_clk_in_regs),
    .D(_03817_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_612_clk_in_regs),
    .D(_03818_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_621_clk_in_regs),
    .D(_03819_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_607_clk_in_regs),
    .D(_03820_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_597_clk_in_regs),
    .D(_03821_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_652_clk_in_regs),
    .D(_03822_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_638_clk_in_regs),
    .D(_03823_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_646_clk_in_regs),
    .D(_03824_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_646_clk_in_regs),
    .D(_03825_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_645_clk_in_regs),
    .D(_03826_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_651_clk_in_regs),
    .D(_03827_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_719_clk_in_regs),
    .D(_03828_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_636_clk_in_regs),
    .D(_03829_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_636_clk_in_regs),
    .D(_03830_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_627_clk_in_regs),
    .D(_03831_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_667_clk_in_regs),
    .D(_03832_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_630_clk_in_regs),
    .D(_03833_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_630_clk_in_regs),
    .D(_03834_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_628_clk_in_regs),
    .D(_03835_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_622_clk_in_regs),
    .D(_03836_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_622_clk_in_regs),
    .D(_03837_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_733_clk_in_regs),
    .D(_03838_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_733_clk_in_regs),
    .D(_03839_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_742_clk_in_regs),
    .D(_03840_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_740_clk_in_regs),
    .D(_03841_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_721_clk_in_regs),
    .D(_03842_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_608_clk_in_regs),
    .D(_03843_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_742_clk_in_regs),
    .D(_03844_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_603_clk_in_regs),
    .D(_03845_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_653_clk_in_regs),
    .D(_03846_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc.base.x_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc_m_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_722_clk_in_regs),
    .D(_03847_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc_m_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc_w_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_723_clk_in_regs),
    .D(_03848_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc_w_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mepc_x_select$_SDFFE_PP0P_  (.CLK(clknet_leaf_731_clk_in_regs),
    .D(_03849_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mepc_x_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.meie.x_data$_SDFFE_PP0P_  (.CLK(clknet_leaf_658_clk_in_regs),
    .D(_03850_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.meie.x_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_658_clk_in_regs),
    .D(_03851_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_638_clk_in_regs),
    .D(_03852_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_637_clk_in_regs),
    .D(_03853_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_648_clk_in_regs),
    .D(_03854_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_617_clk_in_regs),
    .D(_03855_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_617_clk_in_regs),
    .D(_03856_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_659_clk_in_regs),
    .D(_03857_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_678_clk_in_regs),
    .D(_03858_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_643_clk_in_regs),
    .D(_03859_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_644_clk_in_regs),
    .D(_03860_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_665_clk_in_regs),
    .D(_03861_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_650_clk_in_regs),
    .D(_03862_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_640_clk_in_regs),
    .D(_03863_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_680_clk_in_regs),
    .D(_03864_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_649_clk_in_regs),
    .D(_03865_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_666_clk_in_regs),
    .D(_03866_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mfie.x_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.msie.x_data$_SDFFE_PP0P_  (.CLK(clknet_leaf_715_clk_in_regs),
    .D(_03867_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.msie.x_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie.mtie.x_data$_SDFFE_PP0P_  (.CLK(clknet_leaf_715_clk_in_regs),
    .D(_03868_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie.mtie.x_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie_m_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_659_clk_in_regs),
    .D(_03869_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie_m_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie_w_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_715_clk_in_regs),
    .D(_03870_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie_w_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mie_x_select$_SDFFE_PP0P_  (.CLK(clknet_leaf_731_clk_in_regs),
    .D(_03871_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mie_x_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.meip.x_data$_SDFFE_PP0P_  (.CLK(clknet_leaf_655_clk_in_regs),
    .D(_03872_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.meip.x_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_657_clk_in_regs),
    .D(_03873_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_638_clk_in_regs),
    .D(_03874_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_637_clk_in_regs),
    .D(_03875_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_637_clk_in_regs),
    .D(_03876_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_617_clk_in_regs),
    .D(_03877_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_616_clk_in_regs),
    .D(_03878_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_661_clk_in_regs),
    .D(_03879_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_642_clk_in_regs),
    .D(_03880_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_643_clk_in_regs),
    .D(_03881_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_643_clk_in_regs),
    .D(_03882_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_663_clk_in_regs),
    .D(_03883_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_649_clk_in_regs),
    .D(_03884_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_640_clk_in_regs),
    .D(_03885_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_640_clk_in_regs),
    .D(_03886_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_648_clk_in_regs),
    .D(_03887_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_669_clk_in_regs),
    .D(_03888_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mfip.x_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.msip.x_data$_SDFFE_PP0P_  (.CLK(clknet_leaf_655_clk_in_regs),
    .D(_03889_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.msip.x_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip.mtip.x_data$_SDFFE_PP0P_  (.CLK(clknet_leaf_656_clk_in_regs),
    .D(_03890_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip.mtip.x_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip_m_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_665_clk_in_regs),
    .D(_03891_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip_m_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip_w_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_665_clk_in_regs),
    .D(_03892_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip_w_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mip_x_select$_SDFFE_PP0P_  (.CLK(clknet_leaf_731_clk_in_regs),
    .D(_03893_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mip_x_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_664_clk_in_regs),
    .D(_03894_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_604_clk_in_regs),
    .D(_03895_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_718_clk_in_regs),
    .D(_03896_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[12]$_SDFFE_PP1P_  (.CLK(clknet_leaf_610_clk_in_regs),
    .D(_03897_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_615_clk_in_regs),
    .D(_03898_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_605_clk_in_regs),
    .D(_03899_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_607_clk_in_regs),
    .D(_03900_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_659_clk_in_regs),
    .D(_03901_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_641_clk_in_regs),
    .D(_03902_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_643_clk_in_regs),
    .D(_03903_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_643_clk_in_regs),
    .D(_03904_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_661_clk_in_regs),
    .D(_03905_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_665_clk_in_regs),
    .D(_03906_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_650_clk_in_regs),
    .D(_03907_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_640_clk_in_regs),
    .D(_03908_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_640_clk_in_regs),
    .D(_03909_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_617_clk_in_regs),
    .D(_03910_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_666_clk_in_regs),
    .D(_03911_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_735_clk_in_regs),
    .D(_03912_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_716_clk_in_regs),
    .D(_03913_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_733_clk_in_regs),
    .D(_03914_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_739_clk_in_regs),
    .D(_03915_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_740_clk_in_regs),
    .D(_03916_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_717_clk_in_regs),
    .D(_03917_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[8]$_SDFFE_PP1P_  (.CLK(clknet_leaf_610_clk_in_regs),
    .D(_03918_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_609_clk_in_regs),
    .D(_03919_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.ext.x_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.mxl.x_data[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_615_clk_in_regs),
    .D(_03920_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.mxl.x_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa.mxl.x_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_724_clk_in_regs),
    .D(_03921_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa.mxl.x_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa_m_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_666_clk_in_regs),
    .D(_03922_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa_m_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa_w_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_667_clk_in_regs),
    .D(_03923_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa_w_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.misa_x_select$_SDFFE_PP0P_  (.CLK(clknet_leaf_735_clk_in_regs),
    .D(_03924_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.misa_x_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_663_clk_in_regs),
    .D(_03925_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_604_clk_in_regs),
    .D(_03926_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_654_clk_in_regs),
    .D(_03927_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_612_clk_in_regs),
    .D(_03928_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_620_clk_in_regs),
    .D(_03929_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_605_clk_in_regs),
    .D(_03930_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_607_clk_in_regs),
    .D(_03931_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_660_clk_in_regs),
    .D(_03932_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_638_clk_in_regs),
    .D(_03933_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_642_clk_in_regs),
    .D(_03934_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_644_clk_in_regs),
    .D(_03935_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_661_clk_in_regs),
    .D(_03936_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_664_clk_in_regs),
    .D(_03937_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_651_clk_in_regs),
    .D(_03938_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_638_clk_in_regs),
    .D(_03939_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_635_clk_in_regs),
    .D(_03940_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_618_clk_in_regs),
    .D(_03941_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_666_clk_in_regs),
    .D(_03942_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_635_clk_in_regs),
    .D(_03943_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_637_clk_in_regs),
    .D(_03944_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_618_clk_in_regs),
    .D(_03945_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_616_clk_in_regs),
    .D(_03946_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_736_clk_in_regs),
    .D(_03947_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_616_clk_in_regs),
    .D(_03948_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_724_clk_in_regs),
    .D(_03949_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_718_clk_in_regs),
    .D(_03950_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_736_clk_in_regs),
    .D(_03951_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_739_clk_in_regs),
    .D(_03952_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_738_clk_in_regs),
    .D(_03953_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_722_clk_in_regs),
    .D(_03954_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_609_clk_in_regs),
    .D(_03955_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_742_clk_in_regs),
    .D(_03956_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch.$field.x_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch_m_select$_SDFFE_PP0N_  (.CLK(clknet_6_5__leaf_clk_in_regs),
    .D(_03957_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch_m_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch_w_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_659_clk_in_regs),
    .D(_03958_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch_w_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mscratch_x_select$_SDFFE_PP0P_  (.CLK(clknet_leaf_730_clk_in_regs),
    .D(_03959_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mscratch_x_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mstatus.mie.x_data$_SDFFE_PP0P_  (.CLK(clknet_leaf_718_clk_in_regs),
    .D(_03960_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mstatus.mie.x_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mstatus.mpie.x_data$_SDFFE_PP0P_  (.CLK(clknet_leaf_717_clk_in_regs),
    .D(_03961_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mstatus.mpie.x_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mstatus.mpp.x_data[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_719_clk_in_regs),
    .D(_03962_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mstatus.mpp.x_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mstatus.mpp.x_data[1]$_SDFFE_PP1P_  (.CLK(clknet_leaf_720_clk_in_regs),
    .D(_03963_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mstatus.mpp.x_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mstatus_m_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_715_clk_in_regs),
    .D(_03964_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mstatus_m_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mstatus_w_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_715_clk_in_regs),
    .D(_03965_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mstatus_w_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mstatus_x_select$_SDFFE_PP0P_  (.CLK(clknet_leaf_719_clk_in_regs),
    .D(_03966_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mstatus_x_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_663_clk_in_regs),
    .D(_03967_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_603_clk_in_regs),
    .D(_03968_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_653_clk_in_regs),
    .D(_03969_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_612_clk_in_regs),
    .D(_03970_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_620_clk_in_regs),
    .D(_03971_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_606_clk_in_regs),
    .D(_03972_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_597_clk_in_regs),
    .D(_03973_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_616_clk_in_regs),
    .D(_03974_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_638_clk_in_regs),
    .D(_03975_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_647_clk_in_regs),
    .D(_03976_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_647_clk_in_regs),
    .D(_03977_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_662_clk_in_regs),
    .D(_03978_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_645_clk_in_regs),
    .D(_03979_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_651_clk_in_regs),
    .D(_03980_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_636_clk_in_regs),
    .D(_03981_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_636_clk_in_regs),
    .D(_03982_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_628_clk_in_regs),
    .D(_03983_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_663_clk_in_regs),
    .D(_03984_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_636_clk_in_regs),
    .D(_03985_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_629_clk_in_regs),
    .D(_03986_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_628_clk_in_regs),
    .D(_03987_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_619_clk_in_regs),
    .D(_03988_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_735_clk_in_regs),
    .D(_03989_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_615_clk_in_regs),
    .D(_03990_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_724_clk_in_regs),
    .D(_03991_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_719_clk_in_regs),
    .D(_03992_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_733_clk_in_regs),
    .D(_03993_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_742_clk_in_regs),
    .D(_03994_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_740_clk_in_regs),
    .D(_03995_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_722_clk_in_regs),
    .D(_03996_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_608_clk_in_regs),
    .D(_03997_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_609_clk_in_regs),
    .D(_03998_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval.$field.x_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval_m_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_717_clk_in_regs),
    .D(_03999_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval_m_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval_w_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_722_clk_in_regs),
    .D(_04000_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval_w_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtval_x_select$_SDFFE_PP0P_  (.CLK(clknet_leaf_729_clk_in_regs),
    .D(_04001_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtval_x_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_734_clk_in_regs),
    .D(_04002_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_612_clk_in_regs),
    .D(_04003_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_615_clk_in_regs),
    .D(_04004_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_607_clk_in_regs),
    .D(_04005_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_607_clk_in_regs),
    .D(_04006_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_616_clk_in_regs),
    .D(_04007_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_647_clk_in_regs),
    .D(_04008_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_644_clk_in_regs),
    .D(_04009_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_645_clk_in_regs),
    .D(_04010_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_645_clk_in_regs),
    .D(_04011_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_653_clk_in_regs),
    .D(_04012_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_654_clk_in_regs),
    .D(_04013_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_636_clk_in_regs),
    .D(_04014_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[21]$_SDFFE_PP0P_  (.CLK(clknet_6_29__leaf_clk_in_regs),
    .D(_04015_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_618_clk_in_regs),
    .D(_04016_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_667_clk_in_regs),
    .D(_04017_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_637_clk_in_regs),
    .D(_04018_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_637_clk_in_regs),
    .D(_04019_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_618_clk_in_regs),
    .D(_04020_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_620_clk_in_regs),
    .D(_04021_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_615_clk_in_regs),
    .D(_04022_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_733_clk_in_regs),
    .D(_04023_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_733_clk_in_regs),
    .D(_04024_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_741_clk_in_regs),
    .D(_04025_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_740_clk_in_regs),
    .D(_04026_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_722_clk_in_regs),
    .D(_04027_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_608_clk_in_regs),
    .D(_04028_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_742_clk_in_regs),
    .D(_04029_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_611_clk_in_regs),
    .D(_04030_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_654_clk_in_regs),
    .D(_04031_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.base.x_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.mode.x_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_664_clk_in_regs),
    .D(_04032_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.mode.x_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec.mode.x_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_661_clk_in_regs),
    .D(_04033_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec.mode.x_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec_m_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_659_clk_in_regs),
    .D(_04034_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec_m_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec_w_select$_SDFFE_PP0N_  (.CLK(clknet_leaf_659_clk_in_regs),
    .D(_04035_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec_w_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.csr_bank.mtvec_x_select$_SDFFE_PP0P_  (.CLK(clknet_leaf_731_clk_in_regs),
    .D(_04036_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mtvec_x_select ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_658_clk_in_regs),
    .D(_04037_),
    .Q(\inst$top.soc.cpu.exception.m_mie.msie ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[10]$_SDFFE_PP0N_  (.CLK(clknet_leaf_679_clk_in_regs),
    .D(_04038_),
    .Q(\inst$top.soc.cpu.exception.m_mie[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[11]$_SDFFE_PP0N_  (.CLK(clknet_leaf_648_clk_in_regs),
    .D(_04039_),
    .Q(\inst$top.soc.cpu.exception.m_mie[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[12]$_SDFFE_PP0N_  (.CLK(clknet_leaf_666_clk_in_regs),
    .D(_04040_),
    .Q(\inst$top.soc.cpu.exception.m_mie[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[13]$_SDFFE_PP0N_  (.CLK(clknet_leaf_638_clk_in_regs),
    .D(_04041_),
    .Q(\inst$top.soc.cpu.exception.m_mie[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[14]$_SDFFE_PP0N_  (.CLK(clknet_leaf_638_clk_in_regs),
    .D(_04042_),
    .Q(\inst$top.soc.cpu.exception.m_mie[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[15]$_SDFFE_PP0N_  (.CLK(clknet_leaf_648_clk_in_regs),
    .D(_04043_),
    .Q(\inst$top.soc.cpu.exception.m_mie[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[16]$_SDFFE_PP0N_  (.CLK(clknet_leaf_617_clk_in_regs),
    .D(_04044_),
    .Q(\inst$top.soc.cpu.exception.m_mie[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[17]$_SDFFE_PP0N_  (.CLK(clknet_leaf_649_clk_in_regs),
    .D(_04045_),
    .Q(\inst$top.soc.cpu.exception.m_mie[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[18]$_SDFFE_PP0N_  (.CLK(clknet_leaf_659_clk_in_regs),
    .D(_04046_),
    .Q(\inst$top.soc.cpu.exception.m_mie[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_658_clk_in_regs),
    .D(_04047_),
    .Q(\inst$top.soc.cpu.exception.m_mie.mtie ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_658_clk_in_regs),
    .D(_04048_),
    .Q(\inst$top.soc.cpu.exception.m_mie.meie ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_658_clk_in_regs),
    .D(_04049_),
    .Q(\inst$top.soc.cpu.exception.m_mie[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_642_clk_in_regs),
    .D(_04050_),
    .Q(\inst$top.soc.cpu.exception.m_mie[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[5]$_SDFFE_PP0N_  (.CLK(clknet_6_16__leaf_clk_in_regs),
    .D(_04051_),
    .Q(\inst$top.soc.cpu.exception.m_mie[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[6]$_SDFFE_PP0N_  (.CLK(clknet_leaf_644_clk_in_regs),
    .D(_04052_),
    .Q(\inst$top.soc.cpu.exception.m_mie[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[7]$_SDFFE_PP0N_  (.CLK(clknet_leaf_664_clk_in_regs),
    .D(_04053_),
    .Q(\inst$top.soc.cpu.exception.m_mie[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[8]$_SDFFE_PP0N_  (.CLK(clknet_leaf_650_clk_in_regs),
    .D(_04054_),
    .Q(\inst$top.soc.cpu.exception.m_mie[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mie[9]$_SDFFE_PP0N_  (.CLK(clknet_leaf_679_clk_in_regs),
    .D(_04055_),
    .Q(\inst$top.soc.cpu.exception.m_mie[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_655_clk_in_regs),
    .D(_04056_),
    .Q(\inst$top.soc.cpu.exception.m_mip.msip ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[10]$_SDFFE_PP0N_  (.CLK(clknet_leaf_679_clk_in_regs),
    .D(_04057_),
    .Q(\inst$top.soc.cpu.exception.m_mip[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[11]$_SDFFE_PP0N_  (.CLK(clknet_leaf_648_clk_in_regs),
    .D(_04058_),
    .Q(\inst$top.soc.cpu.exception.m_mip[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[12]$_SDFFE_PP0N_  (.CLK(clknet_leaf_664_clk_in_regs),
    .D(_04059_),
    .Q(\inst$top.soc.cpu.exception.m_mip[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[13]$_SDFFE_PP0N_  (.CLK(clknet_leaf_638_clk_in_regs),
    .D(_04060_),
    .Q(\inst$top.soc.cpu.exception.m_mip[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[14]$_SDFFE_PP0N_  (.CLK(clknet_leaf_638_clk_in_regs),
    .D(_04061_),
    .Q(\inst$top.soc.cpu.exception.m_mip[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[15]$_SDFFE_PP0N_  (.CLK(clknet_leaf_648_clk_in_regs),
    .D(_04062_),
    .Q(\inst$top.soc.cpu.exception.m_mip[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[16]$_SDFFE_PP0N_  (.CLK(clknet_leaf_617_clk_in_regs),
    .D(_04063_),
    .Q(\inst$top.soc.cpu.exception.m_mip[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[17]$_SDFFE_PP0N_  (.CLK(clknet_leaf_649_clk_in_regs),
    .D(_04064_),
    .Q(\inst$top.soc.cpu.exception.m_mip[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[18]$_SDFFE_PP0N_  (.CLK(clknet_leaf_660_clk_in_regs),
    .D(_04065_),
    .Q(\inst$top.soc.cpu.exception.m_mip[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_657_clk_in_regs),
    .D(_04066_),
    .Q(\inst$top.soc.cpu.exception.m_mip.mtip ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_656_clk_in_regs),
    .D(_04067_),
    .Q(\inst$top.soc.cpu.exception.m_mip.meip ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_657_clk_in_regs),
    .D(_04068_),
    .Q(\inst$top.soc.cpu.exception.m_mip[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_643_clk_in_regs),
    .D(_04069_),
    .Q(\inst$top.soc.cpu.exception.m_mip[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[5]$_SDFFE_PP0N_  (.CLK(clknet_6_16__leaf_clk_in_regs),
    .D(_04070_),
    .Q(\inst$top.soc.cpu.exception.m_mip[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[6]$_SDFFE_PP0N_  (.CLK(clknet_leaf_643_clk_in_regs),
    .D(_04071_),
    .Q(\inst$top.soc.cpu.exception.m_mip[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[7]$_SDFFE_PP0N_  (.CLK(clknet_leaf_664_clk_in_regs),
    .D(_04072_),
    .Q(\inst$top.soc.cpu.exception.m_mip[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[8]$_SDFFE_PP0N_  (.CLK(clknet_leaf_650_clk_in_regs),
    .D(_04073_),
    .Q(\inst$top.soc.cpu.exception.m_mip[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mip[9]$_SDFFE_PP0N_  (.CLK(clknet_leaf_640_clk_in_regs),
    .D(_04074_),
    .Q(\inst$top.soc.cpu.exception.m_mip[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mstatus[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_715_clk_in_regs),
    .D(_04075_),
    .Q(\inst$top.soc.cpu.exception.m_mstatus.mie ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.m_mstatus[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_716_clk_in_regs),
    .D(_04076_),
    .Q(\inst$top.soc.cpu.exception.m_mstatus.mpie ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$48[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_662_clk_in_regs),
    .D(_04077_),
    .Q(\inst$top.soc.cpu.exception.w_data$48[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$48[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_656_clk_in_regs),
    .D(_04078_),
    .Q(\inst$top.soc.cpu.exception.w_data$48[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$48[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_656_clk_in_regs),
    .D(_04079_),
    .Q(\inst$top.soc.cpu.exception.w_data$48[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$48[31]$_SDFFE_PP0N_  (.CLK(clknet_leaf_722_clk_in_regs),
    .D(_04080_),
    .Q(\inst$top.soc.cpu.exception.w_data$48[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$48[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_656_clk_in_regs),
    .D(_04081_),
    .Q(\inst$top.soc.cpu.exception.w_data$48[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$48[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_720_clk_in_regs),
    .D(_04082_),
    .Q(\inst$top.soc.cpu.exception.w_data$48[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_739_clk_in_regs),
    .D(_04083_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[10]$_SDFFE_PP0N_  (.CLK(clknet_leaf_602_clk_in_regs),
    .D(_04084_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[11]$_SDFFE_PP0N_  (.CLK(clknet_leaf_613_clk_in_regs),
    .D(_04085_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[12]$_SDFFE_PP0N_  (.CLK(clknet_leaf_611_clk_in_regs),
    .D(_04086_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[13]$_SDFFE_PP0N_  (.CLK(clknet_leaf_621_clk_in_regs),
    .D(_04087_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[14]$_SDFFE_PP0N_  (.CLK(clknet_leaf_597_clk_in_regs),
    .D(_04088_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[15]$_SDFFE_PP0N_  (.CLK(clknet_leaf_597_clk_in_regs),
    .D(_04089_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[16]$_SDFFE_PP0N_  (.CLK(clknet_leaf_614_clk_in_regs),
    .D(_04090_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[17]$_SDFFE_PP0N_  (.CLK(clknet_leaf_648_clk_in_regs),
    .D(_04091_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[18]$_SDFFE_PP0N_  (.CLK(clknet_leaf_646_clk_in_regs),
    .D(_04092_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[19]$_SDFFE_PP0N_  (.CLK(clknet_leaf_649_clk_in_regs),
    .D(_04093_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_612_clk_in_regs),
    .D(_04094_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[20]$_SDFFE_PP0N_  (.CLK(clknet_leaf_646_clk_in_regs),
    .D(_04095_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[21]$_SDFFE_PP0N_  (.CLK(clknet_leaf_614_clk_in_regs),
    .D(_04096_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[22]$_SDFFE_PP0N_  (.CLK(clknet_leaf_629_clk_in_regs),
    .D(_04097_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[23]$_SDFFE_PP0N_  (.CLK(clknet_leaf_630_clk_in_regs),
    .D(_04098_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[24]$_SDFFE_PP0N_  (.CLK(clknet_leaf_619_clk_in_regs),
    .D(_04099_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[25]$_SDFFE_PP0N_  (.CLK(clknet_leaf_660_clk_in_regs),
    .D(_04100_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[26]$_SDFFE_PP0N_  (.CLK(clknet_leaf_630_clk_in_regs),
    .D(_04101_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[27]$_SDFFE_PP0N_  (.CLK(clknet_leaf_627_clk_in_regs),
    .D(_04102_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[28]$_SDFFE_PP0N_  (.CLK(clknet_leaf_627_clk_in_regs),
    .D(_04103_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[29]$_SDFFE_PP0N_  (.CLK(clknet_leaf_620_clk_in_regs),
    .D(_04104_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_735_clk_in_regs),
    .D(_04105_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[30]$_SDFFE_PP0N_  (.CLK(clknet_leaf_604_clk_in_regs),
    .D(_04106_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[31]$_SDFFE_PP0N_  (.CLK(clknet_leaf_732_clk_in_regs),
    .D(_04107_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_720_clk_in_regs),
    .D(_04108_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_734_clk_in_regs),
    .D(_04109_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_742_clk_in_regs),
    .D(_04110_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[6]$_SDFFE_PP0N_  (.CLK(clknet_leaf_740_clk_in_regs),
    .D(_04111_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[7]$_SDFFE_PP0N_  (.CLK(clknet_leaf_721_clk_in_regs),
    .D(_04112_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[8]$_SDFFE_PP0N_  (.CLK(clknet_leaf_608_clk_in_regs),
    .D(_04113_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_data$51[9]$_SDFFE_PP0N_  (.CLK(clknet_leaf_743_clk_in_regs),
    .D(_04114_),
    .Q(\inst$top.soc.cpu.exception.w_data$51[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_mret$_SDFFE_PP0N_  (.CLK(clknet_leaf_718_clk_in_regs),
    .D(_04115_),
    .Q(\inst$top.soc.cpu.exception.w_mret ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_mstatus[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_715_clk_in_regs),
    .D(_04116_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mstatus.mpie.w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_mstatus[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_716_clk_in_regs),
    .D(_04117_),
    .Q(\inst$top.soc.cpu.exception.w_mstatus.mpie ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.exception.w_trap$_SDFFE_PP0N_  (.CLK(clknet_leaf_737_clk_in_regs),
    .D(_04118_),
    .Q(\inst$top.soc.cpu.exception.w_trap ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.f.source__valid$_SDFFE_PP0P_  (.CLK(clknet_leaf_776_clk_in_regs),
    .D(_04119_),
    .Q(\inst$top.soc.cpu.f.source__valid ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_774_clk_in_regs),
    .D(_04120_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_769_clk_in_regs),
    .D(_04121_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_11_clk_in_regs),
    .D(_04122_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_768_clk_in_regs),
    .D(_04123_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_14_clk_in_regs),
    .D(_04124_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk_in_regs),
    .D(_04125_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_11_clk_in_regs),
    .D(_04126_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_773_clk_in_regs),
    .D(_04127_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk_in_regs),
    .D(_04128_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_766_clk_in_regs),
    .D(_04129_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_769_clk_in_regs),
    .D(_04130_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_774_clk_in_regs),
    .D(_04131_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_14_clk_in_regs),
    .D(_04132_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_14_clk_in_regs),
    .D(_04133_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_15_clk_in_regs),
    .D(_04134_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk_in_regs),
    .D(_04135_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_16_clk_in_regs),
    .D(_04136_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk_in_regs),
    .D(_04137_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk_in_regs),
    .D(_04138_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_17_clk_in_regs),
    .D(_04139_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_17_clk_in_regs),
    .D(_04140_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_774_clk_in_regs),
    .D(_04141_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[2]$_SDFFE_PP0P_  (.CLK(clknet_6_8__leaf_clk_in_regs),
    .D(_04142_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_772_clk_in_regs),
    .D(_04143_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_770_clk_in_regs),
    .D(_04144_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_765_clk_in_regs),
    .D(_04145_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk_in_regs),
    .D(_04146_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk_in_regs),
    .D(_04147_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk_in_regs),
    .D(_04148_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__adr[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_772_clk_in_regs),
    .D(_04149_),
    .Q(\inst$top.soc.cpu.fetch.ibus__adr[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__cyc$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk_in_regs),
    .D(_04150_),
    .Q(\inst$top.soc.cpu.fetch.ibus__cyc ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus__stb$_SDFFE_PP0P_  (.CLK(clknet_leaf_37_clk_in_regs),
    .D(_04151_),
    .Q(\inst$top.soc.cpu.fetch.ibus__stb ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk_in_regs),
    .D(_04152_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_317_clk_in_regs),
    .D(_04153_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_316_clk_in_regs),
    .D(_04154_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk_in_regs),
    .D(_04155_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk_in_regs),
    .D(_04156_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk_in_regs),
    .D(_04157_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk_in_regs),
    .D(_04158_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_271_clk_in_regs),
    .D(_04159_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_274_clk_in_regs),
    .D(_04160_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk_in_regs),
    .D(_04161_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_312_clk_in_regs),
    .D(_04162_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk_in_regs),
    .D(_04163_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk_in_regs),
    .D(_04164_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk_in_regs),
    .D(_04165_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_272_clk_in_regs),
    .D(_04166_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_38_clk_in_regs),
    .D(_04167_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk_in_regs),
    .D(_04168_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_36_clk_in_regs),
    .D(_04169_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk_in_regs),
    .D(_04170_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk_in_regs),
    .D(_04171_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_31_clk_in_regs),
    .D(_04172_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_36_clk_in_regs),
    .D(_04173_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk_in_regs),
    .D(_04174_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk_in_regs),
    .D(_04175_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk_in_regs),
    .D(_04176_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk_in_regs),
    .D(_04177_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk_in_regs),
    .D(_04178_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_31_clk_in_regs),
    .D(_04179_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk_in_regs),
    .D(_04180_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_313_clk_in_regs),
    .D(_04181_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_316_clk_in_regs),
    .D(_04182_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.fetch.ibus_rdata[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk_in_regs),
    .D(_04183_),
    .Q(\inst$top.soc.cpu.fetch.ibus_rdata[9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk_in_regs),
    .D(net1064),
    .DE(net1377),
    .Q(\inst$top.soc.cpu.gprf.mem[0][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_443_clk_in_regs),
    .D(net995),
    .DE(net1379),
    .Q(\inst$top.soc.cpu.gprf.mem[0][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_412_clk_in_regs),
    .D(net992),
    .DE(net1377),
    .Q(\inst$top.soc.cpu.gprf.mem[0][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_499_clk_in_regs),
    .D(net986),
    .DE(net1378),
    .Q(\inst$top.soc.cpu.gprf.mem[0][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk_in_regs),
    .D(net980),
    .DE(net1377),
    .Q(\inst$top.soc.cpu.gprf.mem[0][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk_in_regs),
    .D(net978),
    .DE(net1378),
    .Q(\inst$top.soc.cpu.gprf.mem[0][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_467_clk_in_regs),
    .D(net889),
    .DE(net1378),
    .Q(\inst$top.soc.cpu.gprf.mem[0][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_494_clk_in_regs),
    .D(net972),
    .DE(net1378),
    .Q(\inst$top.soc.cpu.gprf.mem[0][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_476_clk_in_regs),
    .D(net970),
    .DE(net1378),
    .Q(\inst$top.soc.cpu.gprf.mem[0][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_364_clk_in_regs),
    .D(net965),
    .DE(net1377),
    .Q(\inst$top.soc.cpu.gprf.mem[0][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_465_clk_in_regs),
    .D(net961),
    .DE(net1378),
    .Q(\inst$top.soc.cpu.gprf.mem[0][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk_in_regs),
    .D(net1017),
    .DE(net1377),
    .Q(\inst$top.soc.cpu.gprf.mem[0][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_401_clk_in_regs),
    .D(net954),
    .DE(net1379),
    .Q(\inst$top.soc.cpu.gprf.mem[0][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_463_clk_in_regs),
    .D(net949),
    .DE(net1380),
    .Q(\inst$top.soc.cpu.gprf.mem[0][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_416_clk_in_regs),
    .D(net944),
    .DE(net1377),
    .Q(\inst$top.soc.cpu.gprf.mem[0][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_399_clk_in_regs),
    .D(net940),
    .DE(net1377),
    .Q(\inst$top.soc.cpu.gprf.mem[0][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_499_clk_in_regs),
    .D(net935),
    .DE(net1379),
    .Q(\inst$top.soc.cpu.gprf.mem[0][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk_in_regs),
    .D(net929),
    .DE(net1379),
    .Q(\inst$top.soc.cpu.gprf.mem[0][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk_in_regs),
    .D(net925),
    .DE(net1377),
    .Q(\inst$top.soc.cpu.gprf.mem[0][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk_in_regs),
    .D(net920),
    .DE(net1378),
    .Q(\inst$top.soc.cpu.gprf.mem[0][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk_in_regs),
    .D(net918),
    .DE(net1378),
    .Q(\inst$top.soc.cpu.gprf.mem[0][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_510_clk_in_regs),
    .D(net911),
    .DE(net1379),
    .Q(\inst$top.soc.cpu.gprf.mem[0][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk_in_regs),
    .D(net1062),
    .DE(net1377),
    .Q(\inst$top.soc.cpu.gprf.mem[0][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_430_clk_in_regs),
    .D(net906),
    .DE(net1377),
    .Q(\inst$top.soc.cpu.gprf.mem[0][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_448_clk_in_regs),
    .D(net901),
    .DE(net1379),
    .Q(\inst$top.soc.cpu.gprf.mem[0][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk_in_regs),
    .D(net1056),
    .DE(net1378),
    .Q(\inst$top.soc.cpu.gprf.mem[0][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk_in_regs),
    .D(net1010),
    .DE(net1380),
    .Q(\inst$top.soc.cpu.gprf.mem[0][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk_in_regs),
    .D(net1053),
    .DE(net1379),
    .Q(\inst$top.soc.cpu.gprf.mem[0][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk_in_regs),
    .D(net1048),
    .DE(net1379),
    .Q(\inst$top.soc.cpu.gprf.mem[0][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk_in_regs),
    .D(net890),
    .DE(net1378),
    .Q(\inst$top.soc.cpu.gprf.mem[0][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk_in_regs),
    .D(net1005),
    .DE(net1380),
    .Q(\inst$top.soc.cpu.gprf.mem[0][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_436_clk_in_regs),
    .D(net999),
    .DE(net1379),
    .Q(\inst$top.soc.cpu.gprf.mem[0][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk_in_regs),
    .D(net1065),
    .DE(net1564),
    .Q(\inst$top.soc.cpu.gprf.mem[10][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_444_clk_in_regs),
    .D(net996),
    .DE(net1566),
    .Q(\inst$top.soc.cpu.gprf.mem[10][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_410_clk_in_regs),
    .D(net989),
    .DE(net1564),
    .Q(\inst$top.soc.cpu.gprf.mem[10][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][12]$_DFFE_PP_  (.CLK(clknet_leaf_500_clk_in_regs),
    .D(net985),
    .DE(net1565),
    .Q(\inst$top.soc.cpu.gprf.mem[10][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][13]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk_in_regs),
    .D(net980),
    .DE(net1564),
    .Q(\inst$top.soc.cpu.gprf.mem[10][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][14]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk_in_regs),
    .D(net976),
    .DE(net1565),
    .Q(\inst$top.soc.cpu.gprf.mem[10][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][15]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk_in_regs),
    .D(net887),
    .DE(net1565),
    .Q(\inst$top.soc.cpu.gprf.mem[10][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][16]$_DFFE_PP_  (.CLK(clknet_leaf_495_clk_in_regs),
    .D(net972),
    .DE(net1565),
    .Q(\inst$top.soc.cpu.gprf.mem[10][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][17]$_DFFE_PP_  (.CLK(clknet_leaf_478_clk_in_regs),
    .D(net967),
    .DE(net1565),
    .Q(\inst$top.soc.cpu.gprf.mem[10][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][18]$_DFFE_PP_  (.CLK(clknet_leaf_423_clk_in_regs),
    .D(net964),
    .DE(net1564),
    .Q(\inst$top.soc.cpu.gprf.mem[10][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][19]$_DFFE_PP_  (.CLK(clknet_leaf_472_clk_in_regs),
    .D(net959),
    .DE(net1565),
    .Q(\inst$top.soc.cpu.gprf.mem[10][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk_in_regs),
    .D(net1015),
    .DE(net1564),
    .Q(\inst$top.soc.cpu.gprf.mem[10][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][20]$_DFFE_PP_  (.CLK(clknet_leaf_402_clk_in_regs),
    .D(net953),
    .DE(net1564),
    .Q(\inst$top.soc.cpu.gprf.mem[10][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][21]$_DFFE_PP_  (.CLK(clknet_leaf_488_clk_in_regs),
    .D(net949),
    .DE(net1566),
    .Q(\inst$top.soc.cpu.gprf.mem[10][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][22]$_DFFE_PP_  (.CLK(clknet_leaf_421_clk_in_regs),
    .D(net944),
    .DE(net1564),
    .Q(\inst$top.soc.cpu.gprf.mem[10][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][23]$_DFFE_PP_  (.CLK(clknet_leaf_405_clk_in_regs),
    .D(net939),
    .DE(net1564),
    .Q(\inst$top.soc.cpu.gprf.mem[10][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][24]$_DFFE_PP_  (.CLK(clknet_leaf_503_clk_in_regs),
    .D(net936),
    .DE(net1566),
    .Q(\inst$top.soc.cpu.gprf.mem[10][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][25]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk_in_regs),
    .D(net930),
    .DE(net1566),
    .Q(\inst$top.soc.cpu.gprf.mem[10][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][26]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk_in_regs),
    .D(net925),
    .DE(net1564),
    .Q(\inst$top.soc.cpu.gprf.mem[10][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][27]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk_in_regs),
    .D(net921),
    .DE(net1565),
    .Q(\inst$top.soc.cpu.gprf.mem[10][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][28]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk_in_regs),
    .D(net917),
    .DE(net1565),
    .Q(\inst$top.soc.cpu.gprf.mem[10][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][29]$_DFFE_PP_  (.CLK(clknet_leaf_509_clk_in_regs),
    .D(net911),
    .DE(net1566),
    .Q(\inst$top.soc.cpu.gprf.mem[10][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk_in_regs),
    .D(net1060),
    .DE(net1564),
    .Q(\inst$top.soc.cpu.gprf.mem[10][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][30]$_DFFE_PP_  (.CLK(clknet_leaf_434_clk_in_regs),
    .D(net907),
    .DE(net1567),
    .Q(\inst$top.soc.cpu.gprf.mem[10][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][31]$_DFFE_PP_  (.CLK(clknet_leaf_454_clk_in_regs),
    .D(net901),
    .DE(net1566),
    .Q(\inst$top.soc.cpu.gprf.mem[10][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk_in_regs),
    .D(net1057),
    .DE(net1565),
    .Q(\inst$top.soc.cpu.gprf.mem[10][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk_in_regs),
    .D(net1010),
    .DE(net1567),
    .Q(\inst$top.soc.cpu.gprf.mem[10][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk_in_regs),
    .D(net1052),
    .DE(net1566),
    .Q(\inst$top.soc.cpu.gprf.mem[10][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk_in_regs),
    .D(net1048),
    .DE(net1567),
    .Q(\inst$top.soc.cpu.gprf.mem[10][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk_in_regs),
    .D(net892),
    .DE(net1565),
    .Q(\inst$top.soc.cpu.gprf.mem[10][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk_in_regs),
    .D(net1004),
    .DE(net1567),
    .Q(\inst$top.soc.cpu.gprf.mem[10][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk_in_regs),
    .D(net1000),
    .DE(net1566),
    .Q(\inst$top.soc.cpu.gprf.mem[10][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk_in_regs),
    .D(net1066),
    .DE(net1560),
    .Q(\inst$top.soc.cpu.gprf.mem[11][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_444_clk_in_regs),
    .D(net996),
    .DE(net1562),
    .Q(\inst$top.soc.cpu.gprf.mem[11][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_410_clk_in_regs),
    .D(net990),
    .DE(net1560),
    .Q(\inst$top.soc.cpu.gprf.mem[11][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][12]$_DFFE_PP_  (.CLK(clknet_leaf_500_clk_in_regs),
    .D(net985),
    .DE(net1561),
    .Q(\inst$top.soc.cpu.gprf.mem[11][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][13]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk_in_regs),
    .D(net980),
    .DE(net1560),
    .Q(\inst$top.soc.cpu.gprf.mem[11][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][14]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk_in_regs),
    .D(net976),
    .DE(net1561),
    .Q(\inst$top.soc.cpu.gprf.mem[11][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][15]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk_in_regs),
    .D(net887),
    .DE(net1561),
    .Q(\inst$top.soc.cpu.gprf.mem[11][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][16]$_DFFE_PP_  (.CLK(clknet_leaf_497_clk_in_regs),
    .D(net972),
    .DE(net1561),
    .Q(\inst$top.soc.cpu.gprf.mem[11][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][17]$_DFFE_PP_  (.CLK(clknet_leaf_477_clk_in_regs),
    .D(net967),
    .DE(net1561),
    .Q(\inst$top.soc.cpu.gprf.mem[11][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][18]$_DFFE_PP_  (.CLK(clknet_leaf_423_clk_in_regs),
    .D(net964),
    .DE(net1560),
    .Q(\inst$top.soc.cpu.gprf.mem[11][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][19]$_DFFE_PP_  (.CLK(clknet_leaf_473_clk_in_regs),
    .D(net959),
    .DE(net1561),
    .Q(\inst$top.soc.cpu.gprf.mem[11][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk_in_regs),
    .D(net1015),
    .DE(net1560),
    .Q(\inst$top.soc.cpu.gprf.mem[11][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][20]$_DFFE_PP_  (.CLK(clknet_leaf_400_clk_in_regs),
    .D(net956),
    .DE(net1560),
    .Q(\inst$top.soc.cpu.gprf.mem[11][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][21]$_DFFE_PP_  (.CLK(clknet_leaf_487_clk_in_regs),
    .D(net950),
    .DE(net1562),
    .Q(\inst$top.soc.cpu.gprf.mem[11][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][22]$_DFFE_PP_  (.CLK(clknet_6_52__leaf_clk_in_regs),
    .D(net944),
    .DE(net1560),
    .Q(\inst$top.soc.cpu.gprf.mem[11][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][23]$_DFFE_PP_  (.CLK(clknet_leaf_400_clk_in_regs),
    .D(net939),
    .DE(net1560),
    .Q(\inst$top.soc.cpu.gprf.mem[11][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][24]$_DFFE_PP_  (.CLK(clknet_leaf_501_clk_in_regs),
    .D(net936),
    .DE(net1562),
    .Q(\inst$top.soc.cpu.gprf.mem[11][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][25]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk_in_regs),
    .D(net931),
    .DE(net1562),
    .Q(\inst$top.soc.cpu.gprf.mem[11][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][26]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk_in_regs),
    .D(net925),
    .DE(net1560),
    .Q(\inst$top.soc.cpu.gprf.mem[11][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][27]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk_in_regs),
    .D(net921),
    .DE(net1561),
    .Q(\inst$top.soc.cpu.gprf.mem[11][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][28]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk_in_regs),
    .D(net917),
    .DE(net1561),
    .Q(\inst$top.soc.cpu.gprf.mem[11][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][29]$_DFFE_PP_  (.CLK(clknet_leaf_494_clk_in_regs),
    .D(net913),
    .DE(net1562),
    .Q(\inst$top.soc.cpu.gprf.mem[11][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk_in_regs),
    .D(net1060),
    .DE(net1560),
    .Q(\inst$top.soc.cpu.gprf.mem[11][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][30]$_DFFE_PP_  (.CLK(clknet_leaf_432_clk_in_regs),
    .D(net907),
    .DE(net1563),
    .Q(\inst$top.soc.cpu.gprf.mem[11][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][31]$_DFFE_PP_  (.CLK(clknet_leaf_454_clk_in_regs),
    .D(net901),
    .DE(net1562),
    .Q(\inst$top.soc.cpu.gprf.mem[11][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk_in_regs),
    .D(net1058),
    .DE(net1561),
    .Q(\inst$top.soc.cpu.gprf.mem[11][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk_in_regs),
    .D(net1010),
    .DE(net1563),
    .Q(\inst$top.soc.cpu.gprf.mem[11][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk_in_regs),
    .D(net1052),
    .DE(net1562),
    .Q(\inst$top.soc.cpu.gprf.mem[11][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk_in_regs),
    .D(net1048),
    .DE(net1563),
    .Q(\inst$top.soc.cpu.gprf.mem[11][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk_in_regs),
    .D(net892),
    .DE(net1561),
    .Q(\inst$top.soc.cpu.gprf.mem[11][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk_in_regs),
    .D(net1005),
    .DE(net1563),
    .Q(\inst$top.soc.cpu.gprf.mem[11][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk_in_regs),
    .D(net1001),
    .DE(net1562),
    .Q(\inst$top.soc.cpu.gprf.mem[11][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk_in_regs),
    .D(net1065),
    .DE(net1580),
    .Q(\inst$top.soc.cpu.gprf.mem[12][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_439_clk_in_regs),
    .D(net996),
    .DE(net1581),
    .Q(\inst$top.soc.cpu.gprf.mem[12][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_410_clk_in_regs),
    .D(net989),
    .DE(net1580),
    .Q(\inst$top.soc.cpu.gprf.mem[12][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][12]$_DFFE_PP_  (.CLK(clknet_leaf_482_clk_in_regs),
    .D(net984),
    .DE(net1582),
    .Q(\inst$top.soc.cpu.gprf.mem[12][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][13]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk_in_regs),
    .D(net983),
    .DE(net1580),
    .Q(\inst$top.soc.cpu.gprf.mem[12][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][14]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk_in_regs),
    .D(net976),
    .DE(net1582),
    .Q(\inst$top.soc.cpu.gprf.mem[12][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][15]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk_in_regs),
    .D(net887),
    .DE(net1582),
    .Q(\inst$top.soc.cpu.gprf.mem[12][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][16]$_DFFE_PP_  (.CLK(clknet_leaf_490_clk_in_regs),
    .D(net973),
    .DE(net1581),
    .Q(\inst$top.soc.cpu.gprf.mem[12][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][17]$_DFFE_PP_  (.CLK(clknet_leaf_478_clk_in_regs),
    .D(net967),
    .DE(net1582),
    .Q(\inst$top.soc.cpu.gprf.mem[12][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][18]$_DFFE_PP_  (.CLK(clknet_leaf_423_clk_in_regs),
    .D(net964),
    .DE(net1580),
    .Q(\inst$top.soc.cpu.gprf.mem[12][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][19]$_DFFE_PP_  (.CLK(clknet_leaf_471_clk_in_regs),
    .D(net959),
    .DE(net1582),
    .Q(\inst$top.soc.cpu.gprf.mem[12][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk_in_regs),
    .D(net1016),
    .DE(net1580),
    .Q(\inst$top.soc.cpu.gprf.mem[12][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][20]$_DFFE_PP_  (.CLK(clknet_leaf_403_clk_in_regs),
    .D(net953),
    .DE(net1581),
    .Q(\inst$top.soc.cpu.gprf.mem[12][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][21]$_DFFE_PP_  (.CLK(clknet_leaf_487_clk_in_regs),
    .D(net951),
    .DE(net1582),
    .Q(\inst$top.soc.cpu.gprf.mem[12][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][22]$_DFFE_PP_  (.CLK(clknet_leaf_372_clk_in_regs),
    .D(net944),
    .DE(net1580),
    .Q(\inst$top.soc.cpu.gprf.mem[12][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][23]$_DFFE_PP_  (.CLK(clknet_leaf_406_clk_in_regs),
    .D(net942),
    .DE(net1580),
    .Q(\inst$top.soc.cpu.gprf.mem[12][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][24]$_DFFE_PP_  (.CLK(clknet_leaf_502_clk_in_regs),
    .D(net937),
    .DE(net1582),
    .Q(\inst$top.soc.cpu.gprf.mem[12][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][25]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk_in_regs),
    .D(net931),
    .DE(net1581),
    .Q(\inst$top.soc.cpu.gprf.mem[12][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][26]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk_in_regs),
    .D(net926),
    .DE(net1580),
    .Q(\inst$top.soc.cpu.gprf.mem[12][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][27]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk_in_regs),
    .D(net921),
    .DE(net1581),
    .Q(\inst$top.soc.cpu.gprf.mem[12][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][28]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk_in_regs),
    .D(net918),
    .DE(net1581),
    .Q(\inst$top.soc.cpu.gprf.mem[12][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][29]$_DFFE_PP_  (.CLK(clknet_leaf_492_clk_in_regs),
    .D(net911),
    .DE(net1581),
    .Q(\inst$top.soc.cpu.gprf.mem[12][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk_in_regs),
    .D(net1060),
    .DE(net1580),
    .Q(\inst$top.soc.cpu.gprf.mem[12][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][30]$_DFFE_PP_  (.CLK(clknet_leaf_433_clk_in_regs),
    .D(net907),
    .DE(net1580),
    .Q(\inst$top.soc.cpu.gprf.mem[12][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][31]$_DFFE_PP_  (.CLK(clknet_leaf_455_clk_in_regs),
    .D(net901),
    .DE(net1581),
    .Q(\inst$top.soc.cpu.gprf.mem[12][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk_in_regs),
    .D(net1057),
    .DE(net1582),
    .Q(\inst$top.soc.cpu.gprf.mem[12][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk_in_regs),
    .D(net1010),
    .DE(net1583),
    .Q(\inst$top.soc.cpu.gprf.mem[12][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk_in_regs),
    .D(net1053),
    .DE(net1581),
    .Q(\inst$top.soc.cpu.gprf.mem[12][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk_in_regs),
    .D(net1048),
    .DE(net1581),
    .Q(\inst$top.soc.cpu.gprf.mem[12][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk_in_regs),
    .D(net892),
    .DE(net1583),
    .Q(\inst$top.soc.cpu.gprf.mem[12][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk_in_regs),
    .D(net1004),
    .DE(net1583),
    .Q(\inst$top.soc.cpu.gprf.mem[12][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_458_clk_in_regs),
    .D(net1001),
    .DE(net1582),
    .Q(\inst$top.soc.cpu.gprf.mem[12][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk_in_regs),
    .D(net1065),
    .DE(net1597),
    .Q(\inst$top.soc.cpu.gprf.mem[13][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_439_clk_in_regs),
    .D(net996),
    .DE(net1598),
    .Q(\inst$top.soc.cpu.gprf.mem[13][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_410_clk_in_regs),
    .D(net989),
    .DE(net1597),
    .Q(\inst$top.soc.cpu.gprf.mem[13][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][12]$_DFFE_PP_  (.CLK(clknet_leaf_482_clk_in_regs),
    .D(net984),
    .DE(net1599),
    .Q(\inst$top.soc.cpu.gprf.mem[13][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][13]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk_in_regs),
    .D(net983),
    .DE(net1597),
    .Q(\inst$top.soc.cpu.gprf.mem[13][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][14]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk_in_regs),
    .D(net976),
    .DE(net1599),
    .Q(\inst$top.soc.cpu.gprf.mem[13][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][15]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk_in_regs),
    .D(net887),
    .DE(net1599),
    .Q(\inst$top.soc.cpu.gprf.mem[13][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][16]$_DFFE_PP_  (.CLK(clknet_leaf_491_clk_in_regs),
    .D(net973),
    .DE(net1598),
    .Q(\inst$top.soc.cpu.gprf.mem[13][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][17]$_DFFE_PP_  (.CLK(clknet_leaf_478_clk_in_regs),
    .D(net967),
    .DE(net1599),
    .Q(\inst$top.soc.cpu.gprf.mem[13][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][18]$_DFFE_PP_  (.CLK(clknet_leaf_423_clk_in_regs),
    .D(net965),
    .DE(net1597),
    .Q(\inst$top.soc.cpu.gprf.mem[13][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][19]$_DFFE_PP_  (.CLK(clknet_leaf_471_clk_in_regs),
    .D(net959),
    .DE(net1599),
    .Q(\inst$top.soc.cpu.gprf.mem[13][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk_in_regs),
    .D(net1016),
    .DE(net1597),
    .Q(\inst$top.soc.cpu.gprf.mem[13][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][20]$_DFFE_PP_  (.CLK(clknet_leaf_403_clk_in_regs),
    .D(net953),
    .DE(net1598),
    .Q(\inst$top.soc.cpu.gprf.mem[13][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][21]$_DFFE_PP_  (.CLK(clknet_leaf_487_clk_in_regs),
    .D(net951),
    .DE(net1599),
    .Q(\inst$top.soc.cpu.gprf.mem[13][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][22]$_DFFE_PP_  (.CLK(clknet_leaf_416_clk_in_regs),
    .D(net944),
    .DE(net1597),
    .Q(\inst$top.soc.cpu.gprf.mem[13][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][23]$_DFFE_PP_  (.CLK(clknet_leaf_406_clk_in_regs),
    .D(net942),
    .DE(net1597),
    .Q(\inst$top.soc.cpu.gprf.mem[13][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][24]$_DFFE_PP_  (.CLK(clknet_leaf_482_clk_in_regs),
    .D(net937),
    .DE(net1599),
    .Q(\inst$top.soc.cpu.gprf.mem[13][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][25]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk_in_regs),
    .D(net931),
    .DE(net1598),
    .Q(\inst$top.soc.cpu.gprf.mem[13][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][26]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk_in_regs),
    .D(net926),
    .DE(net1597),
    .Q(\inst$top.soc.cpu.gprf.mem[13][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][27]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk_in_regs),
    .D(net921),
    .DE(net1598),
    .Q(\inst$top.soc.cpu.gprf.mem[13][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][28]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk_in_regs),
    .D(net918),
    .DE(net1598),
    .Q(\inst$top.soc.cpu.gprf.mem[13][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][29]$_DFFE_PP_  (.CLK(clknet_leaf_447_clk_in_regs),
    .D(net911),
    .DE(net1598),
    .Q(\inst$top.soc.cpu.gprf.mem[13][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk_in_regs),
    .D(net1060),
    .DE(net1597),
    .Q(\inst$top.soc.cpu.gprf.mem[13][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][30]$_DFFE_PP_  (.CLK(clknet_leaf_433_clk_in_regs),
    .D(net907),
    .DE(net1597),
    .Q(\inst$top.soc.cpu.gprf.mem[13][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][31]$_DFFE_PP_  (.CLK(clknet_leaf_455_clk_in_regs),
    .D(net901),
    .DE(net1598),
    .Q(\inst$top.soc.cpu.gprf.mem[13][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk_in_regs),
    .D(net1057),
    .DE(net1599),
    .Q(\inst$top.soc.cpu.gprf.mem[13][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk_in_regs),
    .D(net1010),
    .DE(net1600),
    .Q(\inst$top.soc.cpu.gprf.mem[13][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk_in_regs),
    .D(net1053),
    .DE(net1598),
    .Q(\inst$top.soc.cpu.gprf.mem[13][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk_in_regs),
    .D(net1048),
    .DE(net1598),
    .Q(\inst$top.soc.cpu.gprf.mem[13][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk_in_regs),
    .D(net892),
    .DE(net1600),
    .Q(\inst$top.soc.cpu.gprf.mem[13][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk_in_regs),
    .D(net1004),
    .DE(net1600),
    .Q(\inst$top.soc.cpu.gprf.mem[13][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_458_clk_in_regs),
    .D(net1001),
    .DE(net1599),
    .Q(\inst$top.soc.cpu.gprf.mem[13][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk_in_regs),
    .D(net1065),
    .DE(net1588),
    .Q(\inst$top.soc.cpu.gprf.mem[14][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_439_clk_in_regs),
    .D(net996),
    .DE(net1590),
    .Q(\inst$top.soc.cpu.gprf.mem[14][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_410_clk_in_regs),
    .D(net989),
    .DE(net1589),
    .Q(\inst$top.soc.cpu.gprf.mem[14][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][12]$_DFFE_PP_  (.CLK(clknet_leaf_502_clk_in_regs),
    .D(net984),
    .DE(net1591),
    .Q(\inst$top.soc.cpu.gprf.mem[14][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][13]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk_in_regs),
    .D(net983),
    .DE(net1588),
    .Q(\inst$top.soc.cpu.gprf.mem[14][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][14]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk_in_regs),
    .D(net975),
    .DE(net1591),
    .Q(\inst$top.soc.cpu.gprf.mem[14][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][15]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk_in_regs),
    .D(net887),
    .DE(net1591),
    .Q(\inst$top.soc.cpu.gprf.mem[14][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][16]$_DFFE_PP_  (.CLK(clknet_leaf_491_clk_in_regs),
    .D(net973),
    .DE(net1590),
    .Q(\inst$top.soc.cpu.gprf.mem[14][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][17]$_DFFE_PP_  (.CLK(clknet_leaf_479_clk_in_regs),
    .D(net967),
    .DE(net1591),
    .Q(\inst$top.soc.cpu.gprf.mem[14][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][18]$_DFFE_PP_  (.CLK(clknet_leaf_423_clk_in_regs),
    .D(net965),
    .DE(net1589),
    .Q(\inst$top.soc.cpu.gprf.mem[14][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][19]$_DFFE_PP_  (.CLK(clknet_leaf_471_clk_in_regs),
    .D(net959),
    .DE(net1591),
    .Q(\inst$top.soc.cpu.gprf.mem[14][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk_in_regs),
    .D(net1016),
    .DE(net1588),
    .Q(\inst$top.soc.cpu.gprf.mem[14][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][20]$_DFFE_PP_  (.CLK(clknet_leaf_403_clk_in_regs),
    .D(net953),
    .DE(net1590),
    .Q(\inst$top.soc.cpu.gprf.mem[14][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][21]$_DFFE_PP_  (.CLK(clknet_leaf_487_clk_in_regs),
    .D(net951),
    .DE(net1591),
    .Q(\inst$top.soc.cpu.gprf.mem[14][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][22]$_DFFE_PP_  (.CLK(clknet_leaf_416_clk_in_regs),
    .D(net944),
    .DE(net1589),
    .Q(\inst$top.soc.cpu.gprf.mem[14][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][23]$_DFFE_PP_  (.CLK(clknet_leaf_406_clk_in_regs),
    .D(net939),
    .DE(net1589),
    .Q(\inst$top.soc.cpu.gprf.mem[14][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][24]$_DFFE_PP_  (.CLK(clknet_leaf_482_clk_in_regs),
    .D(net937),
    .DE(net1591),
    .Q(\inst$top.soc.cpu.gprf.mem[14][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][25]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk_in_regs),
    .D(net931),
    .DE(net1590),
    .Q(\inst$top.soc.cpu.gprf.mem[14][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][26]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk_in_regs),
    .D(net925),
    .DE(net1588),
    .Q(\inst$top.soc.cpu.gprf.mem[14][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][27]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk_in_regs),
    .D(net921),
    .DE(net1590),
    .Q(\inst$top.soc.cpu.gprf.mem[14][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][28]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk_in_regs),
    .D(net917),
    .DE(net1590),
    .Q(\inst$top.soc.cpu.gprf.mem[14][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][29]$_DFFE_PP_  (.CLK(clknet_leaf_493_clk_in_regs),
    .D(net912),
    .DE(net1590),
    .Q(\inst$top.soc.cpu.gprf.mem[14][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk_in_regs),
    .D(net1060),
    .DE(net1588),
    .Q(\inst$top.soc.cpu.gprf.mem[14][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][30]$_DFFE_PP_  (.CLK(clknet_leaf_433_clk_in_regs),
    .D(net908),
    .DE(net1589),
    .Q(\inst$top.soc.cpu.gprf.mem[14][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][31]$_DFFE_PP_  (.CLK(clknet_leaf_454_clk_in_regs),
    .D(net901),
    .DE(net1590),
    .Q(\inst$top.soc.cpu.gprf.mem[14][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk_in_regs),
    .D(net1058),
    .DE(net1591),
    .Q(\inst$top.soc.cpu.gprf.mem[14][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk_in_regs),
    .D(net1010),
    .DE(net1592),
    .Q(\inst$top.soc.cpu.gprf.mem[14][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk_in_regs),
    .D(net1052),
    .DE(net1590),
    .Q(\inst$top.soc.cpu.gprf.mem[14][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk_in_regs),
    .D(net1048),
    .DE(net1590),
    .Q(\inst$top.soc.cpu.gprf.mem[14][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk_in_regs),
    .D(net892),
    .DE(net1592),
    .Q(\inst$top.soc.cpu.gprf.mem[14][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk_in_regs),
    .D(net1004),
    .DE(net1592),
    .Q(\inst$top.soc.cpu.gprf.mem[14][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_458_clk_in_regs),
    .D(net1001),
    .DE(net1591),
    .Q(\inst$top.soc.cpu.gprf.mem[14][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk_in_regs),
    .D(net1065),
    .DE(net1552),
    .Q(\inst$top.soc.cpu.gprf.mem[15][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_439_clk_in_regs),
    .D(net996),
    .DE(net1553),
    .Q(\inst$top.soc.cpu.gprf.mem[15][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_410_clk_in_regs),
    .D(net989),
    .DE(net1552),
    .Q(\inst$top.soc.cpu.gprf.mem[15][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][12]$_DFFE_PP_  (.CLK(clknet_leaf_502_clk_in_regs),
    .D(net987),
    .DE(net1554),
    .Q(\inst$top.soc.cpu.gprf.mem[15][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][13]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk_in_regs),
    .D(net983),
    .DE(net1552),
    .Q(\inst$top.soc.cpu.gprf.mem[15][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][14]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk_in_regs),
    .D(net975),
    .DE(net1554),
    .Q(\inst$top.soc.cpu.gprf.mem[15][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][15]$_DFFE_PP_  (.CLK(clknet_leaf_471_clk_in_regs),
    .D(net887),
    .DE(net1554),
    .Q(\inst$top.soc.cpu.gprf.mem[15][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][16]$_DFFE_PP_  (.CLK(clknet_leaf_490_clk_in_regs),
    .D(net973),
    .DE(net1554),
    .Q(\inst$top.soc.cpu.gprf.mem[15][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][17]$_DFFE_PP_  (.CLK(clknet_leaf_480_clk_in_regs),
    .D(net967),
    .DE(net1554),
    .Q(\inst$top.soc.cpu.gprf.mem[15][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][18]$_DFFE_PP_  (.CLK(clknet_leaf_424_clk_in_regs),
    .D(net965),
    .DE(net1552),
    .Q(\inst$top.soc.cpu.gprf.mem[15][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][19]$_DFFE_PP_  (.CLK(clknet_leaf_471_clk_in_regs),
    .D(net959),
    .DE(net1554),
    .Q(\inst$top.soc.cpu.gprf.mem[15][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk_in_regs),
    .D(net1016),
    .DE(net1552),
    .Q(\inst$top.soc.cpu.gprf.mem[15][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][20]$_DFFE_PP_  (.CLK(clknet_leaf_402_clk_in_regs),
    .D(net953),
    .DE(net1553),
    .Q(\inst$top.soc.cpu.gprf.mem[15][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][21]$_DFFE_PP_  (.CLK(clknet_leaf_488_clk_in_regs),
    .D(net949),
    .DE(net1554),
    .Q(\inst$top.soc.cpu.gprf.mem[15][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][22]$_DFFE_PP_  (.CLK(clknet_leaf_414_clk_in_regs),
    .D(net944),
    .DE(net1552),
    .Q(\inst$top.soc.cpu.gprf.mem[15][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][23]$_DFFE_PP_  (.CLK(clknet_leaf_405_clk_in_regs),
    .D(net939),
    .DE(net1552),
    .Q(\inst$top.soc.cpu.gprf.mem[15][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][24]$_DFFE_PP_  (.CLK(clknet_leaf_502_clk_in_regs),
    .D(net937),
    .DE(net1554),
    .Q(\inst$top.soc.cpu.gprf.mem[15][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][25]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk_in_regs),
    .D(net931),
    .DE(net1553),
    .Q(\inst$top.soc.cpu.gprf.mem[15][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][26]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk_in_regs),
    .D(net926),
    .DE(net1552),
    .Q(\inst$top.soc.cpu.gprf.mem[15][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][27]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk_in_regs),
    .D(net921),
    .DE(net1553),
    .Q(\inst$top.soc.cpu.gprf.mem[15][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][28]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk_in_regs),
    .D(net917),
    .DE(net1553),
    .Q(\inst$top.soc.cpu.gprf.mem[15][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][29]$_DFFE_PP_  (.CLK(clknet_leaf_493_clk_in_regs),
    .D(net912),
    .DE(net1553),
    .Q(\inst$top.soc.cpu.gprf.mem[15][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk_in_regs),
    .D(net1060),
    .DE(net1552),
    .Q(\inst$top.soc.cpu.gprf.mem[15][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][30]$_DFFE_PP_  (.CLK(clknet_leaf_434_clk_in_regs),
    .D(net908),
    .DE(net1552),
    .Q(\inst$top.soc.cpu.gprf.mem[15][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][31]$_DFFE_PP_  (.CLK(clknet_leaf_455_clk_in_regs),
    .D(net905),
    .DE(net1553),
    .Q(\inst$top.soc.cpu.gprf.mem[15][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk_in_regs),
    .D(net1058),
    .DE(net1554),
    .Q(\inst$top.soc.cpu.gprf.mem[15][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk_in_regs),
    .D(net1010),
    .DE(net1555),
    .Q(\inst$top.soc.cpu.gprf.mem[15][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk_in_regs),
    .D(net1053),
    .DE(net1553),
    .Q(\inst$top.soc.cpu.gprf.mem[15][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk_in_regs),
    .D(net1048),
    .DE(net1553),
    .Q(\inst$top.soc.cpu.gprf.mem[15][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk_in_regs),
    .D(net892),
    .DE(net1554),
    .Q(\inst$top.soc.cpu.gprf.mem[15][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk_in_regs),
    .D(net1004),
    .DE(net1555),
    .Q(\inst$top.soc.cpu.gprf.mem[15][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_458_clk_in_regs),
    .D(net1001),
    .DE(net1553),
    .Q(\inst$top.soc.cpu.gprf.mem[15][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk_in_regs),
    .D(net1065),
    .DE(net1369),
    .Q(\inst$top.soc.cpu.gprf.mem[16][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_441_clk_in_regs),
    .D(net994),
    .DE(net1369),
    .Q(\inst$top.soc.cpu.gprf.mem[16][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_396_clk_in_regs),
    .D(net991),
    .DE(net1369),
    .Q(\inst$top.soc.cpu.gprf.mem[16][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][12]$_DFFE_PP_  (.CLK(clknet_leaf_505_clk_in_regs),
    .D(net985),
    .DE(net1371),
    .Q(\inst$top.soc.cpu.gprf.mem[16][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][13]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk_in_regs),
    .D(net983),
    .DE(net1369),
    .Q(\inst$top.soc.cpu.gprf.mem[16][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][14]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk_in_regs),
    .D(net976),
    .DE(net1371),
    .Q(\inst$top.soc.cpu.gprf.mem[16][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][15]$_DFFE_PP_  (.CLK(clknet_leaf_470_clk_in_regs),
    .D(net887),
    .DE(net1372),
    .Q(\inst$top.soc.cpu.gprf.mem[16][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][16]$_DFFE_PP_  (.CLK(clknet_leaf_506_clk_in_regs),
    .D(net972),
    .DE(net1371),
    .Q(\inst$top.soc.cpu.gprf.mem[16][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][17]$_DFFE_PP_  (.CLK(clknet_leaf_478_clk_in_regs),
    .D(net967),
    .DE(net1372),
    .Q(\inst$top.soc.cpu.gprf.mem[16][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][18]$_DFFE_PP_  (.CLK(clknet_leaf_365_clk_in_regs),
    .D(net963),
    .DE(net1369),
    .Q(\inst$top.soc.cpu.gprf.mem[16][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][19]$_DFFE_PP_  (.CLK(clknet_leaf_472_clk_in_regs),
    .D(net959),
    .DE(net1372),
    .Q(\inst$top.soc.cpu.gprf.mem[16][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk_in_regs),
    .D(net1015),
    .DE(net1369),
    .Q(\inst$top.soc.cpu.gprf.mem[16][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][20]$_DFFE_PP_  (.CLK(clknet_leaf_513_clk_in_regs),
    .D(net956),
    .DE(net1369),
    .Q(\inst$top.soc.cpu.gprf.mem[16][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][21]$_DFFE_PP_  (.CLK(clknet_leaf_450_clk_in_regs),
    .D(net952),
    .DE(net1371),
    .Q(\inst$top.soc.cpu.gprf.mem[16][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][22]$_DFFE_PP_  (.CLK(clknet_leaf_417_clk_in_regs),
    .D(net945),
    .DE(net1369),
    .Q(\inst$top.soc.cpu.gprf.mem[16][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][23]$_DFFE_PP_  (.CLK(clknet_leaf_396_clk_in_regs),
    .D(net942),
    .DE(net1370),
    .Q(\inst$top.soc.cpu.gprf.mem[16][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][24]$_DFFE_PP_  (.CLK(clknet_leaf_503_clk_in_regs),
    .D(net936),
    .DE(net1372),
    .Q(\inst$top.soc.cpu.gprf.mem[16][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][25]$_DFFE_PP_  (.CLK(clknet_leaf_435_clk_in_regs),
    .D(net932),
    .DE(net1370),
    .Q(\inst$top.soc.cpu.gprf.mem[16][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][26]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk_in_regs),
    .D(net926),
    .DE(net1369),
    .Q(\inst$top.soc.cpu.gprf.mem[16][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][27]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk_in_regs),
    .D(net920),
    .DE(net1371),
    .Q(\inst$top.soc.cpu.gprf.mem[16][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][28]$_DFFE_PP_  (.CLK(clknet_leaf_467_clk_in_regs),
    .D(net916),
    .DE(net1372),
    .Q(\inst$top.soc.cpu.gprf.mem[16][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][29]$_DFFE_PP_  (.CLK(clknet_leaf_507_clk_in_regs),
    .D(net913),
    .DE(net1371),
    .Q(\inst$top.soc.cpu.gprf.mem[16][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk_in_regs),
    .D(net1060),
    .DE(net1369),
    .Q(\inst$top.soc.cpu.gprf.mem[16][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][30]$_DFFE_PP_  (.CLK(clknet_leaf_432_clk_in_regs),
    .D(net907),
    .DE(net1370),
    .Q(\inst$top.soc.cpu.gprf.mem[16][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][31]$_DFFE_PP_  (.CLK(clknet_leaf_453_clk_in_regs),
    .D(net902),
    .DE(net1371),
    .Q(\inst$top.soc.cpu.gprf.mem[16][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk_in_regs),
    .D(net1059),
    .DE(net1371),
    .Q(\inst$top.soc.cpu.gprf.mem[16][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk_in_regs),
    .D(net1011),
    .DE(net1370),
    .Q(\inst$top.soc.cpu.gprf.mem[16][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk_in_regs),
    .D(net1054),
    .DE(net1371),
    .Q(\inst$top.soc.cpu.gprf.mem[16][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk_in_regs),
    .D(net1049),
    .DE(net1371),
    .Q(\inst$top.soc.cpu.gprf.mem[16][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk_in_regs),
    .D(net892),
    .DE(net1372),
    .Q(\inst$top.soc.cpu.gprf.mem[16][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk_in_regs),
    .D(net1005),
    .DE(net1370),
    .Q(\inst$top.soc.cpu.gprf.mem[16][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_437_clk_in_regs),
    .D(net999),
    .DE(net1370),
    .Q(\inst$top.soc.cpu.gprf.mem[16][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk_in_regs),
    .D(net1065),
    .DE(net1488),
    .Q(\inst$top.soc.cpu.gprf.mem[17][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_408_clk_in_regs),
    .D(net994),
    .DE(net1488),
    .Q(\inst$top.soc.cpu.gprf.mem[17][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_411_clk_in_regs),
    .D(net991),
    .DE(net1488),
    .Q(\inst$top.soc.cpu.gprf.mem[17][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][12]$_DFFE_PP_  (.CLK(clknet_leaf_505_clk_in_regs),
    .D(net985),
    .DE(net1490),
    .Q(\inst$top.soc.cpu.gprf.mem[17][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][13]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk_in_regs),
    .D(net983),
    .DE(net1488),
    .Q(\inst$top.soc.cpu.gprf.mem[17][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][14]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk_in_regs),
    .D(net976),
    .DE(net1491),
    .Q(\inst$top.soc.cpu.gprf.mem[17][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][15]$_DFFE_PP_  (.CLK(clknet_leaf_469_clk_in_regs),
    .D(net887),
    .DE(net1491),
    .Q(\inst$top.soc.cpu.gprf.mem[17][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][16]$_DFFE_PP_  (.CLK(clknet_leaf_506_clk_in_regs),
    .D(net972),
    .DE(net1490),
    .Q(\inst$top.soc.cpu.gprf.mem[17][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][17]$_DFFE_PP_  (.CLK(clknet_leaf_478_clk_in_regs),
    .D(net967),
    .DE(net1491),
    .Q(\inst$top.soc.cpu.gprf.mem[17][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][18]$_DFFE_PP_  (.CLK(clknet_leaf_365_clk_in_regs),
    .D(net963),
    .DE(net1488),
    .Q(\inst$top.soc.cpu.gprf.mem[17][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][19]$_DFFE_PP_  (.CLK(clknet_leaf_470_clk_in_regs),
    .D(net959),
    .DE(net1491),
    .Q(\inst$top.soc.cpu.gprf.mem[17][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk_in_regs),
    .D(net1015),
    .DE(net1488),
    .Q(\inst$top.soc.cpu.gprf.mem[17][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][20]$_DFFE_PP_  (.CLK(clknet_leaf_513_clk_in_regs),
    .D(net956),
    .DE(net1489),
    .Q(\inst$top.soc.cpu.gprf.mem[17][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][21]$_DFFE_PP_  (.CLK(clknet_leaf_450_clk_in_regs),
    .D(net952),
    .DE(net1490),
    .Q(\inst$top.soc.cpu.gprf.mem[17][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][22]$_DFFE_PP_  (.CLK(clknet_leaf_417_clk_in_regs),
    .D(net945),
    .DE(net1488),
    .Q(\inst$top.soc.cpu.gprf.mem[17][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][23]$_DFFE_PP_  (.CLK(clknet_leaf_396_clk_in_regs),
    .D(net942),
    .DE(net1489),
    .Q(\inst$top.soc.cpu.gprf.mem[17][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][24]$_DFFE_PP_  (.CLK(clknet_leaf_503_clk_in_regs),
    .D(net936),
    .DE(net1491),
    .Q(\inst$top.soc.cpu.gprf.mem[17][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][25]$_DFFE_PP_  (.CLK(clknet_leaf_435_clk_in_regs),
    .D(net932),
    .DE(net1489),
    .Q(\inst$top.soc.cpu.gprf.mem[17][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][26]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk_in_regs),
    .D(net926),
    .DE(net1488),
    .Q(\inst$top.soc.cpu.gprf.mem[17][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][27]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk_in_regs),
    .D(net920),
    .DE(net1490),
    .Q(\inst$top.soc.cpu.gprf.mem[17][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][28]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk_in_regs),
    .D(net916),
    .DE(net1491),
    .Q(\inst$top.soc.cpu.gprf.mem[17][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][29]$_DFFE_PP_  (.CLK(clknet_leaf_507_clk_in_regs),
    .D(net913),
    .DE(net1490),
    .Q(\inst$top.soc.cpu.gprf.mem[17][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk_in_regs),
    .D(net1060),
    .DE(net1488),
    .Q(\inst$top.soc.cpu.gprf.mem[17][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][30]$_DFFE_PP_  (.CLK(clknet_leaf_432_clk_in_regs),
    .D(net907),
    .DE(net1489),
    .Q(\inst$top.soc.cpu.gprf.mem[17][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][31]$_DFFE_PP_  (.CLK(clknet_leaf_459_clk_in_regs),
    .D(net902),
    .DE(net1490),
    .Q(\inst$top.soc.cpu.gprf.mem[17][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk_in_regs),
    .D(net1059),
    .DE(net1490),
    .Q(\inst$top.soc.cpu.gprf.mem[17][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk_in_regs),
    .D(net1011),
    .DE(net1488),
    .Q(\inst$top.soc.cpu.gprf.mem[17][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk_in_regs),
    .D(net1054),
    .DE(net1490),
    .Q(\inst$top.soc.cpu.gprf.mem[17][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk_in_regs),
    .D(net1049),
    .DE(net1490),
    .Q(\inst$top.soc.cpu.gprf.mem[17][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk_in_regs),
    .D(net892),
    .DE(net1491),
    .Q(\inst$top.soc.cpu.gprf.mem[17][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk_in_regs),
    .D(net1005),
    .DE(net1489),
    .Q(\inst$top.soc.cpu.gprf.mem[17][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_437_clk_in_regs),
    .D(net999),
    .DE(net1490),
    .Q(\inst$top.soc.cpu.gprf.mem[17][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk_in_regs),
    .D(net1065),
    .DE(net1492),
    .Q(\inst$top.soc.cpu.gprf.mem[18][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_442_clk_in_regs),
    .D(net994),
    .DE(net1492),
    .Q(\inst$top.soc.cpu.gprf.mem[18][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_395_clk_in_regs),
    .D(net991),
    .DE(net1492),
    .Q(\inst$top.soc.cpu.gprf.mem[18][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][12]$_DFFE_PP_  (.CLK(clknet_leaf_505_clk_in_regs),
    .D(net985),
    .DE(net1494),
    .Q(\inst$top.soc.cpu.gprf.mem[18][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][13]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk_in_regs),
    .D(net980),
    .DE(net1492),
    .Q(\inst$top.soc.cpu.gprf.mem[18][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][14]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk_in_regs),
    .D(net976),
    .DE(net1494),
    .Q(\inst$top.soc.cpu.gprf.mem[18][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][15]$_DFFE_PP_  (.CLK(clknet_leaf_469_clk_in_regs),
    .D(net887),
    .DE(net1495),
    .Q(\inst$top.soc.cpu.gprf.mem[18][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][16]$_DFFE_PP_  (.CLK(clknet_leaf_506_clk_in_regs),
    .D(net972),
    .DE(net1494),
    .Q(\inst$top.soc.cpu.gprf.mem[18][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][17]$_DFFE_PP_  (.CLK(clknet_leaf_478_clk_in_regs),
    .D(net967),
    .DE(net1495),
    .Q(\inst$top.soc.cpu.gprf.mem[18][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][18]$_DFFE_PP_  (.CLK(clknet_leaf_365_clk_in_regs),
    .D(net963),
    .DE(net1492),
    .Q(\inst$top.soc.cpu.gprf.mem[18][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][19]$_DFFE_PP_  (.CLK(clknet_leaf_471_clk_in_regs),
    .D(net959),
    .DE(net1495),
    .Q(\inst$top.soc.cpu.gprf.mem[18][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk_in_regs),
    .D(net1015),
    .DE(net1492),
    .Q(\inst$top.soc.cpu.gprf.mem[18][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][20]$_DFFE_PP_  (.CLK(clknet_leaf_513_clk_in_regs),
    .D(net956),
    .DE(net1493),
    .Q(\inst$top.soc.cpu.gprf.mem[18][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][21]$_DFFE_PP_  (.CLK(clknet_leaf_450_clk_in_regs),
    .D(net952),
    .DE(net1494),
    .Q(\inst$top.soc.cpu.gprf.mem[18][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][22]$_DFFE_PP_  (.CLK(clknet_leaf_417_clk_in_regs),
    .D(net946),
    .DE(net1492),
    .Q(\inst$top.soc.cpu.gprf.mem[18][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][23]$_DFFE_PP_  (.CLK(clknet_leaf_397_clk_in_regs),
    .D(net942),
    .DE(net1493),
    .Q(\inst$top.soc.cpu.gprf.mem[18][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][24]$_DFFE_PP_  (.CLK(clknet_leaf_503_clk_in_regs),
    .D(net936),
    .DE(net1495),
    .Q(\inst$top.soc.cpu.gprf.mem[18][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][25]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk_in_regs),
    .D(net929),
    .DE(net1493),
    .Q(\inst$top.soc.cpu.gprf.mem[18][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][26]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk_in_regs),
    .D(net926),
    .DE(net1492),
    .Q(\inst$top.soc.cpu.gprf.mem[18][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][27]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk_in_regs),
    .D(net923),
    .DE(net1494),
    .Q(\inst$top.soc.cpu.gprf.mem[18][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][28]$_DFFE_PP_  (.CLK(clknet_leaf_460_clk_in_regs),
    .D(net916),
    .DE(net1495),
    .Q(\inst$top.soc.cpu.gprf.mem[18][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][29]$_DFFE_PP_  (.CLK(clknet_leaf_507_clk_in_regs),
    .D(net913),
    .DE(net1494),
    .Q(\inst$top.soc.cpu.gprf.mem[18][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk_in_regs),
    .D(net1060),
    .DE(net1492),
    .Q(\inst$top.soc.cpu.gprf.mem[18][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][30]$_DFFE_PP_  (.CLK(clknet_leaf_433_clk_in_regs),
    .D(net907),
    .DE(net1493),
    .Q(\inst$top.soc.cpu.gprf.mem[18][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][31]$_DFFE_PP_  (.CLK(clknet_leaf_456_clk_in_regs),
    .D(net902),
    .DE(net1494),
    .Q(\inst$top.soc.cpu.gprf.mem[18][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk_in_regs),
    .D(net1059),
    .DE(net1495),
    .Q(\inst$top.soc.cpu.gprf.mem[18][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk_in_regs),
    .D(net1011),
    .DE(net1492),
    .Q(\inst$top.soc.cpu.gprf.mem[18][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk_in_regs),
    .D(net1054),
    .DE(net1494),
    .Q(\inst$top.soc.cpu.gprf.mem[18][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk_in_regs),
    .D(net1050),
    .DE(net1494),
    .Q(\inst$top.soc.cpu.gprf.mem[18][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk_in_regs),
    .D(net892),
    .DE(net1495),
    .Q(\inst$top.soc.cpu.gprf.mem[18][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk_in_regs),
    .D(net1005),
    .DE(net1493),
    .Q(\inst$top.soc.cpu.gprf.mem[18][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_437_clk_in_regs),
    .D(net1000),
    .DE(net1494),
    .Q(\inst$top.soc.cpu.gprf.mem[18][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk_in_regs),
    .D(net1067),
    .DE(net1496),
    .Q(\inst$top.soc.cpu.gprf.mem[19][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_407_clk_in_regs),
    .D(net994),
    .DE(net1496),
    .Q(\inst$top.soc.cpu.gprf.mem[19][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_395_clk_in_regs),
    .D(net991),
    .DE(net1496),
    .Q(\inst$top.soc.cpu.gprf.mem[19][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][12]$_DFFE_PP_  (.CLK(clknet_leaf_505_clk_in_regs),
    .D(net986),
    .DE(net1498),
    .Q(\inst$top.soc.cpu.gprf.mem[19][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][13]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk_in_regs),
    .D(net980),
    .DE(net1496),
    .Q(\inst$top.soc.cpu.gprf.mem[19][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][14]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk_in_regs),
    .D(net976),
    .DE(net1499),
    .Q(\inst$top.soc.cpu.gprf.mem[19][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][15]$_DFFE_PP_  (.CLK(clknet_leaf_470_clk_in_regs),
    .D(net887),
    .DE(net1499),
    .Q(\inst$top.soc.cpu.gprf.mem[19][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][16]$_DFFE_PP_  (.CLK(clknet_leaf_506_clk_in_regs),
    .D(net972),
    .DE(net1498),
    .Q(\inst$top.soc.cpu.gprf.mem[19][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][17]$_DFFE_PP_  (.CLK(clknet_leaf_478_clk_in_regs),
    .D(net967),
    .DE(net1499),
    .Q(\inst$top.soc.cpu.gprf.mem[19][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][18]$_DFFE_PP_  (.CLK(clknet_leaf_366_clk_in_regs),
    .D(net963),
    .DE(net1496),
    .Q(\inst$top.soc.cpu.gprf.mem[19][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][19]$_DFFE_PP_  (.CLK(clknet_leaf_470_clk_in_regs),
    .D(net959),
    .DE(net1499),
    .Q(\inst$top.soc.cpu.gprf.mem[19][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk_in_regs),
    .D(net1015),
    .DE(net1496),
    .Q(\inst$top.soc.cpu.gprf.mem[19][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][20]$_DFFE_PP_  (.CLK(clknet_leaf_513_clk_in_regs),
    .D(net954),
    .DE(net1496),
    .Q(\inst$top.soc.cpu.gprf.mem[19][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][21]$_DFFE_PP_  (.CLK(clknet_leaf_489_clk_in_regs),
    .D(net952),
    .DE(net1498),
    .Q(\inst$top.soc.cpu.gprf.mem[19][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][22]$_DFFE_PP_  (.CLK(clknet_leaf_417_clk_in_regs),
    .D(net946),
    .DE(net1496),
    .Q(\inst$top.soc.cpu.gprf.mem[19][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][23]$_DFFE_PP_  (.CLK(clknet_leaf_397_clk_in_regs),
    .D(net942),
    .DE(net1497),
    .Q(\inst$top.soc.cpu.gprf.mem[19][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][24]$_DFFE_PP_  (.CLK(clknet_leaf_504_clk_in_regs),
    .D(net936),
    .DE(net1499),
    .Q(\inst$top.soc.cpu.gprf.mem[19][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][25]$_DFFE_PP_  (.CLK(clknet_leaf_434_clk_in_regs),
    .D(net932),
    .DE(net1497),
    .Q(\inst$top.soc.cpu.gprf.mem[19][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][26]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk_in_regs),
    .D(net927),
    .DE(net1496),
    .Q(\inst$top.soc.cpu.gprf.mem[19][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][27]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk_in_regs),
    .D(net923),
    .DE(net1498),
    .Q(\inst$top.soc.cpu.gprf.mem[19][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][28]$_DFFE_PP_  (.CLK(clknet_leaf_466_clk_in_regs),
    .D(net916),
    .DE(net1499),
    .Q(\inst$top.soc.cpu.gprf.mem[19][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][29]$_DFFE_PP_  (.CLK(clknet_leaf_507_clk_in_regs),
    .D(net913),
    .DE(net1498),
    .Q(\inst$top.soc.cpu.gprf.mem[19][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk_in_regs),
    .D(net1060),
    .DE(net1496),
    .Q(\inst$top.soc.cpu.gprf.mem[19][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][30]$_DFFE_PP_  (.CLK(clknet_leaf_430_clk_in_regs),
    .D(net906),
    .DE(net1497),
    .Q(\inst$top.soc.cpu.gprf.mem[19][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][31]$_DFFE_PP_  (.CLK(clknet_leaf_456_clk_in_regs),
    .D(net901),
    .DE(net1498),
    .Q(\inst$top.soc.cpu.gprf.mem[19][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk_in_regs),
    .D(net1059),
    .DE(net1498),
    .Q(\inst$top.soc.cpu.gprf.mem[19][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk_in_regs),
    .D(net1012),
    .DE(net1497),
    .Q(\inst$top.soc.cpu.gprf.mem[19][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk_in_regs),
    .D(net1054),
    .DE(net1498),
    .Q(\inst$top.soc.cpu.gprf.mem[19][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk_in_regs),
    .D(net1050),
    .DE(net1498),
    .Q(\inst$top.soc.cpu.gprf.mem[19][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk_in_regs),
    .D(net893),
    .DE(net1499),
    .Q(\inst$top.soc.cpu.gprf.mem[19][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk_in_regs),
    .D(net1005),
    .DE(net1497),
    .Q(\inst$top.soc.cpu.gprf.mem[19][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_457_clk_in_regs),
    .D(net1000),
    .DE(net1498),
    .Q(\inst$top.soc.cpu.gprf.mem[19][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk_in_regs),
    .D(net1064),
    .DE(net1578),
    .Q(\inst$top.soc.cpu.gprf.mem[1][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_439_clk_in_regs),
    .D(net995),
    .DE(net1577),
    .Q(\inst$top.soc.cpu.gprf.mem[1][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_412_clk_in_regs),
    .D(net992),
    .DE(net1578),
    .Q(\inst$top.soc.cpu.gprf.mem[1][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_500_clk_in_regs),
    .D(net986),
    .DE(net1576),
    .Q(\inst$top.soc.cpu.gprf.mem[1][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][13]$_DFFE_PP_  (.CLK(clknet_6_50__leaf_clk_in_regs),
    .D(net980),
    .DE(net1577),
    .Q(\inst$top.soc.cpu.gprf.mem[1][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk_in_regs),
    .D(net978),
    .DE(net1576),
    .Q(\inst$top.soc.cpu.gprf.mem[1][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_467_clk_in_regs),
    .D(net889),
    .DE(net1576),
    .Q(\inst$top.soc.cpu.gprf.mem[1][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_494_clk_in_regs),
    .D(net973),
    .DE(net1576),
    .Q(\inst$top.soc.cpu.gprf.mem[1][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_476_clk_in_regs),
    .D(net970),
    .DE(net1576),
    .Q(\inst$top.soc.cpu.gprf.mem[1][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_364_clk_in_regs),
    .D(net965),
    .DE(net1578),
    .Q(\inst$top.soc.cpu.gprf.mem[1][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_466_clk_in_regs),
    .D(net961),
    .DE(net1576),
    .Q(\inst$top.soc.cpu.gprf.mem[1][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk_in_regs),
    .D(net1017),
    .DE(net1578),
    .Q(\inst$top.soc.cpu.gprf.mem[1][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_511_clk_in_regs),
    .D(net954),
    .DE(net1577),
    .Q(\inst$top.soc.cpu.gprf.mem[1][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_463_clk_in_regs),
    .D(net949),
    .DE(net1579),
    .Q(\inst$top.soc.cpu.gprf.mem[1][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_416_clk_in_regs),
    .D(net944),
    .DE(net1578),
    .Q(\inst$top.soc.cpu.gprf.mem[1][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_398_clk_in_regs),
    .D(net940),
    .DE(net1577),
    .Q(\inst$top.soc.cpu.gprf.mem[1][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_499_clk_in_regs),
    .D(net935),
    .DE(net1579),
    .Q(\inst$top.soc.cpu.gprf.mem[1][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk_in_regs),
    .D(net929),
    .DE(net1577),
    .Q(\inst$top.soc.cpu.gprf.mem[1][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk_in_regs),
    .D(net928),
    .DE(net1578),
    .Q(\inst$top.soc.cpu.gprf.mem[1][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk_in_regs),
    .D(net920),
    .DE(net1576),
    .Q(\inst$top.soc.cpu.gprf.mem[1][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk_in_regs),
    .D(net918),
    .DE(net1576),
    .Q(\inst$top.soc.cpu.gprf.mem[1][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_510_clk_in_regs),
    .D(net911),
    .DE(net1577),
    .Q(\inst$top.soc.cpu.gprf.mem[1][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk_in_regs),
    .D(net1062),
    .DE(net1578),
    .Q(\inst$top.soc.cpu.gprf.mem[1][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_430_clk_in_regs),
    .D(net906),
    .DE(net1578),
    .Q(\inst$top.soc.cpu.gprf.mem[1][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_448_clk_in_regs),
    .D(net901),
    .DE(net1577),
    .Q(\inst$top.soc.cpu.gprf.mem[1][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk_in_regs),
    .D(net1056),
    .DE(net1576),
    .Q(\inst$top.soc.cpu.gprf.mem[1][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk_in_regs),
    .D(net1010),
    .DE(net1578),
    .Q(\inst$top.soc.cpu.gprf.mem[1][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk_in_regs),
    .D(net1053),
    .DE(net1577),
    .Q(\inst$top.soc.cpu.gprf.mem[1][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk_in_regs),
    .D(net1048),
    .DE(net1577),
    .Q(\inst$top.soc.cpu.gprf.mem[1][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk_in_regs),
    .D(net890),
    .DE(net1576),
    .Q(\inst$top.soc.cpu.gprf.mem[1][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk_in_regs),
    .D(net1005),
    .DE(net1578),
    .Q(\inst$top.soc.cpu.gprf.mem[1][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_436_clk_in_regs),
    .D(net999),
    .DE(net1577),
    .Q(\inst$top.soc.cpu.gprf.mem[1][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk_in_regs),
    .D(net1066),
    .DE(net1500),
    .Q(\inst$top.soc.cpu.gprf.mem[20][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_441_clk_in_regs),
    .D(net994),
    .DE(net1500),
    .Q(\inst$top.soc.cpu.gprf.mem[20][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_394_clk_in_regs),
    .D(net992),
    .DE(net1500),
    .Q(\inst$top.soc.cpu.gprf.mem[20][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][12]$_DFFE_PP_  (.CLK(clknet_leaf_504_clk_in_regs),
    .D(net985),
    .DE(net1502),
    .Q(\inst$top.soc.cpu.gprf.mem[20][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][13]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk_in_regs),
    .D(net982),
    .DE(net1500),
    .Q(\inst$top.soc.cpu.gprf.mem[20][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][14]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk_in_regs),
    .D(net976),
    .DE(net1502),
    .Q(\inst$top.soc.cpu.gprf.mem[20][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][15]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk_in_regs),
    .D(net888),
    .DE(net1502),
    .Q(\inst$top.soc.cpu.gprf.mem[20][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][16]$_DFFE_PP_  (.CLK(clknet_leaf_506_clk_in_regs),
    .D(net971),
    .DE(net1502),
    .Q(\inst$top.soc.cpu.gprf.mem[20][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][17]$_DFFE_PP_  (.CLK(clknet_leaf_481_clk_in_regs),
    .D(net969),
    .DE(net1503),
    .Q(\inst$top.soc.cpu.gprf.mem[20][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][18]$_DFFE_PP_  (.CLK(clknet_leaf_363_clk_in_regs),
    .D(net963),
    .DE(net1500),
    .Q(\inst$top.soc.cpu.gprf.mem[20][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][19]$_DFFE_PP_  (.CLK(clknet_leaf_472_clk_in_regs),
    .D(net960),
    .DE(net1503),
    .Q(\inst$top.soc.cpu.gprf.mem[20][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk_in_regs),
    .D(net1015),
    .DE(net1500),
    .Q(\inst$top.soc.cpu.gprf.mem[20][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][20]$_DFFE_PP_  (.CLK(clknet_leaf_512_clk_in_regs),
    .D(net954),
    .DE(net1501),
    .Q(\inst$top.soc.cpu.gprf.mem[20][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][21]$_DFFE_PP_  (.CLK(clknet_leaf_489_clk_in_regs),
    .D(net949),
    .DE(net1502),
    .Q(\inst$top.soc.cpu.gprf.mem[20][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][22]$_DFFE_PP_  (.CLK(clknet_leaf_419_clk_in_regs),
    .D(net946),
    .DE(net1500),
    .Q(\inst$top.soc.cpu.gprf.mem[20][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][23]$_DFFE_PP_  (.CLK(clknet_leaf_397_clk_in_regs),
    .D(net940),
    .DE(net1501),
    .Q(\inst$top.soc.cpu.gprf.mem[20][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][24]$_DFFE_PP_  (.CLK(clknet_leaf_503_clk_in_regs),
    .D(net936),
    .DE(net1503),
    .Q(\inst$top.soc.cpu.gprf.mem[20][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][25]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk_in_regs),
    .D(net931),
    .DE(net1501),
    .Q(\inst$top.soc.cpu.gprf.mem[20][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][26]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk_in_regs),
    .D(net926),
    .DE(net1500),
    .Q(\inst$top.soc.cpu.gprf.mem[20][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][27]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk_in_regs),
    .D(net924),
    .DE(net1502),
    .Q(\inst$top.soc.cpu.gprf.mem[20][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][28]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk_in_regs),
    .D(net916),
    .DE(net1503),
    .Q(\inst$top.soc.cpu.gprf.mem[20][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][29]$_DFFE_PP_  (.CLK(clknet_leaf_512_clk_in_regs),
    .D(net915),
    .DE(net1502),
    .Q(\inst$top.soc.cpu.gprf.mem[20][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk_in_regs),
    .D(net1061),
    .DE(net1500),
    .Q(\inst$top.soc.cpu.gprf.mem[20][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][30]$_DFFE_PP_  (.CLK(clknet_leaf_432_clk_in_regs),
    .D(net908),
    .DE(net1501),
    .Q(\inst$top.soc.cpu.gprf.mem[20][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][31]$_DFFE_PP_  (.CLK(clknet_leaf_455_clk_in_regs),
    .D(net901),
    .DE(net1502),
    .Q(\inst$top.soc.cpu.gprf.mem[20][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk_in_regs),
    .D(net1059),
    .DE(net1503),
    .Q(\inst$top.soc.cpu.gprf.mem[20][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk_in_regs),
    .D(net1012),
    .DE(net1500),
    .Q(\inst$top.soc.cpu.gprf.mem[20][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk_in_regs),
    .D(net1054),
    .DE(net1502),
    .Q(\inst$top.soc.cpu.gprf.mem[20][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk_in_regs),
    .D(net1050),
    .DE(net1501),
    .Q(\inst$top.soc.cpu.gprf.mem[20][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk_in_regs),
    .D(net893),
    .DE(net1503),
    .Q(\inst$top.soc.cpu.gprf.mem[20][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk_in_regs),
    .D(net1007),
    .DE(net1501),
    .Q(\inst$top.soc.cpu.gprf.mem[20][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_456_clk_in_regs),
    .D(net1001),
    .DE(net1502),
    .Q(\inst$top.soc.cpu.gprf.mem[20][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk_in_regs),
    .D(net1066),
    .DE(net1504),
    .Q(\inst$top.soc.cpu.gprf.mem[21][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_441_clk_in_regs),
    .D(net994),
    .DE(net1504),
    .Q(\inst$top.soc.cpu.gprf.mem[21][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_394_clk_in_regs),
    .D(net992),
    .DE(net1504),
    .Q(\inst$top.soc.cpu.gprf.mem[21][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][12]$_DFFE_PP_  (.CLK(clknet_leaf_504_clk_in_regs),
    .D(net985),
    .DE(net1506),
    .Q(\inst$top.soc.cpu.gprf.mem[21][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][13]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk_in_regs),
    .D(net982),
    .DE(net1504),
    .Q(\inst$top.soc.cpu.gprf.mem[21][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][14]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk_in_regs),
    .D(net976),
    .DE(net1506),
    .Q(\inst$top.soc.cpu.gprf.mem[21][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][15]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk_in_regs),
    .D(net888),
    .DE(net1506),
    .Q(\inst$top.soc.cpu.gprf.mem[21][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][16]$_DFFE_PP_  (.CLK(clknet_leaf_508_clk_in_regs),
    .D(net971),
    .DE(net1506),
    .Q(\inst$top.soc.cpu.gprf.mem[21][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][17]$_DFFE_PP_  (.CLK(clknet_leaf_479_clk_in_regs),
    .D(net969),
    .DE(net1507),
    .Q(\inst$top.soc.cpu.gprf.mem[21][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][18]$_DFFE_PP_  (.CLK(clknet_leaf_363_clk_in_regs),
    .D(net963),
    .DE(net1504),
    .Q(\inst$top.soc.cpu.gprf.mem[21][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][19]$_DFFE_PP_  (.CLK(clknet_leaf_472_clk_in_regs),
    .D(net960),
    .DE(net1507),
    .Q(\inst$top.soc.cpu.gprf.mem[21][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk_in_regs),
    .D(net1015),
    .DE(net1504),
    .Q(\inst$top.soc.cpu.gprf.mem[21][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][20]$_DFFE_PP_  (.CLK(clknet_leaf_511_clk_in_regs),
    .D(net954),
    .DE(net1505),
    .Q(\inst$top.soc.cpu.gprf.mem[21][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][21]$_DFFE_PP_  (.CLK(clknet_leaf_489_clk_in_regs),
    .D(net952),
    .DE(net1506),
    .Q(\inst$top.soc.cpu.gprf.mem[21][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][22]$_DFFE_PP_  (.CLK(clknet_leaf_419_clk_in_regs),
    .D(net946),
    .DE(net1504),
    .Q(\inst$top.soc.cpu.gprf.mem[21][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][23]$_DFFE_PP_  (.CLK(clknet_leaf_397_clk_in_regs),
    .D(net940),
    .DE(net1505),
    .Q(\inst$top.soc.cpu.gprf.mem[21][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][24]$_DFFE_PP_  (.CLK(clknet_leaf_503_clk_in_regs),
    .D(net936),
    .DE(net1507),
    .Q(\inst$top.soc.cpu.gprf.mem[21][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][25]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk_in_regs),
    .D(net930),
    .DE(net1505),
    .Q(\inst$top.soc.cpu.gprf.mem[21][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][26]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk_in_regs),
    .D(net926),
    .DE(net1504),
    .Q(\inst$top.soc.cpu.gprf.mem[21][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][27]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk_in_regs),
    .D(net924),
    .DE(net1506),
    .Q(\inst$top.soc.cpu.gprf.mem[21][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][28]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk_in_regs),
    .D(net916),
    .DE(net1507),
    .Q(\inst$top.soc.cpu.gprf.mem[21][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][29]$_DFFE_PP_  (.CLK(clknet_leaf_512_clk_in_regs),
    .D(net915),
    .DE(net1506),
    .Q(\inst$top.soc.cpu.gprf.mem[21][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk_in_regs),
    .D(net1061),
    .DE(net1504),
    .Q(\inst$top.soc.cpu.gprf.mem[21][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][30]$_DFFE_PP_  (.CLK(clknet_leaf_432_clk_in_regs),
    .D(net908),
    .DE(net1505),
    .Q(\inst$top.soc.cpu.gprf.mem[21][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][31]$_DFFE_PP_  (.CLK(clknet_leaf_455_clk_in_regs),
    .D(net901),
    .DE(net1506),
    .Q(\inst$top.soc.cpu.gprf.mem[21][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk_in_regs),
    .D(net1059),
    .DE(net1507),
    .Q(\inst$top.soc.cpu.gprf.mem[21][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk_in_regs),
    .D(net1012),
    .DE(net1504),
    .Q(\inst$top.soc.cpu.gprf.mem[21][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk_in_regs),
    .D(net1054),
    .DE(net1506),
    .Q(\inst$top.soc.cpu.gprf.mem[21][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk_in_regs),
    .D(net1050),
    .DE(net1505),
    .Q(\inst$top.soc.cpu.gprf.mem[21][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk_in_regs),
    .D(net893),
    .DE(net1507),
    .Q(\inst$top.soc.cpu.gprf.mem[21][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk_in_regs),
    .D(net1005),
    .DE(net1505),
    .Q(\inst$top.soc.cpu.gprf.mem[21][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_457_clk_in_regs),
    .D(net1001),
    .DE(net1506),
    .Q(\inst$top.soc.cpu.gprf.mem[21][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk_in_regs),
    .D(net1066),
    .DE(net1508),
    .Q(\inst$top.soc.cpu.gprf.mem[22][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_441_clk_in_regs),
    .D(net994),
    .DE(net1508),
    .Q(\inst$top.soc.cpu.gprf.mem[22][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_394_clk_in_regs),
    .D(net991),
    .DE(net1508),
    .Q(\inst$top.soc.cpu.gprf.mem[22][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][12]$_DFFE_PP_  (.CLK(clknet_leaf_504_clk_in_regs),
    .D(net985),
    .DE(net1510),
    .Q(\inst$top.soc.cpu.gprf.mem[22][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][13]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk_in_regs),
    .D(net982),
    .DE(net1508),
    .Q(\inst$top.soc.cpu.gprf.mem[22][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][14]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk_in_regs),
    .D(net977),
    .DE(net1510),
    .Q(\inst$top.soc.cpu.gprf.mem[22][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][15]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk_in_regs),
    .D(net888),
    .DE(net1511),
    .Q(\inst$top.soc.cpu.gprf.mem[22][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][16]$_DFFE_PP_  (.CLK(clknet_leaf_508_clk_in_regs),
    .D(net971),
    .DE(net1510),
    .Q(\inst$top.soc.cpu.gprf.mem[22][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][17]$_DFFE_PP_  (.CLK(clknet_leaf_481_clk_in_regs),
    .D(net969),
    .DE(net1511),
    .Q(\inst$top.soc.cpu.gprf.mem[22][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][18]$_DFFE_PP_  (.CLK(clknet_leaf_363_clk_in_regs),
    .D(net963),
    .DE(net1508),
    .Q(\inst$top.soc.cpu.gprf.mem[22][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][19]$_DFFE_PP_  (.CLK(clknet_leaf_473_clk_in_regs),
    .D(net960),
    .DE(net1511),
    .Q(\inst$top.soc.cpu.gprf.mem[22][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk_in_regs),
    .D(net1016),
    .DE(net1508),
    .Q(\inst$top.soc.cpu.gprf.mem[22][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][20]$_DFFE_PP_  (.CLK(clknet_leaf_511_clk_in_regs),
    .D(net954),
    .DE(net1509),
    .Q(\inst$top.soc.cpu.gprf.mem[22][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][21]$_DFFE_PP_  (.CLK(clknet_leaf_489_clk_in_regs),
    .D(net952),
    .DE(net1510),
    .Q(\inst$top.soc.cpu.gprf.mem[22][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][22]$_DFFE_PP_  (.CLK(clknet_leaf_419_clk_in_regs),
    .D(net946),
    .DE(net1508),
    .Q(\inst$top.soc.cpu.gprf.mem[22][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][23]$_DFFE_PP_  (.CLK(clknet_leaf_397_clk_in_regs),
    .D(net940),
    .DE(net1509),
    .Q(\inst$top.soc.cpu.gprf.mem[22][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][24]$_DFFE_PP_  (.CLK(clknet_leaf_503_clk_in_regs),
    .D(net936),
    .DE(net1511),
    .Q(\inst$top.soc.cpu.gprf.mem[22][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][25]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk_in_regs),
    .D(net930),
    .DE(net1509),
    .Q(\inst$top.soc.cpu.gprf.mem[22][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][26]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk_in_regs),
    .D(net926),
    .DE(net1508),
    .Q(\inst$top.soc.cpu.gprf.mem[22][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][27]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk_in_regs),
    .D(net923),
    .DE(net1510),
    .Q(\inst$top.soc.cpu.gprf.mem[22][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][28]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk_in_regs),
    .D(net916),
    .DE(net1511),
    .Q(\inst$top.soc.cpu.gprf.mem[22][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][29]$_DFFE_PP_  (.CLK(clknet_leaf_512_clk_in_regs),
    .D(net913),
    .DE(net1510),
    .Q(\inst$top.soc.cpu.gprf.mem[22][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk_in_regs),
    .D(net1061),
    .DE(net1508),
    .Q(\inst$top.soc.cpu.gprf.mem[22][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][30]$_DFFE_PP_  (.CLK(clknet_leaf_431_clk_in_regs),
    .D(net907),
    .DE(net1509),
    .Q(\inst$top.soc.cpu.gprf.mem[22][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][31]$_DFFE_PP_  (.CLK(clknet_leaf_453_clk_in_regs),
    .D(net902),
    .DE(net1510),
    .Q(\inst$top.soc.cpu.gprf.mem[22][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk_in_regs),
    .D(net1059),
    .DE(net1511),
    .Q(\inst$top.soc.cpu.gprf.mem[22][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk_in_regs),
    .D(net1012),
    .DE(net1508),
    .Q(\inst$top.soc.cpu.gprf.mem[22][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk_in_regs),
    .D(net1054),
    .DE(net1510),
    .Q(\inst$top.soc.cpu.gprf.mem[22][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk_in_regs),
    .D(net1050),
    .DE(net1510),
    .Q(\inst$top.soc.cpu.gprf.mem[22][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk_in_regs),
    .D(net893),
    .DE(net1511),
    .Q(\inst$top.soc.cpu.gprf.mem[22][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk_in_regs),
    .D(net1007),
    .DE(net1509),
    .Q(\inst$top.soc.cpu.gprf.mem[22][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_457_clk_in_regs),
    .D(net1000),
    .DE(net1510),
    .Q(\inst$top.soc.cpu.gprf.mem[22][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk_in_regs),
    .D(net1066),
    .DE(net1512),
    .Q(\inst$top.soc.cpu.gprf.mem[23][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_441_clk_in_regs),
    .D(net994),
    .DE(net1512),
    .Q(\inst$top.soc.cpu.gprf.mem[23][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_394_clk_in_regs),
    .D(net992),
    .DE(net1512),
    .Q(\inst$top.soc.cpu.gprf.mem[23][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][12]$_DFFE_PP_  (.CLK(clknet_leaf_504_clk_in_regs),
    .D(net987),
    .DE(net1514),
    .Q(\inst$top.soc.cpu.gprf.mem[23][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][13]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk_in_regs),
    .D(net982),
    .DE(net1512),
    .Q(\inst$top.soc.cpu.gprf.mem[23][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][14]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk_in_regs),
    .D(net977),
    .DE(net1514),
    .Q(\inst$top.soc.cpu.gprf.mem[23][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][15]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk_in_regs),
    .D(net888),
    .DE(net1515),
    .Q(\inst$top.soc.cpu.gprf.mem[23][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][16]$_DFFE_PP_  (.CLK(clknet_leaf_506_clk_in_regs),
    .D(net971),
    .DE(net1514),
    .Q(\inst$top.soc.cpu.gprf.mem[23][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][17]$_DFFE_PP_  (.CLK(clknet_leaf_481_clk_in_regs),
    .D(net969),
    .DE(net1515),
    .Q(\inst$top.soc.cpu.gprf.mem[23][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][18]$_DFFE_PP_  (.CLK(clknet_leaf_364_clk_in_regs),
    .D(net966),
    .DE(net1512),
    .Q(\inst$top.soc.cpu.gprf.mem[23][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][19]$_DFFE_PP_  (.CLK(clknet_leaf_472_clk_in_regs),
    .D(net960),
    .DE(net1515),
    .Q(\inst$top.soc.cpu.gprf.mem[23][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk_in_regs),
    .D(net1016),
    .DE(net1512),
    .Q(\inst$top.soc.cpu.gprf.mem[23][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][20]$_DFFE_PP_  (.CLK(clknet_leaf_512_clk_in_regs),
    .D(net954),
    .DE(net1513),
    .Q(\inst$top.soc.cpu.gprf.mem[23][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][21]$_DFFE_PP_  (.CLK(clknet_leaf_489_clk_in_regs),
    .D(net949),
    .DE(net1514),
    .Q(\inst$top.soc.cpu.gprf.mem[23][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][22]$_DFFE_PP_  (.CLK(clknet_leaf_419_clk_in_regs),
    .D(net946),
    .DE(net1512),
    .Q(\inst$top.soc.cpu.gprf.mem[23][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][23]$_DFFE_PP_  (.CLK(clknet_6_55__leaf_clk_in_regs),
    .D(net940),
    .DE(net1513),
    .Q(\inst$top.soc.cpu.gprf.mem[23][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][24]$_DFFE_PP_  (.CLK(clknet_leaf_503_clk_in_regs),
    .D(net937),
    .DE(net1515),
    .Q(\inst$top.soc.cpu.gprf.mem[23][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][25]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk_in_regs),
    .D(net930),
    .DE(net1513),
    .Q(\inst$top.soc.cpu.gprf.mem[23][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][26]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk_in_regs),
    .D(net926),
    .DE(net1512),
    .Q(\inst$top.soc.cpu.gprf.mem[23][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][27]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk_in_regs),
    .D(net924),
    .DE(net1514),
    .Q(\inst$top.soc.cpu.gprf.mem[23][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][28]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk_in_regs),
    .D(net916),
    .DE(net1515),
    .Q(\inst$top.soc.cpu.gprf.mem[23][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][29]$_DFFE_PP_  (.CLK(clknet_leaf_507_clk_in_regs),
    .D(net913),
    .DE(net1514),
    .Q(\inst$top.soc.cpu.gprf.mem[23][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk_in_regs),
    .D(net1061),
    .DE(net1512),
    .Q(\inst$top.soc.cpu.gprf.mem[23][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][30]$_DFFE_PP_  (.CLK(clknet_leaf_431_clk_in_regs),
    .D(net907),
    .DE(net1513),
    .Q(\inst$top.soc.cpu.gprf.mem[23][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][31]$_DFFE_PP_  (.CLK(clknet_leaf_456_clk_in_regs),
    .D(net902),
    .DE(net1514),
    .Q(\inst$top.soc.cpu.gprf.mem[23][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk_in_regs),
    .D(net1059),
    .DE(net1515),
    .Q(\inst$top.soc.cpu.gprf.mem[23][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk_in_regs),
    .D(net1012),
    .DE(net1512),
    .Q(\inst$top.soc.cpu.gprf.mem[23][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk_in_regs),
    .D(net1054),
    .DE(net1514),
    .Q(\inst$top.soc.cpu.gprf.mem[23][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk_in_regs),
    .D(net1050),
    .DE(net1514),
    .Q(\inst$top.soc.cpu.gprf.mem[23][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk_in_regs),
    .D(net893),
    .DE(net1515),
    .Q(\inst$top.soc.cpu.gprf.mem[23][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk_in_regs),
    .D(net1007),
    .DE(net1513),
    .Q(\inst$top.soc.cpu.gprf.mem[23][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_457_clk_in_regs),
    .D(net1000),
    .DE(net1514),
    .Q(\inst$top.soc.cpu.gprf.mem[23][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk_in_regs),
    .D(net1067),
    .DE(net1516),
    .Q(\inst$top.soc.cpu.gprf.mem[24][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_438_clk_in_regs),
    .D(net995),
    .DE(net1518),
    .Q(\inst$top.soc.cpu.gprf.mem[24][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_418_clk_in_regs),
    .D(net989),
    .DE(net1516),
    .Q(\inst$top.soc.cpu.gprf.mem[24][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][12]$_DFFE_PP_  (.CLK(clknet_leaf_485_clk_in_regs),
    .D(net984),
    .DE(net1517),
    .Q(\inst$top.soc.cpu.gprf.mem[24][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][13]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk_in_regs),
    .D(net980),
    .DE(net1516),
    .Q(\inst$top.soc.cpu.gprf.mem[24][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][14]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk_in_regs),
    .D(net978),
    .DE(net1517),
    .Q(\inst$top.soc.cpu.gprf.mem[24][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][15]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk_in_regs),
    .D(net885),
    .DE(net1517),
    .Q(\inst$top.soc.cpu.gprf.mem[24][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][16]$_DFFE_PP_  (.CLK(clknet_leaf_492_clk_in_regs),
    .D(net971),
    .DE(net1518),
    .Q(\inst$top.soc.cpu.gprf.mem[24][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][17]$_DFFE_PP_  (.CLK(clknet_leaf_476_clk_in_regs),
    .D(net968),
    .DE(net1517),
    .Q(\inst$top.soc.cpu.gprf.mem[24][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][18]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk_in_regs),
    .D(net965),
    .DE(net1516),
    .Q(\inst$top.soc.cpu.gprf.mem[24][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][19]$_DFFE_PP_  (.CLK(clknet_leaf_468_clk_in_regs),
    .D(net958),
    .DE(net1517),
    .Q(\inst$top.soc.cpu.gprf.mem[24][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk_in_regs),
    .D(net1014),
    .DE(net1516),
    .Q(\inst$top.soc.cpu.gprf.mem[24][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][20]$_DFFE_PP_  (.CLK(clknet_leaf_446_clk_in_regs),
    .D(net953),
    .DE(net1518),
    .Q(\inst$top.soc.cpu.gprf.mem[24][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][21]$_DFFE_PP_  (.CLK(clknet_leaf_464_clk_in_regs),
    .D(net950),
    .DE(net1517),
    .Q(\inst$top.soc.cpu.gprf.mem[24][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][22]$_DFFE_PP_  (.CLK(clknet_leaf_421_clk_in_regs),
    .D(net944),
    .DE(net1516),
    .Q(\inst$top.soc.cpu.gprf.mem[24][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][23]$_DFFE_PP_  (.CLK(clknet_leaf_407_clk_in_regs),
    .D(net939),
    .DE(net1516),
    .Q(\inst$top.soc.cpu.gprf.mem[24][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][24]$_DFFE_PP_  (.CLK(clknet_leaf_490_clk_in_regs),
    .D(net934),
    .DE(net1518),
    .Q(\inst$top.soc.cpu.gprf.mem[24][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][25]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk_in_regs),
    .D(net929),
    .DE(net1519),
    .Q(\inst$top.soc.cpu.gprf.mem[24][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][26]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk_in_regs),
    .D(net927),
    .DE(net1516),
    .Q(\inst$top.soc.cpu.gprf.mem[24][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][27]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk_in_regs),
    .D(net921),
    .DE(net1517),
    .Q(\inst$top.soc.cpu.gprf.mem[24][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][28]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk_in_regs),
    .D(net917),
    .DE(net1517),
    .Q(\inst$top.soc.cpu.gprf.mem[24][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][29]$_DFFE_PP_  (.CLK(clknet_leaf_447_clk_in_regs),
    .D(net911),
    .DE(net1518),
    .Q(\inst$top.soc.cpu.gprf.mem[24][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk_in_regs),
    .D(net1061),
    .DE(net1516),
    .Q(\inst$top.soc.cpu.gprf.mem[24][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][30]$_DFFE_PP_  (.CLK(clknet_leaf_428_clk_in_regs),
    .D(net909),
    .DE(net1519),
    .Q(\inst$top.soc.cpu.gprf.mem[24][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][31]$_DFFE_PP_  (.CLK(clknet_leaf_462_clk_in_regs),
    .D(net902),
    .DE(net1518),
    .Q(\inst$top.soc.cpu.gprf.mem[24][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk_in_regs),
    .D(net1057),
    .DE(net1517),
    .Q(\inst$top.soc.cpu.gprf.mem[24][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk_in_regs),
    .D(net1009),
    .DE(net1516),
    .Q(\inst$top.soc.cpu.gprf.mem[24][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk_in_regs),
    .D(net1052),
    .DE(net1518),
    .Q(\inst$top.soc.cpu.gprf.mem[24][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk_in_regs),
    .D(net1049),
    .DE(net1518),
    .Q(\inst$top.soc.cpu.gprf.mem[24][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk_in_regs),
    .D(net890),
    .DE(net1517),
    .Q(\inst$top.soc.cpu.gprf.mem[24][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk_in_regs),
    .D(net1007),
    .DE(net1519),
    .Q(\inst$top.soc.cpu.gprf.mem[24][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk_in_regs),
    .D(net1000),
    .DE(net1518),
    .Q(\inst$top.soc.cpu.gprf.mem[24][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk_in_regs),
    .D(net1067),
    .DE(net1520),
    .Q(\inst$top.soc.cpu.gprf.mem[25][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_438_clk_in_regs),
    .D(net995),
    .DE(net1522),
    .Q(\inst$top.soc.cpu.gprf.mem[25][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_418_clk_in_regs),
    .D(net989),
    .DE(net1520),
    .Q(\inst$top.soc.cpu.gprf.mem[25][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][12]$_DFFE_PP_  (.CLK(clknet_leaf_485_clk_in_regs),
    .D(net984),
    .DE(net1521),
    .Q(\inst$top.soc.cpu.gprf.mem[25][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][13]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk_in_regs),
    .D(net980),
    .DE(net1520),
    .Q(\inst$top.soc.cpu.gprf.mem[25][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][14]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk_in_regs),
    .D(net978),
    .DE(net1521),
    .Q(\inst$top.soc.cpu.gprf.mem[25][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][15]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk_in_regs),
    .D(net885),
    .DE(net1521),
    .Q(\inst$top.soc.cpu.gprf.mem[25][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][16]$_DFFE_PP_  (.CLK(clknet_leaf_492_clk_in_regs),
    .D(net971),
    .DE(net1522),
    .Q(\inst$top.soc.cpu.gprf.mem[25][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][17]$_DFFE_PP_  (.CLK(clknet_leaf_476_clk_in_regs),
    .D(net968),
    .DE(net1521),
    .Q(\inst$top.soc.cpu.gprf.mem[25][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][18]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk_in_regs),
    .D(net965),
    .DE(net1520),
    .Q(\inst$top.soc.cpu.gprf.mem[25][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][19]$_DFFE_PP_  (.CLK(clknet_leaf_474_clk_in_regs),
    .D(net958),
    .DE(net1521),
    .Q(\inst$top.soc.cpu.gprf.mem[25][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk_in_regs),
    .D(net1014),
    .DE(net1520),
    .Q(\inst$top.soc.cpu.gprf.mem[25][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][20]$_DFFE_PP_  (.CLK(clknet_leaf_446_clk_in_regs),
    .D(net953),
    .DE(net1522),
    .Q(\inst$top.soc.cpu.gprf.mem[25][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][21]$_DFFE_PP_  (.CLK(clknet_leaf_464_clk_in_regs),
    .D(net950),
    .DE(net1521),
    .Q(\inst$top.soc.cpu.gprf.mem[25][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][22]$_DFFE_PP_  (.CLK(clknet_leaf_421_clk_in_regs),
    .D(net944),
    .DE(net1520),
    .Q(\inst$top.soc.cpu.gprf.mem[25][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][23]$_DFFE_PP_  (.CLK(clknet_leaf_407_clk_in_regs),
    .D(net939),
    .DE(net1520),
    .Q(\inst$top.soc.cpu.gprf.mem[25][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][24]$_DFFE_PP_  (.CLK(clknet_leaf_490_clk_in_regs),
    .D(net934),
    .DE(net1522),
    .Q(\inst$top.soc.cpu.gprf.mem[25][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][25]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk_in_regs),
    .D(net929),
    .DE(net1523),
    .Q(\inst$top.soc.cpu.gprf.mem[25][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][26]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk_in_regs),
    .D(net927),
    .DE(net1520),
    .Q(\inst$top.soc.cpu.gprf.mem[25][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][27]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk_in_regs),
    .D(net921),
    .DE(net1521),
    .Q(\inst$top.soc.cpu.gprf.mem[25][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][28]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk_in_regs),
    .D(net916),
    .DE(net1521),
    .Q(\inst$top.soc.cpu.gprf.mem[25][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][29]$_DFFE_PP_  (.CLK(clknet_leaf_447_clk_in_regs),
    .D(net911),
    .DE(net1522),
    .Q(\inst$top.soc.cpu.gprf.mem[25][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk_in_regs),
    .D(net1061),
    .DE(net1520),
    .Q(\inst$top.soc.cpu.gprf.mem[25][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][30]$_DFFE_PP_  (.CLK(clknet_leaf_427_clk_in_regs),
    .D(net909),
    .DE(net1523),
    .Q(\inst$top.soc.cpu.gprf.mem[25][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][31]$_DFFE_PP_  (.CLK(clknet_leaf_461_clk_in_regs),
    .D(net902),
    .DE(net1522),
    .Q(\inst$top.soc.cpu.gprf.mem[25][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk_in_regs),
    .D(net1057),
    .DE(net1521),
    .Q(\inst$top.soc.cpu.gprf.mem[25][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk_in_regs),
    .D(net1009),
    .DE(net1520),
    .Q(\inst$top.soc.cpu.gprf.mem[25][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk_in_regs),
    .D(net1052),
    .DE(net1522),
    .Q(\inst$top.soc.cpu.gprf.mem[25][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk_in_regs),
    .D(net1049),
    .DE(net1522),
    .Q(\inst$top.soc.cpu.gprf.mem[25][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk_in_regs),
    .D(net890),
    .DE(net1521),
    .Q(\inst$top.soc.cpu.gprf.mem[25][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk_in_regs),
    .D(net1007),
    .DE(net1523),
    .Q(\inst$top.soc.cpu.gprf.mem[25][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk_in_regs),
    .D(net1000),
    .DE(net1522),
    .Q(\inst$top.soc.cpu.gprf.mem[25][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk_in_regs),
    .D(net1067),
    .DE(net1524),
    .Q(\inst$top.soc.cpu.gprf.mem[26][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_440_clk_in_regs),
    .D(net995),
    .DE(net1526),
    .Q(\inst$top.soc.cpu.gprf.mem[26][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_418_clk_in_regs),
    .D(net989),
    .DE(net1524),
    .Q(\inst$top.soc.cpu.gprf.mem[26][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][12]$_DFFE_PP_  (.CLK(clknet_leaf_484_clk_in_regs),
    .D(net984),
    .DE(net1525),
    .Q(\inst$top.soc.cpu.gprf.mem[26][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][13]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk_in_regs),
    .D(net981),
    .DE(net1524),
    .Q(\inst$top.soc.cpu.gprf.mem[26][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][14]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk_in_regs),
    .D(net978),
    .DE(net1525),
    .Q(\inst$top.soc.cpu.gprf.mem[26][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][15]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk_in_regs),
    .D(net885),
    .DE(net1525),
    .Q(\inst$top.soc.cpu.gprf.mem[26][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][16]$_DFFE_PP_  (.CLK(clknet_leaf_492_clk_in_regs),
    .D(net971),
    .DE(net1526),
    .Q(\inst$top.soc.cpu.gprf.mem[26][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][17]$_DFFE_PP_  (.CLK(clknet_leaf_477_clk_in_regs),
    .D(net968),
    .DE(net1525),
    .Q(\inst$top.soc.cpu.gprf.mem[26][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][18]$_DFFE_PP_  (.CLK(clknet_leaf_425_clk_in_regs),
    .D(net964),
    .DE(net1524),
    .Q(\inst$top.soc.cpu.gprf.mem[26][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][19]$_DFFE_PP_  (.CLK(clknet_leaf_468_clk_in_regs),
    .D(net958),
    .DE(net1525),
    .Q(\inst$top.soc.cpu.gprf.mem[26][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk_in_regs),
    .D(net1014),
    .DE(net1524),
    .Q(\inst$top.soc.cpu.gprf.mem[26][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][20]$_DFFE_PP_  (.CLK(clknet_leaf_445_clk_in_regs),
    .D(net955),
    .DE(net1526),
    .Q(\inst$top.soc.cpu.gprf.mem[26][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][21]$_DFFE_PP_  (.CLK(clknet_leaf_475_clk_in_regs),
    .D(net950),
    .DE(net1525),
    .Q(\inst$top.soc.cpu.gprf.mem[26][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][22]$_DFFE_PP_  (.CLK(clknet_leaf_421_clk_in_regs),
    .D(net947),
    .DE(net1524),
    .Q(\inst$top.soc.cpu.gprf.mem[26][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][23]$_DFFE_PP_  (.CLK(clknet_leaf_406_clk_in_regs),
    .D(net939),
    .DE(net1524),
    .Q(\inst$top.soc.cpu.gprf.mem[26][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][24]$_DFFE_PP_  (.CLK(clknet_leaf_484_clk_in_regs),
    .D(net935),
    .DE(net1526),
    .Q(\inst$top.soc.cpu.gprf.mem[26][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][25]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk_in_regs),
    .D(net929),
    .DE(net1527),
    .Q(\inst$top.soc.cpu.gprf.mem[26][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][26]$_DFFE_PP_  (.CLK(clknet_leaf_426_clk_in_regs),
    .D(net927),
    .DE(net1524),
    .Q(\inst$top.soc.cpu.gprf.mem[26][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][27]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk_in_regs),
    .D(net921),
    .DE(net1525),
    .Q(\inst$top.soc.cpu.gprf.mem[26][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][28]$_DFFE_PP_  (.CLK(clknet_leaf_460_clk_in_regs),
    .D(net917),
    .DE(net1525),
    .Q(\inst$top.soc.cpu.gprf.mem[26][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][29]$_DFFE_PP_  (.CLK(clknet_leaf_447_clk_in_regs),
    .D(net912),
    .DE(net1526),
    .Q(\inst$top.soc.cpu.gprf.mem[26][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk_in_regs),
    .D(net1061),
    .DE(net1524),
    .Q(\inst$top.soc.cpu.gprf.mem[26][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][30]$_DFFE_PP_  (.CLK(clknet_leaf_428_clk_in_regs),
    .D(net907),
    .DE(net1527),
    .Q(\inst$top.soc.cpu.gprf.mem[26][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][31]$_DFFE_PP_  (.CLK(clknet_leaf_461_clk_in_regs),
    .D(net902),
    .DE(net1526),
    .Q(\inst$top.soc.cpu.gprf.mem[26][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk_in_regs),
    .D(net1057),
    .DE(net1525),
    .Q(\inst$top.soc.cpu.gprf.mem[26][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk_in_regs),
    .D(net1009),
    .DE(net1524),
    .Q(\inst$top.soc.cpu.gprf.mem[26][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk_in_regs),
    .D(net1052),
    .DE(net1526),
    .Q(\inst$top.soc.cpu.gprf.mem[26][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk_in_regs),
    .D(net1048),
    .DE(net1526),
    .Q(\inst$top.soc.cpu.gprf.mem[26][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk_in_regs),
    .D(net891),
    .DE(net1525),
    .Q(\inst$top.soc.cpu.gprf.mem[26][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk_in_regs),
    .D(net1007),
    .DE(net1527),
    .Q(\inst$top.soc.cpu.gprf.mem[26][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk_in_regs),
    .D(net1000),
    .DE(net1526),
    .Q(\inst$top.soc.cpu.gprf.mem[26][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk_in_regs),
    .D(net1067),
    .DE(net1528),
    .Q(\inst$top.soc.cpu.gprf.mem[27][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_440_clk_in_regs),
    .D(net995),
    .DE(net1530),
    .Q(\inst$top.soc.cpu.gprf.mem[27][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_409_clk_in_regs),
    .D(net989),
    .DE(net1528),
    .Q(\inst$top.soc.cpu.gprf.mem[27][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][12]$_DFFE_PP_  (.CLK(clknet_leaf_484_clk_in_regs),
    .D(net984),
    .DE(net1529),
    .Q(\inst$top.soc.cpu.gprf.mem[27][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][13]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk_in_regs),
    .D(net981),
    .DE(net1528),
    .Q(\inst$top.soc.cpu.gprf.mem[27][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][14]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk_in_regs),
    .D(net978),
    .DE(net1529),
    .Q(\inst$top.soc.cpu.gprf.mem[27][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][15]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk_in_regs),
    .D(net885),
    .DE(net1529),
    .Q(\inst$top.soc.cpu.gprf.mem[27][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][16]$_DFFE_PP_  (.CLK(clknet_leaf_492_clk_in_regs),
    .D(net971),
    .DE(net1530),
    .Q(\inst$top.soc.cpu.gprf.mem[27][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][17]$_DFFE_PP_  (.CLK(clknet_leaf_477_clk_in_regs),
    .D(net968),
    .DE(net1529),
    .Q(\inst$top.soc.cpu.gprf.mem[27][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][18]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk_in_regs),
    .D(net964),
    .DE(net1528),
    .Q(\inst$top.soc.cpu.gprf.mem[27][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][19]$_DFFE_PP_  (.CLK(clknet_leaf_474_clk_in_regs),
    .D(net958),
    .DE(net1529),
    .Q(\inst$top.soc.cpu.gprf.mem[27][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk_in_regs),
    .D(net1014),
    .DE(net1528),
    .Q(\inst$top.soc.cpu.gprf.mem[27][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][20]$_DFFE_PP_  (.CLK(clknet_leaf_445_clk_in_regs),
    .D(net955),
    .DE(net1530),
    .Q(\inst$top.soc.cpu.gprf.mem[27][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][21]$_DFFE_PP_  (.CLK(clknet_leaf_475_clk_in_regs),
    .D(net950),
    .DE(net1529),
    .Q(\inst$top.soc.cpu.gprf.mem[27][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][22]$_DFFE_PP_  (.CLK(clknet_leaf_421_clk_in_regs),
    .D(net947),
    .DE(net1528),
    .Q(\inst$top.soc.cpu.gprf.mem[27][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][23]$_DFFE_PP_  (.CLK(clknet_leaf_407_clk_in_regs),
    .D(net939),
    .DE(net1528),
    .Q(\inst$top.soc.cpu.gprf.mem[27][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][24]$_DFFE_PP_  (.CLK(clknet_leaf_485_clk_in_regs),
    .D(net934),
    .DE(net1530),
    .Q(\inst$top.soc.cpu.gprf.mem[27][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][25]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk_in_regs),
    .D(net929),
    .DE(net1528),
    .Q(\inst$top.soc.cpu.gprf.mem[27][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][26]$_DFFE_PP_  (.CLK(clknet_leaf_426_clk_in_regs),
    .D(net927),
    .DE(net1531),
    .Q(\inst$top.soc.cpu.gprf.mem[27][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][27]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk_in_regs),
    .D(net922),
    .DE(net1529),
    .Q(\inst$top.soc.cpu.gprf.mem[27][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][28]$_DFFE_PP_  (.CLK(clknet_leaf_461_clk_in_regs),
    .D(net919),
    .DE(net1529),
    .Q(\inst$top.soc.cpu.gprf.mem[27][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][29]$_DFFE_PP_  (.CLK(clknet_leaf_446_clk_in_regs),
    .D(net912),
    .DE(net1530),
    .Q(\inst$top.soc.cpu.gprf.mem[27][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk_in_regs),
    .D(net1063),
    .DE(net1528),
    .Q(\inst$top.soc.cpu.gprf.mem[27][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][30]$_DFFE_PP_  (.CLK(clknet_leaf_428_clk_in_regs),
    .D(net909),
    .DE(net1531),
    .Q(\inst$top.soc.cpu.gprf.mem[27][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][31]$_DFFE_PP_  (.CLK(clknet_leaf_453_clk_in_regs),
    .D(net902),
    .DE(net1530),
    .Q(\inst$top.soc.cpu.gprf.mem[27][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk_in_regs),
    .D(net1057),
    .DE(net1529),
    .Q(\inst$top.soc.cpu.gprf.mem[27][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk_in_regs),
    .D(net1009),
    .DE(net1528),
    .Q(\inst$top.soc.cpu.gprf.mem[27][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk_in_regs),
    .D(net1055),
    .DE(net1530),
    .Q(\inst$top.soc.cpu.gprf.mem[27][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk_in_regs),
    .D(net1050),
    .DE(net1530),
    .Q(\inst$top.soc.cpu.gprf.mem[27][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk_in_regs),
    .D(net892),
    .DE(net1529),
    .Q(\inst$top.soc.cpu.gprf.mem[27][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk_in_regs),
    .D(net1007),
    .DE(net1531),
    .Q(\inst$top.soc.cpu.gprf.mem[27][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk_in_regs),
    .D(net1000),
    .DE(net1530),
    .Q(\inst$top.soc.cpu.gprf.mem[27][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk_in_regs),
    .D(net1067),
    .DE(net1532),
    .Q(\inst$top.soc.cpu.gprf.mem[28][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_440_clk_in_regs),
    .D(net994),
    .DE(net1534),
    .Q(\inst$top.soc.cpu.gprf.mem[28][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_431_clk_in_regs),
    .D(net990),
    .DE(net1532),
    .Q(\inst$top.soc.cpu.gprf.mem[28][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][12]$_DFFE_PP_  (.CLK(clknet_leaf_483_clk_in_regs),
    .D(net987),
    .DE(net1533),
    .Q(\inst$top.soc.cpu.gprf.mem[28][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][13]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk_in_regs),
    .D(net982),
    .DE(net1534),
    .Q(\inst$top.soc.cpu.gprf.mem[28][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][14]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk_in_regs),
    .D(net975),
    .DE(net1533),
    .Q(\inst$top.soc.cpu.gprf.mem[28][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][15]$_DFFE_PP_  (.CLK(clknet_leaf_467_clk_in_regs),
    .D(net885),
    .DE(net1533),
    .Q(\inst$top.soc.cpu.gprf.mem[28][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][16]$_DFFE_PP_  (.CLK(clknet_leaf_491_clk_in_regs),
    .D(net973),
    .DE(net1533),
    .Q(\inst$top.soc.cpu.gprf.mem[28][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][17]$_DFFE_PP_  (.CLK(clknet_leaf_483_clk_in_regs),
    .D(net968),
    .DE(net1533),
    .Q(\inst$top.soc.cpu.gprf.mem[28][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][18]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk_in_regs),
    .D(net963),
    .DE(net1532),
    .Q(\inst$top.soc.cpu.gprf.mem[28][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][19]$_DFFE_PP_  (.CLK(clknet_leaf_475_clk_in_regs),
    .D(net958),
    .DE(net1533),
    .Q(\inst$top.soc.cpu.gprf.mem[28][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk_in_regs),
    .D(net1014),
    .DE(net1532),
    .Q(\inst$top.soc.cpu.gprf.mem[28][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][20]$_DFFE_PP_  (.CLK(clknet_leaf_404_clk_in_regs),
    .D(net956),
    .DE(net1534),
    .Q(\inst$top.soc.cpu.gprf.mem[28][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][21]$_DFFE_PP_  (.CLK(clknet_leaf_463_clk_in_regs),
    .D(net950),
    .DE(net1533),
    .Q(\inst$top.soc.cpu.gprf.mem[28][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][22]$_DFFE_PP_  (.CLK(clknet_leaf_421_clk_in_regs),
    .D(net945),
    .DE(net1532),
    .Q(\inst$top.soc.cpu.gprf.mem[28][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][23]$_DFFE_PP_  (.CLK(clknet_leaf_407_clk_in_regs),
    .D(net939),
    .DE(net1534),
    .Q(\inst$top.soc.cpu.gprf.mem[28][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][24]$_DFFE_PP_  (.CLK(clknet_leaf_490_clk_in_regs),
    .D(net934),
    .DE(net1535),
    .Q(\inst$top.soc.cpu.gprf.mem[28][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][25]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk_in_regs),
    .D(net929),
    .DE(net1532),
    .Q(\inst$top.soc.cpu.gprf.mem[28][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][26]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk_in_regs),
    .D(net927),
    .DE(net1532),
    .Q(\inst$top.soc.cpu.gprf.mem[28][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][27]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk_in_regs),
    .D(net922),
    .DE(net1533),
    .Q(\inst$top.soc.cpu.gprf.mem[28][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][28]$_DFFE_PP_  (.CLK(clknet_leaf_460_clk_in_regs),
    .D(net919),
    .DE(net1535),
    .Q(\inst$top.soc.cpu.gprf.mem[28][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][29]$_DFFE_PP_  (.CLK(clknet_leaf_446_clk_in_regs),
    .D(net915),
    .DE(net1534),
    .Q(\inst$top.soc.cpu.gprf.mem[28][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk_in_regs),
    .D(net1062),
    .DE(net1532),
    .Q(\inst$top.soc.cpu.gprf.mem[28][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][30]$_DFFE_PP_  (.CLK(clknet_leaf_427_clk_in_regs),
    .D(net906),
    .DE(net1532),
    .Q(\inst$top.soc.cpu.gprf.mem[28][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][31]$_DFFE_PP_  (.CLK(clknet_leaf_452_clk_in_regs),
    .D(net903),
    .DE(net1534),
    .Q(\inst$top.soc.cpu.gprf.mem[28][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk_in_regs),
    .D(net1059),
    .DE(net1533),
    .Q(\inst$top.soc.cpu.gprf.mem[28][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk_in_regs),
    .D(net1009),
    .DE(net1532),
    .Q(\inst$top.soc.cpu.gprf.mem[28][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk_in_regs),
    .D(net1054),
    .DE(net1534),
    .Q(\inst$top.soc.cpu.gprf.mem[28][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk_in_regs),
    .D(net1051),
    .DE(net1534),
    .Q(\inst$top.soc.cpu.gprf.mem[28][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk_in_regs),
    .D(net891),
    .DE(net1533),
    .Q(\inst$top.soc.cpu.gprf.mem[28][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk_in_regs),
    .D(net1008),
    .DE(net1535),
    .Q(\inst$top.soc.cpu.gprf.mem[28][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_437_clk_in_regs),
    .D(net999),
    .DE(net1534),
    .Q(\inst$top.soc.cpu.gprf.mem[28][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk_in_regs),
    .D(net1067),
    .DE(net1536),
    .Q(\inst$top.soc.cpu.gprf.mem[29][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_440_clk_in_regs),
    .D(net994),
    .DE(net1538),
    .Q(\inst$top.soc.cpu.gprf.mem[29][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_409_clk_in_regs),
    .D(net990),
    .DE(net1536),
    .Q(\inst$top.soc.cpu.gprf.mem[29][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][12]$_DFFE_PP_  (.CLK(clknet_leaf_483_clk_in_regs),
    .D(net984),
    .DE(net1537),
    .Q(\inst$top.soc.cpu.gprf.mem[29][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][13]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk_in_regs),
    .D(net982),
    .DE(net1536),
    .Q(\inst$top.soc.cpu.gprf.mem[29][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][14]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk_in_regs),
    .D(net975),
    .DE(net1537),
    .Q(\inst$top.soc.cpu.gprf.mem[29][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][15]$_DFFE_PP_  (.CLK(clknet_leaf_468_clk_in_regs),
    .D(net885),
    .DE(net1537),
    .Q(\inst$top.soc.cpu.gprf.mem[29][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][16]$_DFFE_PP_  (.CLK(clknet_leaf_491_clk_in_regs),
    .D(net973),
    .DE(net1537),
    .Q(\inst$top.soc.cpu.gprf.mem[29][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][17]$_DFFE_PP_  (.CLK(clknet_leaf_480_clk_in_regs),
    .D(net968),
    .DE(net1537),
    .Q(\inst$top.soc.cpu.gprf.mem[29][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][18]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk_in_regs),
    .D(net963),
    .DE(net1536),
    .Q(\inst$top.soc.cpu.gprf.mem[29][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][19]$_DFFE_PP_  (.CLK(clknet_leaf_474_clk_in_regs),
    .D(net958),
    .DE(net1537),
    .Q(\inst$top.soc.cpu.gprf.mem[29][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk_in_regs),
    .D(net1017),
    .DE(net1536),
    .Q(\inst$top.soc.cpu.gprf.mem[29][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][20]$_DFFE_PP_  (.CLK(clknet_leaf_404_clk_in_regs),
    .D(net953),
    .DE(net1538),
    .Q(\inst$top.soc.cpu.gprf.mem[29][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][21]$_DFFE_PP_  (.CLK(clknet_leaf_463_clk_in_regs),
    .D(net950),
    .DE(net1537),
    .Q(\inst$top.soc.cpu.gprf.mem[29][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][22]$_DFFE_PP_  (.CLK(clknet_leaf_421_clk_in_regs),
    .D(net945),
    .DE(net1536),
    .Q(\inst$top.soc.cpu.gprf.mem[29][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][23]$_DFFE_PP_  (.CLK(clknet_leaf_407_clk_in_regs),
    .D(net939),
    .DE(net1536),
    .Q(\inst$top.soc.cpu.gprf.mem[29][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][24]$_DFFE_PP_  (.CLK(clknet_leaf_490_clk_in_regs),
    .D(net934),
    .DE(net1538),
    .Q(\inst$top.soc.cpu.gprf.mem[29][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][25]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk_in_regs),
    .D(net929),
    .DE(net1536),
    .Q(\inst$top.soc.cpu.gprf.mem[29][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][26]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk_in_regs),
    .D(net927),
    .DE(net1539),
    .Q(\inst$top.soc.cpu.gprf.mem[29][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][27]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk_in_regs),
    .D(net922),
    .DE(net1537),
    .Q(\inst$top.soc.cpu.gprf.mem[29][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][28]$_DFFE_PP_  (.CLK(clknet_leaf_462_clk_in_regs),
    .D(net919),
    .DE(net1538),
    .Q(\inst$top.soc.cpu.gprf.mem[29][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][29]$_DFFE_PP_  (.CLK(clknet_leaf_446_clk_in_regs),
    .D(net911),
    .DE(net1538),
    .Q(\inst$top.soc.cpu.gprf.mem[29][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk_in_regs),
    .D(net1063),
    .DE(net1536),
    .Q(\inst$top.soc.cpu.gprf.mem[29][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][30]$_DFFE_PP_  (.CLK(clknet_leaf_427_clk_in_regs),
    .D(net906),
    .DE(net1539),
    .Q(\inst$top.soc.cpu.gprf.mem[29][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][31]$_DFFE_PP_  (.CLK(clknet_leaf_452_clk_in_regs),
    .D(net902),
    .DE(net1538),
    .Q(\inst$top.soc.cpu.gprf.mem[29][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk_in_regs),
    .D(net1057),
    .DE(net1537),
    .Q(\inst$top.soc.cpu.gprf.mem[29][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk_in_regs),
    .D(net1013),
    .DE(net1536),
    .Q(\inst$top.soc.cpu.gprf.mem[29][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk_in_regs),
    .D(net1055),
    .DE(net1538),
    .Q(\inst$top.soc.cpu.gprf.mem[29][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk_in_regs),
    .D(net1051),
    .DE(net1538),
    .Q(\inst$top.soc.cpu.gprf.mem[29][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk_in_regs),
    .D(net891),
    .DE(net1537),
    .Q(\inst$top.soc.cpu.gprf.mem[29][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk_in_regs),
    .D(net1004),
    .DE(net1539),
    .Q(\inst$top.soc.cpu.gprf.mem[29][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk_in_regs),
    .D(net1002),
    .DE(net1538),
    .Q(\inst$top.soc.cpu.gprf.mem[29][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk_in_regs),
    .D(net1064),
    .DE(net1593),
    .Q(\inst$top.soc.cpu.gprf.mem[2][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_443_clk_in_regs),
    .D(net995),
    .DE(net1595),
    .Q(\inst$top.soc.cpu.gprf.mem[2][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_412_clk_in_regs),
    .D(net992),
    .DE(net1593),
    .Q(\inst$top.soc.cpu.gprf.mem[2][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_500_clk_in_regs),
    .D(net986),
    .DE(net1594),
    .Q(\inst$top.soc.cpu.gprf.mem[2][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk_in_regs),
    .D(net981),
    .DE(net1595),
    .Q(\inst$top.soc.cpu.gprf.mem[2][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk_in_regs),
    .D(net975),
    .DE(net1594),
    .Q(\inst$top.soc.cpu.gprf.mem[2][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_467_clk_in_regs),
    .D(net885),
    .DE(net1594),
    .Q(\inst$top.soc.cpu.gprf.mem[2][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_494_clk_in_regs),
    .D(net974),
    .DE(net1594),
    .Q(\inst$top.soc.cpu.gprf.mem[2][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_476_clk_in_regs),
    .D(net970),
    .DE(net1594),
    .Q(\inst$top.soc.cpu.gprf.mem[2][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_424_clk_in_regs),
    .D(net965),
    .DE(net1593),
    .Q(\inst$top.soc.cpu.gprf.mem[2][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_465_clk_in_regs),
    .D(net961),
    .DE(net1594),
    .Q(\inst$top.soc.cpu.gprf.mem[2][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk_in_regs),
    .D(net1017),
    .DE(net1593),
    .Q(\inst$top.soc.cpu.gprf.mem[2][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_401_clk_in_regs),
    .D(net954),
    .DE(net1595),
    .Q(\inst$top.soc.cpu.gprf.mem[2][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_462_clk_in_regs),
    .D(net949),
    .DE(net1596),
    .Q(\inst$top.soc.cpu.gprf.mem[2][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_417_clk_in_regs),
    .D(net945),
    .DE(net1593),
    .Q(\inst$top.soc.cpu.gprf.mem[2][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_399_clk_in_regs),
    .D(net942),
    .DE(net1593),
    .Q(\inst$top.soc.cpu.gprf.mem[2][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_496_clk_in_regs),
    .D(net934),
    .DE(net1596),
    .Q(\inst$top.soc.cpu.gprf.mem[2][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk_in_regs),
    .D(net930),
    .DE(net1595),
    .Q(\inst$top.soc.cpu.gprf.mem[2][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk_in_regs),
    .D(net925),
    .DE(net1593),
    .Q(\inst$top.soc.cpu.gprf.mem[2][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk_in_regs),
    .D(net920),
    .DE(net1594),
    .Q(\inst$top.soc.cpu.gprf.mem[2][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk_in_regs),
    .D(net917),
    .DE(net1594),
    .Q(\inst$top.soc.cpu.gprf.mem[2][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_509_clk_in_regs),
    .D(net913),
    .DE(net1595),
    .Q(\inst$top.soc.cpu.gprf.mem[2][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk_in_regs),
    .D(net1062),
    .DE(net1593),
    .Q(\inst$top.soc.cpu.gprf.mem[2][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_429_clk_in_regs),
    .D(net909),
    .DE(net1593),
    .Q(\inst$top.soc.cpu.gprf.mem[2][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_448_clk_in_regs),
    .D(net904),
    .DE(net1595),
    .Q(\inst$top.soc.cpu.gprf.mem[2][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk_in_regs),
    .D(net1056),
    .DE(net1594),
    .Q(\inst$top.soc.cpu.gprf.mem[2][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk_in_regs),
    .D(net1010),
    .DE(net1593),
    .Q(\inst$top.soc.cpu.gprf.mem[2][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk_in_regs),
    .D(net1053),
    .DE(net1595),
    .Q(\inst$top.soc.cpu.gprf.mem[2][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk_in_regs),
    .D(net1051),
    .DE(net1595),
    .Q(\inst$top.soc.cpu.gprf.mem[2][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk_in_regs),
    .D(net890),
    .DE(net1594),
    .Q(\inst$top.soc.cpu.gprf.mem[2][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk_in_regs),
    .D(net1005),
    .DE(net1596),
    .Q(\inst$top.soc.cpu.gprf.mem[2][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_436_clk_in_regs),
    .D(net1002),
    .DE(net1595),
    .Q(\inst$top.soc.cpu.gprf.mem[2][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk_in_regs),
    .D(net1067),
    .DE(net1540),
    .Q(\inst$top.soc.cpu.gprf.mem[30][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_440_clk_in_regs),
    .D(net995),
    .DE(net1542),
    .Q(\inst$top.soc.cpu.gprf.mem[30][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_408_clk_in_regs),
    .D(net990),
    .DE(net1540),
    .Q(\inst$top.soc.cpu.gprf.mem[30][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][12]$_DFFE_PP_  (.CLK(clknet_leaf_483_clk_in_regs),
    .D(net984),
    .DE(net1541),
    .Q(\inst$top.soc.cpu.gprf.mem[30][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][13]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk_in_regs),
    .D(net982),
    .DE(net1540),
    .Q(\inst$top.soc.cpu.gprf.mem[30][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][14]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk_in_regs),
    .D(net975),
    .DE(net1541),
    .Q(\inst$top.soc.cpu.gprf.mem[30][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][15]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk_in_regs),
    .D(net886),
    .DE(net1541),
    .Q(\inst$top.soc.cpu.gprf.mem[30][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][16]$_DFFE_PP_  (.CLK(clknet_leaf_491_clk_in_regs),
    .D(net971),
    .DE(net1542),
    .Q(\inst$top.soc.cpu.gprf.mem[30][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][17]$_DFFE_PP_  (.CLK(clknet_leaf_479_clk_in_regs),
    .D(net968),
    .DE(net1541),
    .Q(\inst$top.soc.cpu.gprf.mem[30][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][18]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk_in_regs),
    .D(net965),
    .DE(net1540),
    .Q(\inst$top.soc.cpu.gprf.mem[30][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][19]$_DFFE_PP_  (.CLK(clknet_leaf_474_clk_in_regs),
    .D(net958),
    .DE(net1541),
    .Q(\inst$top.soc.cpu.gprf.mem[30][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk_in_regs),
    .D(net1017),
    .DE(net1540),
    .Q(\inst$top.soc.cpu.gprf.mem[30][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][20]$_DFFE_PP_  (.CLK(clknet_leaf_404_clk_in_regs),
    .D(net953),
    .DE(net1542),
    .Q(\inst$top.soc.cpu.gprf.mem[30][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][21]$_DFFE_PP_  (.CLK(clknet_leaf_463_clk_in_regs),
    .D(net950),
    .DE(net1541),
    .Q(\inst$top.soc.cpu.gprf.mem[30][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][22]$_DFFE_PP_  (.CLK(clknet_leaf_421_clk_in_regs),
    .D(net945),
    .DE(net1540),
    .Q(\inst$top.soc.cpu.gprf.mem[30][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][23]$_DFFE_PP_  (.CLK(clknet_leaf_407_clk_in_regs),
    .D(net941),
    .DE(net1540),
    .Q(\inst$top.soc.cpu.gprf.mem[30][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][24]$_DFFE_PP_  (.CLK(clknet_leaf_490_clk_in_regs),
    .D(net934),
    .DE(net1541),
    .Q(\inst$top.soc.cpu.gprf.mem[30][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][25]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk_in_regs),
    .D(net929),
    .DE(net1540),
    .Q(\inst$top.soc.cpu.gprf.mem[30][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][26]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk_in_regs),
    .D(net927),
    .DE(net1540),
    .Q(\inst$top.soc.cpu.gprf.mem[30][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][27]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk_in_regs),
    .D(net922),
    .DE(net1541),
    .Q(\inst$top.soc.cpu.gprf.mem[30][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][28]$_DFFE_PP_  (.CLK(clknet_leaf_461_clk_in_regs),
    .D(net917),
    .DE(net1542),
    .Q(\inst$top.soc.cpu.gprf.mem[30][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][29]$_DFFE_PP_  (.CLK(clknet_leaf_446_clk_in_regs),
    .D(net911),
    .DE(net1542),
    .Q(\inst$top.soc.cpu.gprf.mem[30][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk_in_regs),
    .D(net1063),
    .DE(net1540),
    .Q(\inst$top.soc.cpu.gprf.mem[30][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][30]$_DFFE_PP_  (.CLK(clknet_leaf_427_clk_in_regs),
    .D(net906),
    .DE(net1543),
    .Q(\inst$top.soc.cpu.gprf.mem[30][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][31]$_DFFE_PP_  (.CLK(clknet_leaf_453_clk_in_regs),
    .D(net903),
    .DE(net1542),
    .Q(\inst$top.soc.cpu.gprf.mem[30][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk_in_regs),
    .D(net1057),
    .DE(net1541),
    .Q(\inst$top.soc.cpu.gprf.mem[30][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk_in_regs),
    .D(net1009),
    .DE(net1543),
    .Q(\inst$top.soc.cpu.gprf.mem[30][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk_in_regs),
    .D(net1053),
    .DE(net1542),
    .Q(\inst$top.soc.cpu.gprf.mem[30][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk_in_regs),
    .D(net1050),
    .DE(net1542),
    .Q(\inst$top.soc.cpu.gprf.mem[30][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk_in_regs),
    .D(net893),
    .DE(net1541),
    .Q(\inst$top.soc.cpu.gprf.mem[30][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk_in_regs),
    .D(net1004),
    .DE(net1543),
    .Q(\inst$top.soc.cpu.gprf.mem[30][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk_in_regs),
    .D(net1002),
    .DE(net1542),
    .Q(\inst$top.soc.cpu.gprf.mem[30][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk_in_regs),
    .D(net1064),
    .DE(net1544),
    .Q(\inst$top.soc.cpu.gprf.mem[31][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_440_clk_in_regs),
    .D(net997),
    .DE(net1544),
    .Q(\inst$top.soc.cpu.gprf.mem[31][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_418_clk_in_regs),
    .D(net990),
    .DE(net1544),
    .Q(\inst$top.soc.cpu.gprf.mem[31][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][12]$_DFFE_PP_  (.CLK(clknet_leaf_484_clk_in_regs),
    .D(net984),
    .DE(net1545),
    .Q(\inst$top.soc.cpu.gprf.mem[31][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][13]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk_in_regs),
    .D(net982),
    .DE(net1544),
    .Q(\inst$top.soc.cpu.gprf.mem[31][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][14]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk_in_regs),
    .D(net975),
    .DE(net1545),
    .Q(\inst$top.soc.cpu.gprf.mem[31][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][15]$_DFFE_PP_  (.CLK(clknet_leaf_469_clk_in_regs),
    .D(net886),
    .DE(net1545),
    .Q(\inst$top.soc.cpu.gprf.mem[31][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][16]$_DFFE_PP_  (.CLK(clknet_leaf_492_clk_in_regs),
    .D(net971),
    .DE(net1546),
    .Q(\inst$top.soc.cpu.gprf.mem[31][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][17]$_DFFE_PP_  (.CLK(clknet_leaf_483_clk_in_regs),
    .D(net968),
    .DE(net1545),
    .Q(\inst$top.soc.cpu.gprf.mem[31][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][18]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk_in_regs),
    .D(net963),
    .DE(net1544),
    .Q(\inst$top.soc.cpu.gprf.mem[31][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][19]$_DFFE_PP_  (.CLK(clknet_leaf_475_clk_in_regs),
    .D(net958),
    .DE(net1545),
    .Q(\inst$top.soc.cpu.gprf.mem[31][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk_in_regs),
    .D(net1014),
    .DE(net1544),
    .Q(\inst$top.soc.cpu.gprf.mem[31][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][20]$_DFFE_PP_  (.CLK(clknet_leaf_404_clk_in_regs),
    .D(net956),
    .DE(net1546),
    .Q(\inst$top.soc.cpu.gprf.mem[31][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][21]$_DFFE_PP_  (.CLK(clknet_leaf_452_clk_in_regs),
    .D(net949),
    .DE(net1545),
    .Q(\inst$top.soc.cpu.gprf.mem[31][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][22]$_DFFE_PP_  (.CLK(clknet_leaf_417_clk_in_regs),
    .D(net945),
    .DE(net1544),
    .Q(\inst$top.soc.cpu.gprf.mem[31][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][23]$_DFFE_PP_  (.CLK(clknet_leaf_404_clk_in_regs),
    .D(net941),
    .DE(net1544),
    .Q(\inst$top.soc.cpu.gprf.mem[31][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][24]$_DFFE_PP_  (.CLK(clknet_leaf_496_clk_in_regs),
    .D(net934),
    .DE(net1545),
    .Q(\inst$top.soc.cpu.gprf.mem[31][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][25]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk_in_regs),
    .D(net933),
    .DE(net1544),
    .Q(\inst$top.soc.cpu.gprf.mem[31][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][26]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk_in_regs),
    .D(net927),
    .DE(net1547),
    .Q(\inst$top.soc.cpu.gprf.mem[31][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][27]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk_in_regs),
    .D(net922),
    .DE(net1545),
    .Q(\inst$top.soc.cpu.gprf.mem[31][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][28]$_DFFE_PP_  (.CLK(clknet_leaf_462_clk_in_regs),
    .D(net917),
    .DE(net1546),
    .Q(\inst$top.soc.cpu.gprf.mem[31][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][29]$_DFFE_PP_  (.CLK(clknet_leaf_446_clk_in_regs),
    .D(net911),
    .DE(net1546),
    .Q(\inst$top.soc.cpu.gprf.mem[31][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk_in_regs),
    .D(net1062),
    .DE(net1544),
    .Q(\inst$top.soc.cpu.gprf.mem[31][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][30]$_DFFE_PP_  (.CLK(clknet_leaf_426_clk_in_regs),
    .D(net910),
    .DE(net1547),
    .Q(\inst$top.soc.cpu.gprf.mem[31][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][31]$_DFFE_PP_  (.CLK(clknet_leaf_454_clk_in_regs),
    .D(net903),
    .DE(net1546),
    .Q(\inst$top.soc.cpu.gprf.mem[31][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk_in_regs),
    .D(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[3] ),
    .DE(net1545),
    .Q(\inst$top.soc.cpu.gprf.mem[31][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk_in_regs),
    .D(net1013),
    .DE(net1547),
    .Q(\inst$top.soc.cpu.gprf.mem[31][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk_in_regs),
    .D(net1055),
    .DE(net1546),
    .Q(\inst$top.soc.cpu.gprf.mem[31][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk_in_regs),
    .D(net1051),
    .DE(net1546),
    .Q(\inst$top.soc.cpu.gprf.mem[31][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk_in_regs),
    .D(net891),
    .DE(net1545),
    .Q(\inst$top.soc.cpu.gprf.mem[31][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk_in_regs),
    .D(net1007),
    .DE(net1547),
    .Q(\inst$top.soc.cpu.gprf.mem[31][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_457_clk_in_regs),
    .D(net1000),
    .DE(net1546),
    .Q(\inst$top.soc.cpu.gprf.mem[31][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk_in_regs),
    .D(net1064),
    .DE(net1558),
    .Q(\inst$top.soc.cpu.gprf.mem[3][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_442_clk_in_regs),
    .D(net995),
    .DE(net1557),
    .Q(\inst$top.soc.cpu.gprf.mem[3][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_412_clk_in_regs),
    .D(net992),
    .DE(net1558),
    .Q(\inst$top.soc.cpu.gprf.mem[3][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_498_clk_in_regs),
    .D(net986),
    .DE(net1556),
    .Q(\inst$top.soc.cpu.gprf.mem[3][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk_in_regs),
    .D(net981),
    .DE(net1557),
    .Q(\inst$top.soc.cpu.gprf.mem[3][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk_in_regs),
    .D(net978),
    .DE(net1556),
    .Q(\inst$top.soc.cpu.gprf.mem[3][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_467_clk_in_regs),
    .D(net885),
    .DE(net1556),
    .Q(\inst$top.soc.cpu.gprf.mem[3][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_497_clk_in_regs),
    .D(net972),
    .DE(net1556),
    .Q(\inst$top.soc.cpu.gprf.mem[3][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_476_clk_in_regs),
    .D(net970),
    .DE(net1556),
    .Q(\inst$top.soc.cpu.gprf.mem[3][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_424_clk_in_regs),
    .D(net965),
    .DE(net1558),
    .Q(\inst$top.soc.cpu.gprf.mem[3][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_465_clk_in_regs),
    .D(net961),
    .DE(net1556),
    .Q(\inst$top.soc.cpu.gprf.mem[3][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk_in_regs),
    .D(net1017),
    .DE(net1558),
    .Q(\inst$top.soc.cpu.gprf.mem[3][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_511_clk_in_regs),
    .D(net954),
    .DE(net1557),
    .Q(\inst$top.soc.cpu.gprf.mem[3][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_452_clk_in_regs),
    .D(net949),
    .DE(net1559),
    .Q(\inst$top.soc.cpu.gprf.mem[3][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_417_clk_in_regs),
    .D(net945),
    .DE(net1558),
    .Q(\inst$top.soc.cpu.gprf.mem[3][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_397_clk_in_regs),
    .D(net940),
    .DE(net1557),
    .Q(\inst$top.soc.cpu.gprf.mem[3][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_498_clk_in_regs),
    .D(net935),
    .DE(net1559),
    .Q(\inst$top.soc.cpu.gprf.mem[3][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk_in_regs),
    .D(net930),
    .DE(net1557),
    .Q(\inst$top.soc.cpu.gprf.mem[3][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk_in_regs),
    .D(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[26] ),
    .DE(net1558),
    .Q(\inst$top.soc.cpu.gprf.mem[3][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk_in_regs),
    .D(net920),
    .DE(net1556),
    .Q(\inst$top.soc.cpu.gprf.mem[3][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_459_clk_in_regs),
    .D(net918),
    .DE(net1556),
    .Q(\inst$top.soc.cpu.gprf.mem[3][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_510_clk_in_regs),
    .D(net913),
    .DE(net1557),
    .Q(\inst$top.soc.cpu.gprf.mem[3][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk_in_regs),
    .D(net1063),
    .DE(net1558),
    .Q(\inst$top.soc.cpu.gprf.mem[3][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_419_clk_in_regs),
    .D(net906),
    .DE(net1558),
    .Q(\inst$top.soc.cpu.gprf.mem[3][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_448_clk_in_regs),
    .D(net905),
    .DE(net1557),
    .Q(\inst$top.soc.cpu.gprf.mem[3][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk_in_regs),
    .D(net1056),
    .DE(net1556),
    .Q(\inst$top.soc.cpu.gprf.mem[3][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk_in_regs),
    .D(net1010),
    .DE(net1558),
    .Q(\inst$top.soc.cpu.gprf.mem[3][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk_in_regs),
    .D(net1054),
    .DE(net1557),
    .Q(\inst$top.soc.cpu.gprf.mem[3][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk_in_regs),
    .D(net1051),
    .DE(net1557),
    .Q(\inst$top.soc.cpu.gprf.mem[3][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk_in_regs),
    .D(net890),
    .DE(net1556),
    .Q(\inst$top.soc.cpu.gprf.mem[3][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk_in_regs),
    .D(net1006),
    .DE(net1558),
    .Q(\inst$top.soc.cpu.gprf.mem[3][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_435_clk_in_regs),
    .D(net999),
    .DE(net1557),
    .Q(\inst$top.soc.cpu.gprf.mem[3][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk_in_regs),
    .D(net1064),
    .DE(net1486),
    .Q(\inst$top.soc.cpu.gprf.mem[4][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_442_clk_in_regs),
    .D(net995),
    .DE(net1485),
    .Q(\inst$top.soc.cpu.gprf.mem[4][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_411_clk_in_regs),
    .D(net989),
    .DE(net1486),
    .Q(\inst$top.soc.cpu.gprf.mem[4][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_498_clk_in_regs),
    .D(net986),
    .DE(net1484),
    .Q(\inst$top.soc.cpu.gprf.mem[4][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk_in_regs),
    .D(net981),
    .DE(net1485),
    .Q(\inst$top.soc.cpu.gprf.mem[4][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk_in_regs),
    .D(net978),
    .DE(net1484),
    .Q(\inst$top.soc.cpu.gprf.mem[4][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk_in_regs),
    .D(net889),
    .DE(net1484),
    .Q(\inst$top.soc.cpu.gprf.mem[4][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_497_clk_in_regs),
    .D(net972),
    .DE(net1484),
    .Q(\inst$top.soc.cpu.gprf.mem[4][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_486_clk_in_regs),
    .D(net970),
    .DE(net1484),
    .Q(\inst$top.soc.cpu.gprf.mem[4][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_425_clk_in_regs),
    .D(net964),
    .DE(net1486),
    .Q(\inst$top.soc.cpu.gprf.mem[4][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_464_clk_in_regs),
    .D(net961),
    .DE(net1484),
    .Q(\inst$top.soc.cpu.gprf.mem[4][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk_in_regs),
    .D(net1014),
    .DE(net1486),
    .Q(\inst$top.soc.cpu.gprf.mem[4][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_510_clk_in_regs),
    .D(net954),
    .DE(net1485),
    .Q(\inst$top.soc.cpu.gprf.mem[4][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_451_clk_in_regs),
    .D(net952),
    .DE(net1487),
    .Q(\inst$top.soc.cpu.gprf.mem[4][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_415_clk_in_regs),
    .D(net947),
    .DE(net1486),
    .Q(\inst$top.soc.cpu.gprf.mem[4][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_398_clk_in_regs),
    .D(net940),
    .DE(net1485),
    .Q(\inst$top.soc.cpu.gprf.mem[4][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_497_clk_in_regs),
    .D(net934),
    .DE(net1487),
    .Q(\inst$top.soc.cpu.gprf.mem[4][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk_in_regs),
    .D(net930),
    .DE(net1485),
    .Q(\inst$top.soc.cpu.gprf.mem[4][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk_in_regs),
    .D(net925),
    .DE(net1486),
    .Q(\inst$top.soc.cpu.gprf.mem[4][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk_in_regs),
    .D(net920),
    .DE(net1484),
    .Q(\inst$top.soc.cpu.gprf.mem[4][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk_in_regs),
    .D(net918),
    .DE(net1484),
    .Q(\inst$top.soc.cpu.gprf.mem[4][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_509_clk_in_regs),
    .D(net913),
    .DE(net1485),
    .Q(\inst$top.soc.cpu.gprf.mem[4][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk_in_regs),
    .D(net1062),
    .DE(net1486),
    .Q(\inst$top.soc.cpu.gprf.mem[4][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_429_clk_in_regs),
    .D(net906),
    .DE(net1486),
    .Q(\inst$top.soc.cpu.gprf.mem[4][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_449_clk_in_regs),
    .D(net903),
    .DE(net1487),
    .Q(\inst$top.soc.cpu.gprf.mem[4][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk_in_regs),
    .D(net1056),
    .DE(net1484),
    .Q(\inst$top.soc.cpu.gprf.mem[4][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk_in_regs),
    .D(net1009),
    .DE(net1486),
    .Q(\inst$top.soc.cpu.gprf.mem[4][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk_in_regs),
    .D(net1053),
    .DE(net1485),
    .Q(\inst$top.soc.cpu.gprf.mem[4][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk_in_regs),
    .D(net1051),
    .DE(net1485),
    .Q(\inst$top.soc.cpu.gprf.mem[4][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk_in_regs),
    .D(net890),
    .DE(net1484),
    .Q(\inst$top.soc.cpu.gprf.mem[4][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk_in_regs),
    .D(net1004),
    .DE(net1486),
    .Q(\inst$top.soc.cpu.gprf.mem[4][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_435_clk_in_regs),
    .D(net999),
    .DE(net1485),
    .Q(\inst$top.soc.cpu.gprf.mem[4][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk_in_regs),
    .D(net1064),
    .DE(net1375),
    .Q(\inst$top.soc.cpu.gprf.mem[5][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_445_clk_in_regs),
    .D(net996),
    .DE(net1374),
    .Q(\inst$top.soc.cpu.gprf.mem[5][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_410_clk_in_regs),
    .D(net990),
    .DE(net1375),
    .Q(\inst$top.soc.cpu.gprf.mem[5][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_498_clk_in_regs),
    .D(net986),
    .DE(net1373),
    .Q(\inst$top.soc.cpu.gprf.mem[5][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk_in_regs),
    .D(net981),
    .DE(net1374),
    .Q(\inst$top.soc.cpu.gprf.mem[5][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk_in_regs),
    .D(net978),
    .DE(net1373),
    .Q(\inst$top.soc.cpu.gprf.mem[5][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk_in_regs),
    .D(net885),
    .DE(net1373),
    .Q(\inst$top.soc.cpu.gprf.mem[5][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_497_clk_in_regs),
    .D(net972),
    .DE(net1373),
    .Q(\inst$top.soc.cpu.gprf.mem[5][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_486_clk_in_regs),
    .D(net970),
    .DE(net1373),
    .Q(\inst$top.soc.cpu.gprf.mem[5][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_425_clk_in_regs),
    .D(net964),
    .DE(net1375),
    .Q(\inst$top.soc.cpu.gprf.mem[5][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_465_clk_in_regs),
    .D(net961),
    .DE(net1373),
    .Q(\inst$top.soc.cpu.gprf.mem[5][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk_in_regs),
    .D(net1014),
    .DE(net1375),
    .Q(\inst$top.soc.cpu.gprf.mem[5][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_510_clk_in_regs),
    .D(net955),
    .DE(net1374),
    .Q(\inst$top.soc.cpu.gprf.mem[5][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_451_clk_in_regs),
    .D(net949),
    .DE(net1376),
    .Q(\inst$top.soc.cpu.gprf.mem[5][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_414_clk_in_regs),
    .D(net947),
    .DE(net1375),
    .Q(\inst$top.soc.cpu.gprf.mem[5][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_398_clk_in_regs),
    .D(net940),
    .DE(net1374),
    .Q(\inst$top.soc.cpu.gprf.mem[5][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_497_clk_in_regs),
    .D(net934),
    .DE(net1376),
    .Q(\inst$top.soc.cpu.gprf.mem[5][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk_in_regs),
    .D(net930),
    .DE(net1374),
    .Q(\inst$top.soc.cpu.gprf.mem[5][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk_in_regs),
    .D(net925),
    .DE(net1375),
    .Q(\inst$top.soc.cpu.gprf.mem[5][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk_in_regs),
    .D(net920),
    .DE(net1373),
    .Q(\inst$top.soc.cpu.gprf.mem[5][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk_in_regs),
    .D(net918),
    .DE(net1373),
    .Q(\inst$top.soc.cpu.gprf.mem[5][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_508_clk_in_regs),
    .D(net914),
    .DE(net1376),
    .Q(\inst$top.soc.cpu.gprf.mem[5][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk_in_regs),
    .D(net1062),
    .DE(net1375),
    .Q(\inst$top.soc.cpu.gprf.mem[5][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_429_clk_in_regs),
    .D(net906),
    .DE(net1375),
    .Q(\inst$top.soc.cpu.gprf.mem[5][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_449_clk_in_regs),
    .D(net903),
    .DE(net1374),
    .Q(\inst$top.soc.cpu.gprf.mem[5][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk_in_regs),
    .D(net1056),
    .DE(net1373),
    .Q(\inst$top.soc.cpu.gprf.mem[5][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk_in_regs),
    .D(net1009),
    .DE(net1375),
    .Q(\inst$top.soc.cpu.gprf.mem[5][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk_in_regs),
    .D(net1053),
    .DE(net1374),
    .Q(\inst$top.soc.cpu.gprf.mem[5][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk_in_regs),
    .D(net1051),
    .DE(net1374),
    .Q(\inst$top.soc.cpu.gprf.mem[5][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk_in_regs),
    .D(net890),
    .DE(net1373),
    .Q(\inst$top.soc.cpu.gprf.mem[5][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk_in_regs),
    .D(net1004),
    .DE(net1375),
    .Q(\inst$top.soc.cpu.gprf.mem[5][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_434_clk_in_regs),
    .D(net999),
    .DE(net1374),
    .Q(\inst$top.soc.cpu.gprf.mem[5][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk_in_regs),
    .D(net1064),
    .DE(net1550),
    .Q(\inst$top.soc.cpu.gprf.mem[6][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_442_clk_in_regs),
    .D(net997),
    .DE(net1549),
    .Q(\inst$top.soc.cpu.gprf.mem[6][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_411_clk_in_regs),
    .D(net991),
    .DE(net1550),
    .Q(\inst$top.soc.cpu.gprf.mem[6][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_498_clk_in_regs),
    .D(net986),
    .DE(net1548),
    .Q(\inst$top.soc.cpu.gprf.mem[6][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk_in_regs),
    .D(net981),
    .DE(net1549),
    .Q(\inst$top.soc.cpu.gprf.mem[6][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk_in_regs),
    .D(net975),
    .DE(net1548),
    .Q(\inst$top.soc.cpu.gprf.mem[6][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk_in_regs),
    .D(net885),
    .DE(net1548),
    .Q(\inst$top.soc.cpu.gprf.mem[6][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_497_clk_in_regs),
    .D(net974),
    .DE(net1548),
    .Q(\inst$top.soc.cpu.gprf.mem[6][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_486_clk_in_regs),
    .D(net970),
    .DE(net1548),
    .Q(\inst$top.soc.cpu.gprf.mem[6][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_424_clk_in_regs),
    .D(net964),
    .DE(net1550),
    .Q(\inst$top.soc.cpu.gprf.mem[6][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_465_clk_in_regs),
    .D(net958),
    .DE(net1548),
    .Q(\inst$top.soc.cpu.gprf.mem[6][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk_in_regs),
    .D(net1014),
    .DE(net1550),
    .Q(\inst$top.soc.cpu.gprf.mem[6][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_510_clk_in_regs),
    .D(net955),
    .DE(net1549),
    .Q(\inst$top.soc.cpu.gprf.mem[6][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_451_clk_in_regs),
    .D(net951),
    .DE(net1551),
    .Q(\inst$top.soc.cpu.gprf.mem[6][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_415_clk_in_regs),
    .D(net945),
    .DE(net1550),
    .Q(\inst$top.soc.cpu.gprf.mem[6][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_398_clk_in_regs),
    .D(net940),
    .DE(net1549),
    .Q(\inst$top.soc.cpu.gprf.mem[6][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_496_clk_in_regs),
    .D(net935),
    .DE(net1551),
    .Q(\inst$top.soc.cpu.gprf.mem[6][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk_in_regs),
    .D(net930),
    .DE(net1549),
    .Q(\inst$top.soc.cpu.gprf.mem[6][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk_in_regs),
    .D(net925),
    .DE(net1550),
    .Q(\inst$top.soc.cpu.gprf.mem[6][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk_in_regs),
    .D(net920),
    .DE(net1548),
    .Q(\inst$top.soc.cpu.gprf.mem[6][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk_in_regs),
    .D(net918),
    .DE(net1548),
    .Q(\inst$top.soc.cpu.gprf.mem[6][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_509_clk_in_regs),
    .D(net914),
    .DE(net1549),
    .Q(\inst$top.soc.cpu.gprf.mem[6][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk_in_regs),
    .D(net1062),
    .DE(net1550),
    .Q(\inst$top.soc.cpu.gprf.mem[6][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][30]$_DFFE_PP_  (.CLK(clknet_6_54__leaf_clk_in_regs),
    .D(net910),
    .DE(net1550),
    .Q(\inst$top.soc.cpu.gprf.mem[6][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_449_clk_in_regs),
    .D(net904),
    .DE(net1549),
    .Q(\inst$top.soc.cpu.gprf.mem[6][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk_in_regs),
    .D(net1056),
    .DE(net1548),
    .Q(\inst$top.soc.cpu.gprf.mem[6][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk_in_regs),
    .D(net1009),
    .DE(net1550),
    .Q(\inst$top.soc.cpu.gprf.mem[6][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk_in_regs),
    .D(net1052),
    .DE(net1549),
    .Q(\inst$top.soc.cpu.gprf.mem[6][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk_in_regs),
    .D(net1048),
    .DE(net1549),
    .Q(\inst$top.soc.cpu.gprf.mem[6][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk_in_regs),
    .D(net890),
    .DE(net1548),
    .Q(\inst$top.soc.cpu.gprf.mem[6][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk_in_regs),
    .D(net1006),
    .DE(net1550),
    .Q(\inst$top.soc.cpu.gprf.mem[6][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_435_clk_in_regs),
    .D(net999),
    .DE(net1549),
    .Q(\inst$top.soc.cpu.gprf.mem[6][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk_in_regs),
    .D(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[0] ),
    .DE(net1570),
    .Q(\inst$top.soc.cpu.gprf.mem[7][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_442_clk_in_regs),
    .D(net996),
    .DE(net1569),
    .Q(\inst$top.soc.cpu.gprf.mem[7][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_411_clk_in_regs),
    .D(net991),
    .DE(net1570),
    .Q(\inst$top.soc.cpu.gprf.mem[7][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_498_clk_in_regs),
    .D(net986),
    .DE(net1568),
    .Q(\inst$top.soc.cpu.gprf.mem[7][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk_in_regs),
    .D(net981),
    .DE(net1569),
    .Q(\inst$top.soc.cpu.gprf.mem[7][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk_in_regs),
    .D(net975),
    .DE(net1568),
    .Q(\inst$top.soc.cpu.gprf.mem[7][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk_in_regs),
    .D(net889),
    .DE(net1568),
    .Q(\inst$top.soc.cpu.gprf.mem[7][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_497_clk_in_regs),
    .D(net974),
    .DE(net1568),
    .Q(\inst$top.soc.cpu.gprf.mem[7][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_486_clk_in_regs),
    .D(net970),
    .DE(net1568),
    .Q(\inst$top.soc.cpu.gprf.mem[7][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_423_clk_in_regs),
    .D(net964),
    .DE(net1570),
    .Q(\inst$top.soc.cpu.gprf.mem[7][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_465_clk_in_regs),
    .D(net958),
    .DE(net1568),
    .Q(\inst$top.soc.cpu.gprf.mem[7][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk_in_regs),
    .D(net1014),
    .DE(net1570),
    .Q(\inst$top.soc.cpu.gprf.mem[7][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_512_clk_in_regs),
    .D(net955),
    .DE(net1569),
    .Q(\inst$top.soc.cpu.gprf.mem[7][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_450_clk_in_regs),
    .D(net952),
    .DE(net1571),
    .Q(\inst$top.soc.cpu.gprf.mem[7][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_415_clk_in_regs),
    .D(net945),
    .DE(net1570),
    .Q(\inst$top.soc.cpu.gprf.mem[7][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_513_clk_in_regs),
    .D(net941),
    .DE(net1569),
    .Q(\inst$top.soc.cpu.gprf.mem[7][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_498_clk_in_regs),
    .D(net935),
    .DE(net1571),
    .Q(\inst$top.soc.cpu.gprf.mem[7][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk_in_regs),
    .D(net930),
    .DE(net1569),
    .Q(\inst$top.soc.cpu.gprf.mem[7][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk_in_regs),
    .D(net928),
    .DE(net1570),
    .Q(\inst$top.soc.cpu.gprf.mem[7][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk_in_regs),
    .D(net920),
    .DE(net1568),
    .Q(\inst$top.soc.cpu.gprf.mem[7][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk_in_regs),
    .D(net918),
    .DE(net1568),
    .Q(\inst$top.soc.cpu.gprf.mem[7][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_509_clk_in_regs),
    .D(net914),
    .DE(net1569),
    .Q(\inst$top.soc.cpu.gprf.mem[7][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk_in_regs),
    .D(net1062),
    .DE(net1570),
    .Q(\inst$top.soc.cpu.gprf.mem[7][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_429_clk_in_regs),
    .D(net906),
    .DE(net1570),
    .Q(\inst$top.soc.cpu.gprf.mem[7][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_449_clk_in_regs),
    .D(net903),
    .DE(net1571),
    .Q(\inst$top.soc.cpu.gprf.mem[7][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk_in_regs),
    .D(net1056),
    .DE(net1568),
    .Q(\inst$top.soc.cpu.gprf.mem[7][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk_in_regs),
    .D(net1009),
    .DE(net1570),
    .Q(\inst$top.soc.cpu.gprf.mem[7][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk_in_regs),
    .D(net1052),
    .DE(net1569),
    .Q(\inst$top.soc.cpu.gprf.mem[7][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk_in_regs),
    .D(net1051),
    .DE(net1569),
    .Q(\inst$top.soc.cpu.gprf.mem[7][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk_in_regs),
    .D(net890),
    .DE(net1568),
    .Q(\inst$top.soc.cpu.gprf.mem[7][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk_in_regs),
    .D(net1006),
    .DE(net1570),
    .Q(\inst$top.soc.cpu.gprf.mem[7][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_435_clk_in_regs),
    .D(net999),
    .DE(net1569),
    .Q(\inst$top.soc.cpu.gprf.mem[7][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk_in_regs),
    .D(net1065),
    .DE(net1584),
    .Q(\inst$top.soc.cpu.gprf.mem[8][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_444_clk_in_regs),
    .D(net996),
    .DE(net1586),
    .Q(\inst$top.soc.cpu.gprf.mem[8][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_406_clk_in_regs),
    .D(net990),
    .DE(net1584),
    .Q(\inst$top.soc.cpu.gprf.mem[8][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][12]$_DFFE_PP_  (.CLK(clknet_leaf_500_clk_in_regs),
    .D(net985),
    .DE(net1585),
    .Q(\inst$top.soc.cpu.gprf.mem[8][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][13]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk_in_regs),
    .D(net980),
    .DE(net1584),
    .Q(\inst$top.soc.cpu.gprf.mem[8][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][14]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk_in_regs),
    .D(net975),
    .DE(net1585),
    .Q(\inst$top.soc.cpu.gprf.mem[8][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][15]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk_in_regs),
    .D(net886),
    .DE(net1585),
    .Q(\inst$top.soc.cpu.gprf.mem[8][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][16]$_DFFE_PP_  (.CLK(clknet_leaf_495_clk_in_regs),
    .D(net973),
    .DE(net1585),
    .Q(\inst$top.soc.cpu.gprf.mem[8][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][17]$_DFFE_PP_  (.CLK(clknet_leaf_477_clk_in_regs),
    .D(net968),
    .DE(net1585),
    .Q(\inst$top.soc.cpu.gprf.mem[8][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][18]$_DFFE_PP_  (.CLK(clknet_leaf_426_clk_in_regs),
    .D(net964),
    .DE(net1584),
    .Q(\inst$top.soc.cpu.gprf.mem[8][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][19]$_DFFE_PP_  (.CLK(clknet_leaf_474_clk_in_regs),
    .D(net960),
    .DE(net1585),
    .Q(\inst$top.soc.cpu.gprf.mem[8][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk_in_regs),
    .D(net1015),
    .DE(net1584),
    .Q(\inst$top.soc.cpu.gprf.mem[8][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][20]$_DFFE_PP_  (.CLK(clknet_leaf_400_clk_in_regs),
    .D(net956),
    .DE(net1584),
    .Q(\inst$top.soc.cpu.gprf.mem[8][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][21]$_DFFE_PP_  (.CLK(clknet_leaf_488_clk_in_regs),
    .D(net950),
    .DE(net1586),
    .Q(\inst$top.soc.cpu.gprf.mem[8][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][22]$_DFFE_PP_  (.CLK(clknet_leaf_366_clk_in_regs),
    .D(net948),
    .DE(net1584),
    .Q(\inst$top.soc.cpu.gprf.mem[8][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][23]$_DFFE_PP_  (.CLK(clknet_leaf_400_clk_in_regs),
    .D(net941),
    .DE(net1584),
    .Q(\inst$top.soc.cpu.gprf.mem[8][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][24]$_DFFE_PP_  (.CLK(clknet_leaf_501_clk_in_regs),
    .D(net936),
    .DE(net1586),
    .Q(\inst$top.soc.cpu.gprf.mem[8][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][25]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk_in_regs),
    .D(net931),
    .DE(net1586),
    .Q(\inst$top.soc.cpu.gprf.mem[8][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][26]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk_in_regs),
    .D(net925),
    .DE(net1584),
    .Q(\inst$top.soc.cpu.gprf.mem[8][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][27]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk_in_regs),
    .D(net921),
    .DE(net1585),
    .Q(\inst$top.soc.cpu.gprf.mem[8][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][28]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk_in_regs),
    .D(net916),
    .DE(net1585),
    .Q(\inst$top.soc.cpu.gprf.mem[8][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][29]$_DFFE_PP_  (.CLK(clknet_leaf_493_clk_in_regs),
    .D(net912),
    .DE(net1586),
    .Q(\inst$top.soc.cpu.gprf.mem[8][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk_in_regs),
    .D(net1061),
    .DE(net1584),
    .Q(\inst$top.soc.cpu.gprf.mem[8][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][30]$_DFFE_PP_  (.CLK(clknet_leaf_434_clk_in_regs),
    .D(net908),
    .DE(net1587),
    .Q(\inst$top.soc.cpu.gprf.mem[8][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][31]$_DFFE_PP_  (.CLK(clknet_leaf_448_clk_in_regs),
    .D(net904),
    .DE(net1586),
    .Q(\inst$top.soc.cpu.gprf.mem[8][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk_in_regs),
    .D(net1056),
    .DE(net1585),
    .Q(\inst$top.soc.cpu.gprf.mem[8][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk_in_regs),
    .D(net1011),
    .DE(net1587),
    .Q(\inst$top.soc.cpu.gprf.mem[8][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk_in_regs),
    .D(net1052),
    .DE(net1586),
    .Q(\inst$top.soc.cpu.gprf.mem[8][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk_in_regs),
    .D(net1049),
    .DE(net1586),
    .Q(\inst$top.soc.cpu.gprf.mem[8][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk_in_regs),
    .D(net891),
    .DE(net1585),
    .Q(\inst$top.soc.cpu.gprf.mem[8][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk_in_regs),
    .D(net1005),
    .DE(net1587),
    .Q(\inst$top.soc.cpu.gprf.mem[8][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk_in_regs),
    .D(net1001),
    .DE(net1586),
    .Q(\inst$top.soc.cpu.gprf.mem[8][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk_in_regs),
    .D(net1065),
    .DE(net1572),
    .Q(\inst$top.soc.cpu.gprf.mem[9][0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_444_clk_in_regs),
    .D(net997),
    .DE(net1574),
    .Q(\inst$top.soc.cpu.gprf.mem[9][10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_408_clk_in_regs),
    .D(net990),
    .DE(net1572),
    .Q(\inst$top.soc.cpu.gprf.mem[9][11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][12]$_DFFE_PP_  (.CLK(clknet_leaf_500_clk_in_regs),
    .D(net985),
    .DE(net1573),
    .Q(\inst$top.soc.cpu.gprf.mem[9][12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][13]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk_in_regs),
    .D(net980),
    .DE(net1572),
    .Q(\inst$top.soc.cpu.gprf.mem[9][13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][14]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk_in_regs),
    .D(net977),
    .DE(net1573),
    .Q(\inst$top.soc.cpu.gprf.mem[9][14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][15]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk_in_regs),
    .D(net886),
    .DE(net1573),
    .Q(\inst$top.soc.cpu.gprf.mem[9][15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][16]$_DFFE_PP_  (.CLK(clknet_leaf_495_clk_in_regs),
    .D(net973),
    .DE(net1573),
    .Q(\inst$top.soc.cpu.gprf.mem[9][16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][17]$_DFFE_PP_  (.CLK(clknet_leaf_477_clk_in_regs),
    .D(net968),
    .DE(net1573),
    .Q(\inst$top.soc.cpu.gprf.mem[9][17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][18]$_DFFE_PP_  (.CLK(clknet_leaf_426_clk_in_regs),
    .D(net966),
    .DE(net1572),
    .Q(\inst$top.soc.cpu.gprf.mem[9][18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][19]$_DFFE_PP_  (.CLK(clknet_leaf_473_clk_in_regs),
    .D(net960),
    .DE(net1573),
    .Q(\inst$top.soc.cpu.gprf.mem[9][19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk_in_regs),
    .D(net1015),
    .DE(net1572),
    .Q(\inst$top.soc.cpu.gprf.mem[9][1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][20]$_DFFE_PP_  (.CLK(clknet_leaf_402_clk_in_regs),
    .D(net953),
    .DE(net1572),
    .Q(\inst$top.soc.cpu.gprf.mem[9][20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][21]$_DFFE_PP_  (.CLK(clknet_leaf_487_clk_in_regs),
    .D(net950),
    .DE(net1574),
    .Q(\inst$top.soc.cpu.gprf.mem[9][21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][22]$_DFFE_PP_  (.CLK(clknet_leaf_366_clk_in_regs),
    .D(net948),
    .DE(net1572),
    .Q(\inst$top.soc.cpu.gprf.mem[9][22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][23]$_DFFE_PP_  (.CLK(clknet_leaf_405_clk_in_regs),
    .D(net941),
    .DE(net1572),
    .Q(\inst$top.soc.cpu.gprf.mem[9][23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][24]$_DFFE_PP_  (.CLK(clknet_leaf_482_clk_in_regs),
    .D(net938),
    .DE(net1574),
    .Q(\inst$top.soc.cpu.gprf.mem[9][24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][25]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk_in_regs),
    .D(net931),
    .DE(net1574),
    .Q(\inst$top.soc.cpu.gprf.mem[9][25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][26]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk_in_regs),
    .D(net925),
    .DE(net1572),
    .Q(\inst$top.soc.cpu.gprf.mem[9][26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][27]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk_in_regs),
    .D(net922),
    .DE(net1573),
    .Q(\inst$top.soc.cpu.gprf.mem[9][27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][28]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk_in_regs),
    .D(net917),
    .DE(net1573),
    .Q(\inst$top.soc.cpu.gprf.mem[9][28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][29]$_DFFE_PP_  (.CLK(clknet_leaf_493_clk_in_regs),
    .D(net912),
    .DE(net1574),
    .Q(\inst$top.soc.cpu.gprf.mem[9][29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk_in_regs),
    .D(net1061),
    .DE(net1572),
    .Q(\inst$top.soc.cpu.gprf.mem[9][2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][30]$_DFFE_PP_  (.CLK(clknet_leaf_434_clk_in_regs),
    .D(net908),
    .DE(net1575),
    .Q(\inst$top.soc.cpu.gprf.mem[9][30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][31]$_DFFE_PP_  (.CLK(clknet_leaf_448_clk_in_regs),
    .D(net904),
    .DE(net1574),
    .Q(\inst$top.soc.cpu.gprf.mem[9][31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk_in_regs),
    .D(net1056),
    .DE(net1573),
    .Q(\inst$top.soc.cpu.gprf.mem[9][3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk_in_regs),
    .D(net1011),
    .DE(net1575),
    .Q(\inst$top.soc.cpu.gprf.mem[9][4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk_in_regs),
    .D(net1052),
    .DE(net1574),
    .Q(\inst$top.soc.cpu.gprf.mem[9][5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk_in_regs),
    .D(net1049),
    .DE(net1574),
    .Q(\inst$top.soc.cpu.gprf.mem[9][6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk_in_regs),
    .D(net891),
    .DE(net1573),
    .Q(\inst$top.soc.cpu.gprf.mem[9][7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk_in_regs),
    .D(net1004),
    .DE(net1575),
    .Q(\inst$top.soc.cpu.gprf.mem[9][8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk_in_regs),
    .D(net1001),
    .DE(net1574),
    .Q(\inst$top.soc.cpu.gprf.mem[9][9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[0]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk_in_regs),
    .D(_00032_),
    .DE(net706),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[10]$_DFFE_PP_  (.CLK(clknet_leaf_408_clk_in_regs),
    .D(_00033_),
    .DE(net715),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[11]$_DFFE_PP_  (.CLK(clknet_leaf_412_clk_in_regs),
    .D(_00034_),
    .DE(net715),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[12]$_DFFE_PP_  (.CLK(clknet_leaf_497_clk_in_regs),
    .D(_00035_),
    .DE(net719),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[13]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk_in_regs),
    .D(_00036_),
    .DE(net716),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[14]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk_in_regs),
    .D(_00037_),
    .DE(net720),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[15]$_DFFE_PP_  (.CLK(clknet_leaf_438_clk_in_regs),
    .D(_00038_),
    .DE(net718),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[16]$_DFFE_PP_  (.CLK(clknet_leaf_508_clk_in_regs),
    .D(_00039_),
    .DE(net719),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[17]$_DFFE_PP_  (.CLK(clknet_leaf_445_clk_in_regs),
    .D(_00040_),
    .DE(net718),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[18]$_DFFE_PP_  (.CLK(clknet_leaf_366_clk_in_regs),
    .D(_00041_),
    .DE(net714),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[19]$_DFFE_PP_  (.CLK(clknet_leaf_449_clk_in_regs),
    .D(_00042_),
    .DE(net719),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[1]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk_in_regs),
    .D(_00043_),
    .DE(net706),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[20]$_DFFE_PP_  (.CLK(clknet_leaf_400_clk_in_regs),
    .D(_00044_),
    .DE(net716),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[21]$_DFFE_PP_  (.CLK(clknet_leaf_444_clk_in_regs),
    .D(_00045_),
    .DE(net718),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[22]$_DFFE_PP_  (.CLK(clknet_leaf_372_clk_in_regs),
    .D(_00046_),
    .DE(net713),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[23]$_DFFE_PP_  (.CLK(clknet_leaf_399_clk_in_regs),
    .D(_00047_),
    .DE(net715),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[24]$_DFFE_PP_  (.CLK(clknet_leaf_496_clk_in_regs),
    .D(_00048_),
    .DE(net719),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[25]$_DFFE_PP_  (.CLK(clknet_leaf_407_clk_in_regs),
    .D(_00049_),
    .DE(net716),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[26]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk_in_regs),
    .D(_00050_),
    .DE(net714),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[27]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk_in_regs),
    .D(_00051_),
    .DE(net720),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[28]$_DFFE_PP_  (.CLK(clknet_leaf_461_clk_in_regs),
    .D(_00052_),
    .DE(net719),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[29]$_DFFE_PP_  (.CLK(clknet_leaf_403_clk_in_regs),
    .D(_00053_),
    .DE(net718),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[2]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk_in_regs),
    .D(_00054_),
    .DE(net706),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[30]$_DFFE_PP_  (.CLK(clknet_leaf_419_clk_in_regs),
    .D(_00055_),
    .DE(net715),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[31]$_DFFE_PP_  (.CLK(clknet_leaf_441_clk_in_regs),
    .D(_00056_),
    .DE(net715),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[3]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk_in_regs),
    .D(_00057_),
    .DE(net717),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[4]$_DFFE_PP_  (.CLK(clknet_6_40__leaf_clk_in_regs),
    .D(_00058_),
    .DE(net706),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk_in_regs),
    .D(_00059_),
    .DE(net717),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[6]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk_in_regs),
    .D(_00060_),
    .DE(net716),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[7]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk_in_regs),
    .D(_00061_),
    .DE(net717),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[8]$_DFFE_PP_  (.CLK(clknet_leaf_427_clk_in_regs),
    .D(_00062_),
    .DE(net716),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp1__data[9]$_DFFE_PP_  (.CLK(clknet_leaf_426_clk_in_regs),
    .D(_00063_),
    .DE(net715),
    .Q(\inst$top.soc.cpu.gprf.mem_rp1__data[9] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[0]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk_in_regs),
    .D(_00000_),
    .DE(net706),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[0] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[10]$_DFFE_PP_  (.CLK(clknet_leaf_371_clk_in_regs),
    .D(_00001_),
    .DE(net712),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[10] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[11]$_DFFE_PP_  (.CLK(clknet_leaf_412_clk_in_regs),
    .D(_00002_),
    .DE(net715),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[11] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[12]$_DFFE_PP_  (.CLK(clknet_leaf_508_clk_in_regs),
    .D(_00003_),
    .DE(net719),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[12] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[13]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk_in_regs),
    .D(_00004_),
    .DE(net716),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[13] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[14]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk_in_regs),
    .D(_00005_),
    .DE(net717),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[14] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[15]$_DFFE_PP_  (.CLK(clknet_leaf_460_clk_in_regs),
    .D(_00006_),
    .DE(net717),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[15] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[16]$_DFFE_PP_  (.CLK(clknet_leaf_446_clk_in_regs),
    .D(_00007_),
    .DE(net718),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[16] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[17]$_DFFE_PP_  (.CLK(clknet_leaf_489_clk_in_regs),
    .D(_00008_),
    .DE(net719),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[17] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[18]$_DFFE_PP_  (.CLK(clknet_leaf_367_clk_in_regs),
    .D(_00009_),
    .DE(net712),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[18] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[19]$_DFFE_PP_  (.CLK(clknet_leaf_463_clk_in_regs),
    .D(_00010_),
    .DE(net718),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[19] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[1]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk_in_regs),
    .D(_00011_),
    .DE(net706),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[1] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[20]$_DFFE_PP_  (.CLK(clknet_leaf_405_clk_in_regs),
    .D(_00012_),
    .DE(net715),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[20] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[21]$_DFFE_PP_  (.CLK(clknet_leaf_449_clk_in_regs),
    .D(_00013_),
    .DE(net718),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[21] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[22]$_DFFE_PP_  (.CLK(clknet_leaf_371_clk_in_regs),
    .D(_00014_),
    .DE(net712),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[22] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[23]$_DFFE_PP_  (.CLK(clknet_leaf_395_clk_in_regs),
    .D(_00015_),
    .DE(net715),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[23] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[24]$_DFFE_PP_  (.CLK(clknet_leaf_497_clk_in_regs),
    .D(_00016_),
    .DE(net718),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[24] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[25]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk_in_regs),
    .D(_00017_),
    .DE(net706),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[25] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[26]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk_in_regs),
    .D(_00018_),
    .DE(net714),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[26] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[27]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk_in_regs),
    .D(_00019_),
    .DE(net717),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[27] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[28]$_DFFE_PP_  (.CLK(clknet_leaf_460_clk_in_regs),
    .D(_00020_),
    .DE(net717),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[28] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[29]$_DFFE_PP_  (.CLK(clknet_leaf_510_clk_in_regs),
    .D(_00021_),
    .DE(net718),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[29] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[2]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk_in_regs),
    .D(_00022_),
    .DE(net706),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[2] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[30]$_DFFE_PP_  (.CLK(clknet_leaf_428_clk_in_regs),
    .D(_00023_),
    .DE(net716),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[30] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[31]$_DFFE_PP_  (.CLK(clknet_leaf_439_clk_in_regs),
    .D(_00024_),
    .DE(net718),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[31] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[3]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk_in_regs),
    .D(_00025_),
    .DE(net717),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[3] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[4]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk_in_regs),
    .D(_00026_),
    .DE(net714),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[4] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk_in_regs),
    .D(_00027_),
    .DE(net717),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[5] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[6]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk_in_regs),
    .D(_00028_),
    .DE(net716),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[6] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[7]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk_in_regs),
    .D(_00029_),
    .DE(net717),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[7] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[8]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk_in_regs),
    .D(_00030_),
    .DE(net716),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[8] ));
 sky130_fd_sc_hd__edfxtp_1 \inst$top.soc.cpu.gprf.mem_rp2__data[9]$_DFFE_PP_  (.CLK(clknet_leaf_434_clk_in_regs),
    .D(_00031_),
    .DE(net715),
    .Q(\inst$top.soc.cpu.gprf.mem_rp2__data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_302_clk_in_regs),
    .D(_04184_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_351_clk_in_regs),
    .D(_04185_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_348_clk_in_regs),
    .D(_04186_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_373_clk_in_regs),
    .D(_04187_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_351_clk_in_regs),
    .D(_04188_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_358_clk_in_regs),
    .D(_04189_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_353_clk_in_regs),
    .D(_04190_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_381_clk_in_regs),
    .D(_04191_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_370_clk_in_regs),
    .D(_04192_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_353_clk_in_regs),
    .D(_04193_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_351_clk_in_regs),
    .D(_04194_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_339_clk_in_regs),
    .D(_04195_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_388_clk_in_regs),
    .D(_04196_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_373_clk_in_regs),
    .D(_04197_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_375_clk_in_regs),
    .D(_04198_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_388_clk_in_regs),
    .D(_04199_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_375_clk_in_regs),
    .D(_04200_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_381_clk_in_regs),
    .D(_04201_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_303_clk_in_regs),
    .D(_04202_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_363_clk_in_regs),
    .D(_04203_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_365_clk_in_regs),
    .D(_04204_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_388_clk_in_regs),
    .D(_04205_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_340_clk_in_regs),
    .D(_04206_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_353_clk_in_regs),
    .D(_04207_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_354_clk_in_regs),
    .D(_04208_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_341_clk_in_regs),
    .D(_04209_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_339_clk_in_regs),
    .D(_04210_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_302_clk_in_regs),
    .D(_04211_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_363_clk_in_regs),
    .D(_04212_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_356_clk_in_regs),
    .D(_04213_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_367_clk_in_regs),
    .D(_04214_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_data[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_360_clk_in_regs),
    .D(_04215_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass1_raw$_SDFFE_PP0P_  (.CLK(clknet_leaf_304_clk_in_regs),
    .D(_04216_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass1_raw ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_299_clk_in_regs),
    .D(_04217_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_353_clk_in_regs),
    .D(_04218_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_349_clk_in_regs),
    .D(_04219_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_371_clk_in_regs),
    .D(_04220_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[13]$_SDFFE_PP0P_  (.CLK(clknet_6_40__leaf_clk_in_regs),
    .D(_04221_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_299_clk_in_regs),
    .D(_04222_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_303_clk_in_regs),
    .D(_04223_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_379_clk_in_regs),
    .D(_04224_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_367_clk_in_regs),
    .D(_04225_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_302_clk_in_regs),
    .D(_04226_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_359_clk_in_regs),
    .D(_04227_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_303_clk_in_regs),
    .D(_04228_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_372_clk_in_regs),
    .D(_04229_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_371_clk_in_regs),
    .D(_04230_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_373_clk_in_regs),
    .D(_04231_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_379_clk_in_regs),
    .D(_04232_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_371_clk_in_regs),
    .D(_04233_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_305_clk_in_regs),
    .D(_04234_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_304_clk_in_regs),
    .D(_04235_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_305_clk_in_regs),
    .D(_04236_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_362_clk_in_regs),
    .D(_04237_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_373_clk_in_regs),
    .D(_04238_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_304_clk_in_regs),
    .D(_04239_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_358_clk_in_regs),
    .D(_04240_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_356_clk_in_regs),
    .D(_04241_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_304_clk_in_regs),
    .D(_04242_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_303_clk_in_regs),
    .D(_04243_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_299_clk_in_regs),
    .D(_04244_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_296_clk_in_regs),
    .D(_04245_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_305_clk_in_regs),
    .D(_04246_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_361_clk_in_regs),
    .D(_04247_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_data[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_362_clk_in_regs),
    .D(_04248_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.gprf.x_bypass2_raw$_SDFFE_PP0P_  (.CLK(clknet_leaf_300_clk_in_regs),
    .D(_04249_),
    .Q(\inst$top.soc.cpu.gprf.x_bypass2_raw ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_771_clk_in_regs),
    .D(_04250_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_768_clk_in_regs),
    .D(_04251_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_14_clk_in_regs),
    .D(_04252_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk_in_regs),
    .D(_04253_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_14_clk_in_regs),
    .D(_04254_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk_in_regs),
    .D(_04255_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk_in_regs),
    .D(_04256_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_769_clk_in_regs),
    .D(_04257_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_769_clk_in_regs),
    .D(_04258_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_770_clk_in_regs),
    .D(_04259_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_769_clk_in_regs),
    .D(_04260_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_772_clk_in_regs),
    .D(_04261_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_14_clk_in_regs),
    .D(_04262_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[21]$_SDFFE_PP0P_  (.CLK(clknet_6_25__leaf_clk_in_regs),
    .D(_04263_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_17_clk_in_regs),
    .D(_04264_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk_in_regs),
    .D(_04265_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk_in_regs),
    .D(_04266_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk_in_regs),
    .D(_04267_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_17_clk_in_regs),
    .D(_04268_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk_in_regs),
    .D(_04269_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_17_clk_in_regs),
    .D(_04270_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_771_clk_in_regs),
    .D(_04271_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_770_clk_in_regs),
    .D(_04272_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_772_clk_in_regs),
    .D(_04273_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_770_clk_in_regs),
    .D(_04274_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_765_clk_in_regs),
    .D(_04275_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk_in_regs),
    .D(_04276_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk_in_regs),
    .D(_04277_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk_in_regs),
    .D(_04278_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__adr[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_769_clk_in_regs),
    .D(_04279_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__adr[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__cyc$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk_in_regs),
    .D(_04280_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__cyc ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_72_clk_in_regs),
    .D(_04281_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk_in_regs),
    .D(_04282_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_67_clk_in_regs),
    .D(_04283_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk_in_regs),
    .D(_04284_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_44_clk_in_regs),
    .D(_04285_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_56_clk_in_regs),
    .D(_04286_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_55_clk_in_regs),
    .D(_04287_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk_in_regs),
    .D(_04288_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk_in_regs),
    .D(_04289_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk_in_regs),
    .D(_04290_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_317_clk_in_regs),
    .D(_04291_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_67_clk_in_regs),
    .D(_04292_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_45_clk_in_regs),
    .D(_04293_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_38_clk_in_regs),
    .D(_04294_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_45_clk_in_regs),
    .D(_04295_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk_in_regs),
    .D(_04296_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk_in_regs),
    .D(_04297_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk_in_regs),
    .D(_04298_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_71_clk_in_regs),
    .D(_04299_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_45_clk_in_regs),
    .D(_04300_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_72_clk_in_regs),
    .D(_04301_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_50_clk_in_regs),
    .D(_04302_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_38_clk_in_regs),
    .D(_04303_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_37_clk_in_regs),
    .D(_04304_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_44_clk_in_regs),
    .D(_04305_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk_in_regs),
    .D(_04306_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk_in_regs),
    .D(_04307_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_72_clk_in_regs),
    .D(_04308_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk_in_regs),
    .D(_04309_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_70_clk_in_regs),
    .D(_04310_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_38_clk_in_regs),
    .D(_04311_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__dat_w[9]$_SDFFE_PP0P_  (.CLK(clknet_6_32__leaf_clk_in_regs),
    .D(_04312_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__dat_w[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__sel[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk_in_regs),
    .D(_04313_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__sel[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__sel[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk_in_regs),
    .D(_04314_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__sel[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__sel[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_330_clk_in_regs),
    .D(_04315_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__sel[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_38_clk_in_regs),
    .D(_04316_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__sel[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__stb$_SDFFE_PP0P_  (.CLK(clknet_leaf_36_clk_in_regs),
    .D(_04317_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__stb ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.dbus__we$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk_in_regs),
    .D(_04318_),
    .Q(\inst$top.soc.cpu.loadstore.dbus__we ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk_in_regs),
    .D(_04319_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_317_clk_in_regs),
    .D(_04320_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_313_clk_in_regs),
    .D(_04321_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_313_clk_in_regs),
    .D(_04322_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_310_clk_in_regs),
    .D(_04323_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_273_clk_in_regs),
    .D(_04324_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_272_clk_in_regs),
    .D(_04325_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_271_clk_in_regs),
    .D(_04326_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_274_clk_in_regs),
    .D(_04327_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_87_clk_in_regs),
    .D(_04328_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_275_clk_in_regs),
    .D(_04329_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk_in_regs),
    .D(_04330_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_272_clk_in_regs),
    .D(_04331_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_272_clk_in_regs),
    .D(_04332_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_272_clk_in_regs),
    .D(_04333_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_311_clk_in_regs),
    .D(_04334_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_273_clk_in_regs),
    .D(_04335_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_309_clk_in_regs),
    .D(_04336_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_311_clk_in_regs),
    .D(_04337_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk_in_regs),
    .D(_04338_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk_in_regs),
    .D(_04339_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_273_clk_in_regs),
    .D(_04340_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk_in_regs),
    .D(_04341_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_276_clk_in_regs),
    .D(_04342_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_314_clk_in_regs),
    .D(_04343_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk_in_regs),
    .D(_04344_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk_in_regs),
    .D(_04345_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_314_clk_in_regs),
    .D(_04346_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_310_clk_in_regs),
    .D(_04347_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_314_clk_in_regs),
    .D(_04348_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_313_clk_in_regs),
    .D(_04349_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.loadstore.m_load_data[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_309_clk_in_regs),
    .D(_04350_),
    .Q(\inst$top.soc.cpu.loadstore.m_load_data[9] ));
 sky130_fd_sc_hd__dfxtp_2 \inst$top.soc.cpu.m.source__valid$_SDFF_PP0_  (.CLK(clknet_leaf_728_clk_in_regs),
    .D(_04351_),
    .Q(\inst$top.soc.cpu.m.source__valid ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_low$_SDFFE_PP0N_  (.CLK(clknet_leaf_346_clk_in_regs),
    .D(_04352_),
    .Q(\inst$top.soc.cpu.multiplier.m_low ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_561_clk_in_regs),
    .D(_04353_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[10]$_SDFFE_PP0N_  (.CLK(clknet_leaf_545_clk_in_regs),
    .D(_04354_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[11]$_SDFFE_PP0N_  (.CLK(clknet_leaf_545_clk_in_regs),
    .D(_04355_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[12]$_SDFFE_PP0N_  (.CLK(clknet_leaf_544_clk_in_regs),
    .D(_04356_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[13]$_SDFFE_PP0N_  (.CLK(clknet_6_23__leaf_clk_in_regs),
    .D(_04357_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[14]$_SDFFE_PP0N_  (.CLK(clknet_leaf_544_clk_in_regs),
    .D(_04358_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[15]$_SDFFE_PP0N_  (.CLK(clknet_leaf_544_clk_in_regs),
    .D(_04359_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[16]$_SDFFE_PP0N_  (.CLK(clknet_leaf_535_clk_in_regs),
    .D(_04360_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[17]$_SDFFE_PP0N_  (.CLK(clknet_leaf_535_clk_in_regs),
    .D(_04361_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[18]$_SDFFE_PP0N_  (.CLK(clknet_leaf_535_clk_in_regs),
    .D(_04362_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[19]$_SDFFE_PP0N_  (.CLK(clknet_leaf_534_clk_in_regs),
    .D(_04363_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_554_clk_in_regs),
    .D(_04364_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[20]$_SDFFE_PP0N_  (.CLK(clknet_leaf_527_clk_in_regs),
    .D(_04365_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[21]$_SDFFE_PP0N_  (.CLK(clknet_leaf_528_clk_in_regs),
    .D(_04366_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[22]$_SDFFE_PP0N_  (.CLK(clknet_leaf_529_clk_in_regs),
    .D(_04367_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[23]$_SDFFE_PP0N_  (.CLK(clknet_leaf_525_clk_in_regs),
    .D(_04368_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[24]$_SDFFE_PP0N_  (.CLK(clknet_leaf_527_clk_in_regs),
    .D(_04369_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[25]$_SDFFE_PP0N_  (.CLK(clknet_leaf_525_clk_in_regs),
    .D(_04370_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[26]$_SDFFE_PP0N_  (.CLK(clknet_6_47__leaf_clk_in_regs),
    .D(_04371_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[27]$_SDFFE_PP0N_  (.CLK(clknet_6_23__leaf_clk_in_regs),
    .D(_04372_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[28]$_SDFFE_PP0N_  (.CLK(clknet_leaf_515_clk_in_regs),
    .D(_04373_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[29]$_SDFFE_PP0N_  (.CLK(clknet_leaf_515_clk_in_regs),
    .D(_04374_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_554_clk_in_regs),
    .D(_04375_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[30]$_SDFFE_PP0N_  (.CLK(clknet_leaf_515_clk_in_regs),
    .D(_04376_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[31]$_SDFFE_PP0N_  (.CLK(clknet_6_53__leaf_clk_in_regs),
    .D(_04377_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[32]$_SDFFE_PP0N_  (.CLK(clknet_leaf_519_clk_in_regs),
    .D(_04378_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[32] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[33]$_SDFFE_PP0N_  (.CLK(clknet_leaf_542_clk_in_regs),
    .D(_04379_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[33] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[34]$_SDFFE_PP0N_  (.CLK(clknet_6_53__leaf_clk_in_regs),
    .D(_04380_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[34] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[35]$_SDFFE_PP0N_  (.CLK(clknet_leaf_554_clk_in_regs),
    .D(_04381_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[35] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[36]$_SDFFE_PP0N_  (.CLK(clknet_6_22__leaf_clk_in_regs),
    .D(_04382_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[36] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[37]$_SDFFE_PP0N_  (.CLK(clknet_6_53__leaf_clk_in_regs),
    .D(_04383_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[37] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[38]$_SDFFE_PP0N_  (.CLK(clknet_leaf_538_clk_in_regs),
    .D(_04384_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[38] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[39]$_SDFFE_PP0N_  (.CLK(clknet_leaf_544_clk_in_regs),
    .D(_04385_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[39] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_555_clk_in_regs),
    .D(_04386_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[40]$_SDFFE_PP0N_  (.CLK(clknet_leaf_533_clk_in_regs),
    .D(_04387_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[40] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[41]$_SDFFE_PP0N_  (.CLK(clknet_leaf_535_clk_in_regs),
    .D(_04388_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[41] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[42]$_SDFFE_PP0N_  (.CLK(clknet_leaf_538_clk_in_regs),
    .D(_04389_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[42] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[43]$_SDFFE_PP0N_  (.CLK(clknet_leaf_538_clk_in_regs),
    .D(_04390_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[43] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[44]$_SDFFE_PP0N_  (.CLK(clknet_leaf_532_clk_in_regs),
    .D(_04391_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[44] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[45]$_SDFFE_PP0N_  (.CLK(clknet_leaf_537_clk_in_regs),
    .D(_04392_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[45] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[46]$_SDFFE_PP0N_  (.CLK(clknet_leaf_536_clk_in_regs),
    .D(_04393_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[46] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[47]$_SDFFE_PP0N_  (.CLK(clknet_leaf_537_clk_in_regs),
    .D(_04394_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[47] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[48]$_SDFFE_PP0N_  (.CLK(clknet_leaf_536_clk_in_regs),
    .D(_04395_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[48] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[49]$_SDFFE_PP0N_  (.CLK(clknet_leaf_529_clk_in_regs),
    .D(_04396_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[49] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_555_clk_in_regs),
    .D(_04397_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[50]$_SDFFE_PP0N_  (.CLK(clknet_leaf_536_clk_in_regs),
    .D(_04398_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[50] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[51]$_SDFFE_PP0N_  (.CLK(clknet_leaf_534_clk_in_regs),
    .D(_04399_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[51] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[52]$_SDFFE_PP0N_  (.CLK(clknet_leaf_530_clk_in_regs),
    .D(_04400_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[52] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[53]$_SDFFE_PP0N_  (.CLK(clknet_leaf_533_clk_in_regs),
    .D(_04401_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[53] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[54]$_SDFFE_PP0N_  (.CLK(clknet_leaf_530_clk_in_regs),
    .D(_04402_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[54] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[55]$_SDFFE_PP0N_  (.CLK(clknet_leaf_528_clk_in_regs),
    .D(_04403_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[55] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[56]$_SDFFE_PP0N_  (.CLK(clknet_leaf_531_clk_in_regs),
    .D(_04404_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[56] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[57]$_SDFFE_PP0N_  (.CLK(clknet_6_53__leaf_clk_in_regs),
    .D(_04405_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[57] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[58]$_SDFFE_PP0N_  (.CLK(clknet_leaf_532_clk_in_regs),
    .D(_04406_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[58] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[59]$_SDFFE_PP0N_  (.CLK(clknet_6_23__leaf_clk_in_regs),
    .D(_04407_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[59] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_555_clk_in_regs),
    .D(_04408_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[60]$_SDFFE_PP0N_  (.CLK(clknet_leaf_531_clk_in_regs),
    .D(_04409_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[60] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[61]$_SDFFE_PP0N_  (.CLK(clknet_leaf_531_clk_in_regs),
    .D(_04410_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[61] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[62]$_SDFFE_PP0N_  (.CLK(clknet_leaf_529_clk_in_regs),
    .D(_04411_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[62] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[63]$_SDFFE_PP0N_  (.CLK(clknet_leaf_542_clk_in_regs),
    .D(_04412_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[63] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[6]$_SDFFE_PP0N_  (.CLK(clknet_leaf_543_clk_in_regs),
    .D(_04413_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[7]$_SDFFE_PP0N_  (.CLK(clknet_leaf_543_clk_in_regs),
    .D(_04414_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[8]$_SDFFE_PP0N_  (.CLK(clknet_leaf_543_clk_in_regs),
    .D(_04415_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.m_prod[9]$_SDFFE_PP0N_  (.CLK(clknet_leaf_545_clk_in_regs),
    .D(_04416_),
    .Q(\inst$top.soc.cpu.multiplier.m_prod[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_561_clk_in_regs),
    .D(_04417_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[10]$_SDFFE_PP0N_  (.CLK(clknet_leaf_350_clk_in_regs),
    .D(_04418_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[11]$_SDFFE_PP0N_  (.CLK(clknet_leaf_562_clk_in_regs),
    .D(_04419_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[12]$_SDFFE_PP0N_  (.CLK(clknet_6_46__leaf_clk_in_regs),
    .D(_04420_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[13]$_SDFFE_PP0N_  (.CLK(clknet_leaf_561_clk_in_regs),
    .D(_04421_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[14]$_SDFFE_PP0N_  (.CLK(clknet_leaf_561_clk_in_regs),
    .D(_04422_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[15]$_SDFFE_PP0N_  (.CLK(clknet_6_22__leaf_clk_in_regs),
    .D(_04423_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[16]$_SDFFE_PP0N_  (.CLK(clknet_leaf_559_clk_in_regs),
    .D(_04424_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[17]$_SDFFE_PP0N_  (.CLK(clknet_leaf_560_clk_in_regs),
    .D(_04425_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[18]$_SDFFE_PP0N_  (.CLK(clknet_6_45__leaf_clk_in_regs),
    .D(_04426_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[19]$_SDFFE_PP0N_  (.CLK(clknet_leaf_559_clk_in_regs),
    .D(_04427_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_557_clk_in_regs),
    .D(_04428_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[20]$_SDFFE_PP0N_  (.CLK(clknet_leaf_560_clk_in_regs),
    .D(_04429_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[21]$_SDFFE_PP0N_  (.CLK(clknet_leaf_520_clk_in_regs),
    .D(_04430_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[22]$_SDFFE_PP0N_  (.CLK(clknet_leaf_519_clk_in_regs),
    .D(_04431_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[23]$_SDFFE_PP0N_  (.CLK(clknet_leaf_520_clk_in_regs),
    .D(_04432_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[24]$_SDFFE_PP0N_  (.CLK(clknet_6_46__leaf_clk_in_regs),
    .D(_04433_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[25]$_SDFFE_PP0N_  (.CLK(clknet_leaf_520_clk_in_regs),
    .D(_04434_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[26]$_SDFFE_PP0N_  (.CLK(clknet_6_22__leaf_clk_in_regs),
    .D(_04435_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[27]$_SDFFE_PP0N_  (.CLK(clknet_leaf_557_clk_in_regs),
    .D(_04436_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[28]$_SDFFE_PP0N_  (.CLK(clknet_leaf_368_clk_in_regs),
    .D(_04437_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[29]$_SDFFE_PP0N_  (.CLK(clknet_leaf_520_clk_in_regs),
    .D(_04438_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[2]$_SDFFE_PP0N_  (.CLK(clknet_6_22__leaf_clk_in_regs),
    .D(_04439_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[30]$_SDFFE_PP0N_  (.CLK(clknet_leaf_560_clk_in_regs),
    .D(_04440_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[31]$_SDFFE_PP0N_  (.CLK(clknet_leaf_557_clk_in_regs),
    .D(_04441_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_347_clk_in_regs),
    .D(_04442_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_347_clk_in_regs),
    .D(_04443_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_561_clk_in_regs),
    .D(_04444_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[6]$_SDFFE_PP0N_  (.CLK(clknet_leaf_383_clk_in_regs),
    .D(_04445_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[7]$_SDFFE_PP0N_  (.CLK(clknet_leaf_348_clk_in_regs),
    .D(_04446_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[8]$_SDFFE_PP0N_  (.CLK(clknet_leaf_384_clk_in_regs),
    .D(_04447_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.w_result[9]$_SDFFE_PP0N_  (.CLK(clknet_leaf_359_clk_in_regs),
    .D(_04448_),
    .Q(\inst$top.soc.cpu.multiplier.w_result[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.x_low$_SDFFE_PP0P_  (.CLK(clknet_leaf_341_clk_in_regs),
    .D(_04449_),
    .Q(\inst$top.soc.cpu.multiplier.x_low ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.x_src1_signed$_SDFFE_PP0P_  (.CLK(clknet_leaf_343_clk_in_regs),
    .D(_04450_),
    .Q(\inst$top.soc.cpu.multiplier.x_src1_signed ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.multiplier.x_src2_signed$_SDFFE_PP0P_  (.CLK(clknet_leaf_575_clk_in_regs),
    .D(_04451_),
    .Q(\inst$top.soc.cpu.multiplier.x_src2_signed ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_direction$_SDFFE_PP0N_  (.CLK(clknet_leaf_391_clk_in_regs),
    .D(_04452_),
    .Q(\inst$top.soc.cpu.shifter.m_direction ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_413_clk_in_regs),
    .D(_04453_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[10]$_SDFFE_PP0N_  (.CLK(clknet_leaf_391_clk_in_regs),
    .D(_04454_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[11]$_SDFFE_PP0N_  (.CLK(clknet_leaf_390_clk_in_regs),
    .D(_04455_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[12]$_SDFFE_PP0N_  (.CLK(clknet_leaf_390_clk_in_regs),
    .D(_04456_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[13]$_SDFFE_PP0N_  (.CLK(clknet_leaf_389_clk_in_regs),
    .D(_04457_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[14]$_SDFFE_PP0N_  (.CLK(clknet_leaf_374_clk_in_regs),
    .D(_04458_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[15]$_SDFFE_PP0N_  (.CLK(clknet_leaf_414_clk_in_regs),
    .D(_04459_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[16]$_SDFFE_PP0N_  (.CLK(clknet_leaf_383_clk_in_regs),
    .D(_04460_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[17]$_SDFFE_PP0N_  (.CLK(clknet_leaf_390_clk_in_regs),
    .D(_04461_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[18]$_SDFFE_PP0N_  (.CLK(clknet_leaf_385_clk_in_regs),
    .D(_04462_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[19]$_SDFFE_PP0N_  (.CLK(clknet_leaf_388_clk_in_regs),
    .D(_04463_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_414_clk_in_regs),
    .D(_04464_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[20]$_SDFFE_PP0N_  (.CLK(clknet_leaf_387_clk_in_regs),
    .D(_16380_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[21]$_SDFFE_PP0N_  (.CLK(clknet_leaf_392_clk_in_regs),
    .D(_16384_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[22]$_SDFFE_PP0N_  (.CLK(clknet_leaf_389_clk_in_regs),
    .D(_16388_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[23]$_SDFFE_PP0N_  (.CLK(clknet_leaf_390_clk_in_regs),
    .D(_04468_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[24]$_SDFFE_PP0N_  (.CLK(clknet_leaf_393_clk_in_regs),
    .D(_04469_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[25]$_SDFFE_PP0N_  (.CLK(clknet_leaf_387_clk_in_regs),
    .D(_04470_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[26]$_SDFFE_PP0N_  (.CLK(clknet_leaf_387_clk_in_regs),
    .D(_04471_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[27]$_SDFFE_PP0N_  (.CLK(clknet_leaf_392_clk_in_regs),
    .D(_04472_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[28]$_SDFFE_PP0N_  (.CLK(clknet_leaf_390_clk_in_regs),
    .D(_04473_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[29]$_SDFFE_PP0N_  (.CLK(clknet_leaf_413_clk_in_regs),
    .D(_04474_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_374_clk_in_regs),
    .D(_04475_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[30]$_SDFFE_PP0N_  (.CLK(clknet_leaf_375_clk_in_regs),
    .D(_16411_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[31]$_SDFFE_PP0N_  (.CLK(clknet_leaf_374_clk_in_regs),
    .D(_04477_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_390_clk_in_regs),
    .D(_04478_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_389_clk_in_regs),
    .D(_04479_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_393_clk_in_regs),
    .D(_04480_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[6]$_SDFFE_PP0N_  (.CLK(clknet_leaf_391_clk_in_regs),
    .D(_04481_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[7]$_SDFFE_PP0N_  (.CLK(clknet_leaf_390_clk_in_regs),
    .D(_04482_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[8]$_SDFFE_PP0N_  (.CLK(clknet_leaf_412_clk_in_regs),
    .D(_04483_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.shifter.m_result$7[9]$_SDFFE_PP0N_  (.CLK(clknet_leaf_392_clk_in_regs),
    .D(_04484_),
    .Q(\inst$top.soc.cpu.shifter.m_result$7[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[100]$_SDFFE_PP0P_  (.CLK(clknet_leaf_319_clk_in_regs),
    .D(_04485_),
    .Q(\inst$top.soc.cpu.sink__payload$12[100] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[101]$_SDFFE_PP0P_  (.CLK(clknet_leaf_342_clk_in_regs),
    .D(_04486_),
    .Q(\inst$top.soc.cpu.sink__payload$12[101] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[102]$_SDFFE_PP0P_  (.CLK(clknet_leaf_342_clk_in_regs),
    .D(_04487_),
    .Q(\inst$top.soc.cpu.sink__payload$12[102] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[103]$_SDFFE_PP0P_  (.CLK(clknet_leaf_345_clk_in_regs),
    .D(_04488_),
    .Q(\inst$top.soc.cpu.sink__payload$12[103] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[104]$_SDFFE_PP0P_  (.CLK(clknet_leaf_580_clk_in_regs),
    .D(_04489_),
    .Q(\inst$top.soc.cpu.sink__payload$12[104] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[105]$_SDFFE_PP0P_  (.CLK(clknet_leaf_578_clk_in_regs),
    .D(_04490_),
    .Q(\inst$top.soc.cpu.sink__payload$12[105] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[106]$_SDFFE_PP0P_  (.CLK(clknet_leaf_324_clk_in_regs),
    .D(_04491_),
    .Q(\inst$top.soc.cpu.d.sink__payload.rd_we ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[107]$_SDFFE_PP0P_  (.CLK(clknet_leaf_588_clk_in_regs),
    .D(_04492_),
    .Q(\inst$top.soc.cpu.d.sink__payload.rs1_re ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[108]$_SDFFE_PP0P_  (.CLK(clknet_leaf_333_clk_in_regs),
    .D(_04493_),
    .Q(\inst$top.soc.cpu.d.sink__payload.rs2_re ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_755_clk_in_regs),
    .D(_04494_),
    .Q(\inst$top.soc.cpu.sink__payload$12[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[111]$_SDFFE_PP0P_  (.CLK(clknet_leaf_327_clk_in_regs),
    .D(_04495_),
    .Q(\inst$top.soc.cpu.sink__payload$12[111] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[112]$_SDFFE_PP0P_  (.CLK(clknet_6_39__leaf_clk_in_regs),
    .D(_04496_),
    .Q(\inst$top.soc.cpu.sink__payload$12[112] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[113]$_SDFFE_PP0P_  (.CLK(clknet_leaf_327_clk_in_regs),
    .D(_04497_),
    .Q(\inst$top.soc.cpu.sink__payload$12[113] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[114]$_SDFFE_PP0P_  (.CLK(clknet_leaf_327_clk_in_regs),
    .D(_04498_),
    .Q(\inst$top.soc.cpu.sink__payload$12[114] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[115]$_SDFFE_PP0P_  (.CLK(clknet_leaf_332_clk_in_regs),
    .D(_04499_),
    .Q(\inst$top.soc.cpu.sink__payload$12[115] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[116]$_SDFFE_PP0P_  (.CLK(clknet_leaf_334_clk_in_regs),
    .D(_04500_),
    .Q(\inst$top.soc.cpu.sink__payload$12[116] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[117]$_SDFFE_PP0P_  (.CLK(clknet_leaf_333_clk_in_regs),
    .D(_04501_),
    .Q(\inst$top.soc.cpu.sink__payload$12[117] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[118]$_SDFFE_PP0P_  (.CLK(clknet_leaf_335_clk_in_regs),
    .D(_04502_),
    .Q(\inst$top.soc.cpu.sink__payload$12[118] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[119]$_SDFFE_PP0P_  (.CLK(clknet_leaf_337_clk_in_regs),
    .D(_04503_),
    .Q(\inst$top.soc.cpu.sink__payload$12[119] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_590_clk_in_regs),
    .D(_04504_),
    .Q(\inst$top.soc.cpu.sink__payload$12[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[120]$_SDFFE_PP0P_  (.CLK(clknet_leaf_344_clk_in_regs),
    .D(_04505_),
    .Q(\inst$top.soc.cpu.sink__payload$12[120] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[121]$_SDFFE_PP0P_  (.CLK(clknet_leaf_337_clk_in_regs),
    .D(_04506_),
    .Q(\inst$top.soc.cpu.sink__payload$12[121] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[122]$_SDFFE_PP0P_  (.CLK(clknet_leaf_329_clk_in_regs),
    .D(_04507_),
    .Q(\inst$top.soc.cpu.sink__payload$12[122] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[123]$_SDFFE_PP0P_  (.CLK(clknet_leaf_332_clk_in_regs),
    .D(_04508_),
    .Q(\inst$top.soc.cpu.sink__payload$12[123] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[124]$_SDFFE_PP0P_  (.CLK(clknet_leaf_325_clk_in_regs),
    .D(_04509_),
    .Q(\inst$top.soc.cpu.sink__payload$12[124] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[125]$_SDFFE_PP0P_  (.CLK(clknet_leaf_324_clk_in_regs),
    .D(_04510_),
    .Q(\inst$top.soc.cpu.sink__payload$12[125] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[126]$_SDFFE_PP0P_  (.CLK(clknet_leaf_325_clk_in_regs),
    .D(_04511_),
    .Q(\inst$top.soc.cpu.sink__payload$12[126] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[127]$_SDFFE_PP0P_  (.CLK(clknet_leaf_319_clk_in_regs),
    .D(_04512_),
    .Q(\inst$top.soc.cpu.sink__payload$12[127] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[128]$_SDFFE_PP0P_  (.CLK(clknet_leaf_325_clk_in_regs),
    .D(_04513_),
    .Q(\inst$top.soc.cpu.sink__payload$12[128] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[129]$_SDFFE_PP0P_  (.CLK(clknet_leaf_332_clk_in_regs),
    .D(_04514_),
    .Q(\inst$top.soc.cpu.sink__payload$12[129] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_593_clk_in_regs),
    .D(_04515_),
    .Q(\inst$top.soc.cpu.sink__payload$12[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[130]$_SDFFE_PP0P_  (.CLK(clknet_leaf_328_clk_in_regs),
    .D(_04516_),
    .Q(\inst$top.soc.cpu.sink__payload$12[130] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[131]$_SDFFE_PP0P_  (.CLK(clknet_leaf_328_clk_in_regs),
    .D(_04517_),
    .Q(\inst$top.soc.cpu.sink__payload$12[131] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[132]$_SDFFE_PP0P_  (.CLK(clknet_leaf_327_clk_in_regs),
    .D(_04518_),
    .Q(\inst$top.soc.cpu.sink__payload$12[132] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[133]$_SDFFE_PP0P_  (.CLK(clknet_leaf_330_clk_in_regs),
    .D(_04519_),
    .Q(\inst$top.soc.cpu.sink__payload$12[133] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[134]$_SDFFE_PP0P_  (.CLK(clknet_leaf_329_clk_in_regs),
    .D(_04520_),
    .Q(\inst$top.soc.cpu.sink__payload$12[134] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[135]$_SDFFE_PP0P_  (.CLK(clknet_leaf_331_clk_in_regs),
    .D(_04521_),
    .Q(\inst$top.soc.cpu.sink__payload$12[135] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[136]$_SDFFE_PP0P_  (.CLK(clknet_leaf_330_clk_in_regs),
    .D(_04522_),
    .Q(\inst$top.soc.cpu.sink__payload$12[136] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[137]$_SDFFE_PP0P_  (.CLK(clknet_leaf_331_clk_in_regs),
    .D(_04523_),
    .Q(\inst$top.soc.cpu.sink__payload$12[137] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[138]$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk_in_regs),
    .D(_04524_),
    .Q(\inst$top.soc.cpu.sink__payload$12[138] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[139]$_SDFFE_PP0P_  (.CLK(clknet_leaf_333_clk_in_regs),
    .D(_04525_),
    .Q(\inst$top.soc.cpu.sink__payload$12[139] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_589_clk_in_regs),
    .D(_04526_),
    .Q(\inst$top.soc.cpu.sink__payload$12[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[140]$_SDFFE_PP0P_  (.CLK(clknet_leaf_340_clk_in_regs),
    .D(_04527_),
    .Q(\inst$top.soc.cpu.sink__payload$12[140] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[141]$_SDFFE_PP0P_  (.CLK(clknet_leaf_340_clk_in_regs),
    .D(_04528_),
    .Q(\inst$top.soc.cpu.d.sink__payload.bypass_x ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[142]$_SDFFE_PP0P_  (.CLK(clknet_leaf_340_clk_in_regs),
    .D(_04529_),
    .Q(\inst$top.soc.cpu.d.sink__payload.bypass_m ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[143]$_SDFFE_PP0P_  (.CLK(clknet_leaf_329_clk_in_regs),
    .D(_04530_),
    .Q(\inst$top.soc.cpu.sink__payload$12[143] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[144]$_SDFFE_PP0P_  (.CLK(clknet_leaf_330_clk_in_regs),
    .D(_04531_),
    .Q(\inst$top.soc.cpu.sink__payload$12[144] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[146]$_SDFFE_PP0P_  (.CLK(clknet_leaf_343_clk_in_regs),
    .D(_04532_),
    .Q(\inst$top.soc.cpu.d.sink__payload.lui ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[147]$_SDFFE_PP0P_  (.CLK(clknet_leaf_343_clk_in_regs),
    .D(_04533_),
    .Q(\inst$top.soc.cpu.d.sink__payload.auipc ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[148]$_SDFFE_PP0P_  (.CLK(clknet_leaf_335_clk_in_regs),
    .D(_04534_),
    .Q(\inst$top.soc.cpu.d.sink__payload.load ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[149]$_SDFFE_PP0P_  (.CLK(clknet_leaf_332_clk_in_regs),
    .D(_04535_),
    .Q(\inst$top.soc.cpu.d.sink__payload.store ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_754_clk_in_regs),
    .D(_04536_),
    .Q(\inst$top.soc.cpu.sink__payload$12[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[150]$_SDFFE_PP0P_  (.CLK(clknet_leaf_574_clk_in_regs),
    .D(_04537_),
    .Q(\inst$top.soc.cpu.adder$307.x_sub ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[151]$_SDFFE_PP0P_  (.CLK(clknet_leaf_584_clk_in_regs),
    .D(_04538_),
    .Q(\inst$top.soc.cpu.d.sink__payload.logic ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[152]$_SDFFE_PP0P_  (.CLK(clknet_leaf_343_clk_in_regs),
    .D(_04539_),
    .Q(\inst$top.soc.cpu.d.sink__payload.multiply ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[153]$_SDFFE_PP0P_  (.CLK(clknet_leaf_585_clk_in_regs),
    .D(_04540_),
    .Q(\inst$top.soc.cpu.d.sink__payload.divide ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[154]$_SDFFE_PP0P_  (.CLK(clknet_leaf_344_clk_in_regs),
    .D(_04541_),
    .Q(\inst$top.soc.cpu.d.sink__payload.shift ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[155]$_SDFFE_PP0P_  (.CLK(clknet_leaf_391_clk_in_regs),
    .D(_04542_),
    .Q(\inst$top.soc.cpu.d.sink__payload.direction ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[156]$_SDFFE_PP0P_  (.CLK(clknet_6_31__leaf_clk_in_regs),
    .D(_04543_),
    .Q(\inst$top.soc.cpu.d.sink__payload.sext ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[157]$_SDFFE_PP0P_  (.CLK(clknet_leaf_586_clk_in_regs),
    .D(_04544_),
    .Q(\inst$top.soc.cpu.d.sink__payload.jump ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[158]$_SDFFE_PP0P_  (.CLK(clknet_6_27__leaf_clk_in_regs),
    .D(_04545_),
    .Q(\inst$top.soc.cpu.d.sink__payload.compare ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[159]$_SDFFE_PP0P_  (.CLK(clknet_leaf_344_clk_in_regs),
    .D(_04546_),
    .Q(\inst$top.soc.cpu.d.sink__payload.branch ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_334_clk_in_regs),
    .D(_04547_),
    .Q(\inst$top.soc.cpu.sink__payload$12[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[160]$_SDFFE_PP0P_  (.CLK(clknet_leaf_730_clk_in_regs),
    .D(_04548_),
    .Q(\inst$top.soc.cpu.sink__payload$12[109] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[161]$_SDFFE_PP0P_  (.CLK(clknet_leaf_586_clk_in_regs),
    .D(_04549_),
    .Q(\inst$top.soc.cpu.sink__payload$12[110] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[162]$_SDFFE_PP0P_  (.CLK(clknet_leaf_728_clk_in_regs),
    .D(_04550_),
    .Q(\inst$top.soc.cpu.sink__payload$12[162] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[163]$_SDFFE_PP0P_  (.CLK(clknet_leaf_728_clk_in_regs),
    .D(_04551_),
    .Q(\inst$top.soc.cpu.sink__payload$12[163] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[164]$_SDFFE_PP0P_  (.CLK(clknet_leaf_726_clk_in_regs),
    .D(_04552_),
    .Q(\inst$top.soc.cpu.sink__payload$12[164] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[165]$_SDFFE_PP0P_  (.CLK(clknet_leaf_748_clk_in_regs),
    .D(_04553_),
    .Q(\inst$top.soc.cpu.sink__payload$12[165] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[166]$_SDFFE_PP0P_  (.CLK(clknet_leaf_749_clk_in_regs),
    .D(_04554_),
    .Q(\inst$top.soc.cpu.sink__payload$12[166] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[167]$_SDFFE_PP0P_  (.CLK(clknet_leaf_727_clk_in_regs),
    .D(_04555_),
    .Q(\inst$top.soc.cpu.sink__payload$12[167] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[168]$_SDFFE_PP0P_  (.CLK(clknet_leaf_753_clk_in_regs),
    .D(_04556_),
    .Q(\inst$top.soc.cpu.sink__payload$12[168] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[169]$_SDFFE_PP0P_  (.CLK(clknet_leaf_753_clk_in_regs),
    .D(_04557_),
    .Q(\inst$top.soc.cpu.sink__payload$12[169] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_333_clk_in_regs),
    .D(_04558_),
    .Q(\inst$top.soc.cpu.sink__payload$12[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[170]$_SDFFE_PP0P_  (.CLK(clknet_leaf_756_clk_in_regs),
    .D(_04559_),
    .Q(\inst$top.soc.cpu.sink__payload$12[170] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[171]$_SDFFE_PP0P_  (.CLK(clknet_leaf_750_clk_in_regs),
    .D(_04560_),
    .Q(\inst$top.soc.cpu.sink__payload$12[171] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[172]$_SDFFE_PP0P_  (.CLK(clknet_leaf_753_clk_in_regs),
    .D(_04561_),
    .Q(\inst$top.soc.cpu.sink__payload$12[172] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[173]$_SDFFE_PP0P_  (.CLK(clknet_leaf_755_clk_in_regs),
    .D(_04562_),
    .Q(\inst$top.soc.cpu.sink__payload$12[173] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[174]$_SDFFE_PP0P_  (.CLK(clknet_leaf_756_clk_in_regs),
    .D(_04563_),
    .Q(\inst$top.soc.cpu.sink__payload$12[174] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[175]$_SDFFE_PP0P_  (.CLK(clknet_leaf_594_clk_in_regs),
    .D(_04564_),
    .Q(\inst$top.soc.cpu.sink__payload$12[175] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[176]$_SDFFE_PP0P_  (.CLK(clknet_leaf_753_clk_in_regs),
    .D(_04565_),
    .Q(\inst$top.soc.cpu.sink__payload$12[176] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[177]$_SDFFE_PP0P_  (.CLK(clknet_leaf_753_clk_in_regs),
    .D(_04566_),
    .Q(\inst$top.soc.cpu.sink__payload$12[177] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[178]$_SDFFE_PP0P_  (.CLK(clknet_leaf_764_clk_in_regs),
    .D(_04567_),
    .Q(\inst$top.soc.cpu.sink__payload$12[178] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[179]$_SDFFE_PP0P_  (.CLK(clknet_leaf_726_clk_in_regs),
    .D(_04568_),
    .Q(\inst$top.soc.cpu.sink__payload$12[179] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk_in_regs),
    .D(_04569_),
    .Q(\inst$top.soc.cpu.sink__payload$12[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[180]$_SDFFE_PP0P_  (.CLK(clknet_leaf_751_clk_in_regs),
    .D(_04570_),
    .Q(\inst$top.soc.cpu.sink__payload$12[180] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[181]$_SDFFE_PP0P_  (.CLK(clknet_leaf_762_clk_in_regs),
    .D(_04571_),
    .Q(\inst$top.soc.cpu.sink__payload$12[181] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[182]$_SDFFE_PP0P_  (.CLK(clknet_leaf_755_clk_in_regs),
    .D(_04572_),
    .Q(\inst$top.soc.cpu.sink__payload$12[182] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[183]$_SDFFE_PP0P_  (.CLK(clknet_leaf_757_clk_in_regs),
    .D(_04573_),
    .Q(\inst$top.soc.cpu.sink__payload$12[183] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[184]$_SDFFE_PP0P_  (.CLK(clknet_leaf_757_clk_in_regs),
    .D(_04574_),
    .Q(\inst$top.soc.cpu.sink__payload$12[184] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[185]$_SDFFE_PP0P_  (.CLK(clknet_leaf_779_clk_in_regs),
    .D(_04575_),
    .Q(\inst$top.soc.cpu.sink__payload$12[185] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[186]$_SDFFE_PP0P_  (.CLK(clknet_leaf_589_clk_in_regs),
    .D(_04576_),
    .Q(\inst$top.soc.cpu.sink__payload$12[186] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[187]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk_in_regs),
    .D(_04577_),
    .Q(\inst$top.soc.cpu.sink__payload$12[187] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[188]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk_in_regs),
    .D(_04578_),
    .Q(\inst$top.soc.cpu.sink__payload$12[188] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[189]$_SDFFE_PP0P_  (.CLK(clknet_leaf_758_clk_in_regs),
    .D(_04579_),
    .Q(\inst$top.soc.cpu.sink__payload$12[189] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_764_clk_in_regs),
    .D(_04580_),
    .Q(\inst$top.soc.cpu.sink__payload$12[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[190]$_SDFFE_PP0P_  (.CLK(clknet_leaf_758_clk_in_regs),
    .D(_04581_),
    .Q(\inst$top.soc.cpu.sink__payload$12[190] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[191]$_SDFFE_PP0P_  (.CLK(clknet_leaf_779_clk_in_regs),
    .D(_04582_),
    .Q(\inst$top.soc.cpu.sink__payload$12[191] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[192]$_SDFFE_PP0P_  (.CLK(clknet_6_12__leaf_clk_in_regs),
    .D(_04583_),
    .Q(\inst$top.soc.cpu.d.sink__payload.branch_predict_taken ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[193]$_SDFFE_PP0P_  (.CLK(clknet_leaf_758_clk_in_regs),
    .D(_04584_),
    .Q(\inst$top.soc.cpu.d.sink__payload.fence_i ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[194]$_SDFFE_PP0P_  (.CLK(clknet_leaf_343_clk_in_regs),
    .D(_04585_),
    .Q(\inst$top.soc.cpu.d.sink__payload.csr_re ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[195]$_SDFFE_PP0P_  (.CLK(clknet_leaf_334_clk_in_regs),
    .D(_04586_),
    .Q(\inst$top.soc.cpu.d.sink__payload.csr_we ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[196]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk_in_regs),
    .D(_04587_),
    .Q(\inst$top.soc.cpu.d.sink__payload.csr_fmt_i ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[197]$_SDFFE_PP0P_  (.CLK(clknet_leaf_585_clk_in_regs),
    .D(_04588_),
    .Q(\inst$top.soc.cpu.d.sink__payload.csr_set ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[198]$_SDFFE_PP0P_  (.CLK(clknet_leaf_584_clk_in_regs),
    .D(_04589_),
    .Q(\inst$top.soc.cpu.d.sink__payload.csr_clear ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[199]$_SDFFE_PP0P_  (.CLK(clknet_leaf_586_clk_in_regs),
    .D(_04590_),
    .Q(\inst$top.soc.cpu.d.sink__payload.ecall ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk_in_regs),
    .D(_04591_),
    .Q(\inst$top.soc.cpu.sink__payload$12[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[200]$_SDFFE_PP0P_  (.CLK(clknet_leaf_588_clk_in_regs),
    .D(_04592_),
    .Q(\inst$top.soc.cpu.d.sink__payload.ebreak ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[201]$_SDFFE_PP0P_  (.CLK(clknet_leaf_591_clk_in_regs),
    .D(_04593_),
    .Q(\inst$top.soc.cpu.d.sink__payload.mret ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_777_clk_in_regs),
    .D(_04594_),
    .Q(\inst$top.soc.cpu.sink__payload$12[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_767_clk_in_regs),
    .D(_04595_),
    .Q(\inst$top.soc.cpu.sink__payload$12[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk_in_regs),
    .D(_04596_),
    .Q(\inst$top.soc.cpu.sink__payload$12[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk_in_regs),
    .D(_04597_),
    .Q(\inst$top.soc.cpu.sink__payload$12[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk_in_regs),
    .D(_04598_),
    .Q(\inst$top.soc.cpu.sink__payload$12[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk_in_regs),
    .D(_04599_),
    .Q(\inst$top.soc.cpu.sink__payload$12[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk_in_regs),
    .D(_04600_),
    .Q(\inst$top.soc.cpu.sink__payload$12[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk_in_regs),
    .D(_04601_),
    .Q(\inst$top.soc.cpu.sink__payload$12[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk_in_regs),
    .D(_04602_),
    .Q(\inst$top.soc.cpu.sink__payload$12[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk_in_regs),
    .D(_04603_),
    .Q(\inst$top.soc.cpu.sink__payload$12[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_728_clk_in_regs),
    .D(_04604_),
    .Q(\inst$top.soc.cpu.sink__payload$12[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_334_clk_in_regs),
    .D(_04605_),
    .Q(\inst$top.soc.cpu.sink__payload$12[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_334_clk_in_regs),
    .D(_04606_),
    .Q(\inst$top.soc.cpu.sink__payload$12[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[32]$_SDFFE_PP0P_  (.CLK(clknet_leaf_587_clk_in_regs),
    .D(_04607_),
    .Q(\inst$top.soc.cpu.sink__payload$12[32] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[33]$_SDFFE_PP0P_  (.CLK(clknet_leaf_744_clk_in_regs),
    .D(_04608_),
    .Q(\inst$top.soc.cpu.sink__payload$12[33] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[34]$_SDFFE_PP0P_  (.CLK(clknet_leaf_750_clk_in_regs),
    .D(_04609_),
    .Q(\inst$top.soc.cpu.sink__payload$12[34] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[35]$_SDFFE_PP0P_  (.CLK(clknet_leaf_750_clk_in_regs),
    .D(_04610_),
    .Q(\inst$top.soc.cpu.sink__payload$12[35] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[36]$_SDFFE_PP0P_  (.CLK(clknet_leaf_753_clk_in_regs),
    .D(_04611_),
    .Q(\inst$top.soc.cpu.sink__payload$12[36] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[37]$_SDFFE_PP0P_  (.CLK(clknet_leaf_748_clk_in_regs),
    .D(_04612_),
    .Q(\inst$top.soc.cpu.sink__payload$12[37] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[38]$_SDFFE_PP0P_  (.CLK(clknet_leaf_749_clk_in_regs),
    .D(_04613_),
    .Q(\inst$top.soc.cpu.sink__payload$12[38] ));
 sky130_fd_sc_hd__dfxtp_2 \inst$top.soc.cpu.sink__payload$12[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_727_clk_in_regs),
    .D(_04614_),
    .Q(\inst$top.soc.cpu.sink__payload$12[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_726_clk_in_regs),
    .D(_04615_),
    .Q(\inst$top.soc.cpu.sink__payload$12[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[52]$_SDFFE_PP0P_  (.CLK(clknet_leaf_614_clk_in_regs),
    .D(_04616_),
    .Q(\inst$top.soc.cpu.sink__payload$12[52] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[53]$_SDFFE_PP0P_  (.CLK(clknet_leaf_586_clk_in_regs),
    .D(_04617_),
    .Q(\inst$top.soc.cpu.sink__payload$12[53] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[54]$_SDFFE_PP0P_  (.CLK(clknet_leaf_576_clk_in_regs),
    .D(_04618_),
    .Q(\inst$top.soc.cpu.sink__payload$12[54] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[55]$_SDFFE_PP0P_  (.CLK(clknet_leaf_623_clk_in_regs),
    .D(_04619_),
    .Q(\inst$top.soc.cpu.sink__payload$12[55] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[56]$_SDFFE_PP0P_  (.CLK(clknet_leaf_624_clk_in_regs),
    .D(_04620_),
    .Q(\inst$top.soc.cpu.sink__payload$12[56] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[57]$_SDFFE_PP0P_  (.CLK(clknet_leaf_725_clk_in_regs),
    .D(_04621_),
    .Q(\inst$top.soc.cpu.sink__payload$12[57] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[58]$_SDFFE_PP0P_  (.CLK(clknet_leaf_588_clk_in_regs),
    .D(_04622_),
    .Q(\inst$top.soc.cpu.sink__payload$12[58] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[59]$_SDFFE_PP0P_  (.CLK(clknet_leaf_589_clk_in_regs),
    .D(_04623_),
    .Q(\inst$top.soc.cpu.sink__payload$12[59] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_751_clk_in_regs),
    .D(_04624_),
    .Q(\inst$top.soc.cpu.sink__payload$12[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[60]$_SDFFE_PP0P_  (.CLK(clknet_leaf_588_clk_in_regs),
    .D(_04625_),
    .Q(\inst$top.soc.cpu.sink__payload$12[60] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[61]$_SDFFE_PP0P_  (.CLK(clknet_leaf_591_clk_in_regs),
    .D(_04626_),
    .Q(\inst$top.soc.cpu.sink__payload$12[61] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[62]$_SDFFE_PP0P_  (.CLK(clknet_leaf_587_clk_in_regs),
    .D(_04627_),
    .Q(\inst$top.soc.cpu.sink__payload$12[62] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[63]$_SDFFE_PP0P_  (.CLK(clknet_leaf_729_clk_in_regs),
    .D(_04628_),
    .Q(\inst$top.soc.cpu.sink__payload$12[63] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_744_clk_in_regs),
    .D(_04629_),
    .Q(\inst$top.soc.cpu.sink__payload$12[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_593_clk_in_regs),
    .D(_04630_),
    .Q(\inst$top.soc.cpu.sink__payload$12[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_754_clk_in_regs),
    .D(_04631_),
    .Q(\inst$top.soc.cpu.sink__payload$12[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[95]$_SDFFE_PP0P_  (.CLK(clknet_leaf_588_clk_in_regs),
    .D(_04632_),
    .Q(\inst$top.soc.cpu.d.sink__payload.illegal ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[96]$_SDFFE_PP0P_  (.CLK(clknet_leaf_320_clk_in_regs),
    .D(_04633_),
    .Q(\inst$top.soc.cpu.sink__payload$12[39] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[97]$_SDFFE_PP0P_  (.CLK(clknet_leaf_322_clk_in_regs),
    .D(_04634_),
    .Q(\inst$top.soc.cpu.sink__payload$12[40] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[98]$_SDFFE_PP0P_  (.CLK(clknet_leaf_319_clk_in_regs),
    .D(_04635_),
    .Q(\inst$top.soc.cpu.sink__payload$12[41] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[99]$_SDFFE_PP0P_  (.CLK(clknet_leaf_319_clk_in_regs),
    .D(_04636_),
    .Q(\inst$top.soc.cpu.sink__payload$12[42] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$12[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_596_clk_in_regs),
    .D(_04637_),
    .Q(\inst$top.soc.cpu.sink__payload$12[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[100]$_SDFFE_PP0N_  (.CLK(clknet_leaf_323_clk_in_regs),
    .D(_04638_),
    .Q(\inst$top.soc.cpu.sink__payload$18[100] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[101]$_SDFFE_PP0N_  (.CLK(clknet_leaf_322_clk_in_regs),
    .D(_04639_),
    .Q(\inst$top.soc.cpu.sink__payload$18[101] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[102]$_SDFFE_PP0N_  (.CLK(clknet_leaf_323_clk_in_regs),
    .D(_04640_),
    .Q(\inst$top.soc.cpu.sink__payload$18[102] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[103]$_SDFFE_PP0N_  (.CLK(clknet_leaf_323_clk_in_regs),
    .D(_04641_),
    .Q(\inst$top.soc.cpu.sink__payload$18[103] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[104]$_SDFFE_PP0N_  (.CLK(clknet_leaf_324_clk_in_regs),
    .D(_04642_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.rd_we ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[105]$_SDFFE_PP0N_  (.CLK(clknet_leaf_339_clk_in_regs),
    .D(_04643_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.bypass_m ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[106]$_SDFFE_PP0N_  (.CLK(clknet_leaf_573_clk_in_regs),
    .D(_04644_),
    .Q(\inst$top.soc.cpu.sink__payload$18[106] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[107]$_SDFFE_PP0N_  (.CLK(clknet_6_27__leaf_clk_in_regs),
    .D(_04645_),
    .Q(\inst$top.soc.cpu.sink__payload$18[107] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[108]$_SDFFE_PP0N_  (.CLK(clknet_leaf_318_clk_in_regs),
    .D(_04646_),
    .Q(\inst$top.soc.cpu.sink__payload$18[108] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[109]$_SDFFE_PP0N_  (.CLK(clknet_leaf_579_clk_in_regs),
    .D(_04647_),
    .Q(\inst$top.soc.cpu.sink__payload$18[109] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[10]$_SDFFE_PP0N_  (.CLK(clknet_leaf_598_clk_in_regs),
    .D(_04648_),
    .Q(\inst$top.soc.cpu.sink__payload$18[10] ));
 sky130_fd_sc_hd__dfxtp_2 \inst$top.soc.cpu.sink__payload$18[110]$_SDFFE_PP0N_  (.CLK(clknet_leaf_347_clk_in_regs),
    .D(_04649_),
    .Q(\inst$top.soc.cpu.sink__payload$18[110] ));
 sky130_fd_sc_hd__dfxtp_2 \inst$top.soc.cpu.sink__payload$18[111]$_SDFFE_PP0N_  (.CLK(clknet_leaf_580_clk_in_regs),
    .D(_04650_),
    .Q(\inst$top.soc.cpu.sink__payload$18[111] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[112]$_SDFFE_PP0N_  (.CLK(clknet_leaf_577_clk_in_regs),
    .D(_04651_),
    .Q(\inst$top.soc.cpu.sink__payload$18[112] ));
 sky130_fd_sc_hd__dfxtp_2 \inst$top.soc.cpu.sink__payload$18[113]$_SDFFE_PP0N_  (.CLK(clknet_leaf_345_clk_in_regs),
    .D(_04652_),
    .Q(\inst$top.soc.cpu.sink__payload$18[113] ));
 sky130_fd_sc_hd__dfxtp_2 \inst$top.soc.cpu.sink__payload$18[114]$_SDFFE_PP0N_  (.CLK(clknet_leaf_350_clk_in_regs),
    .D(_04653_),
    .Q(\inst$top.soc.cpu.sink__payload$18[114] ));
 sky130_fd_sc_hd__dfxtp_2 \inst$top.soc.cpu.sink__payload$18[115]$_SDFFE_PP0N_  (.CLK(clknet_leaf_378_clk_in_regs),
    .D(_04654_),
    .Q(\inst$top.soc.cpu.sink__payload$18[115] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[116]$_SDFFE_PP0N_  (.CLK(clknet_leaf_580_clk_in_regs),
    .D(_04655_),
    .Q(\inst$top.soc.cpu.sink__payload$18[116] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[117]$_SDFFE_PP0N_  (.CLK(clknet_leaf_352_clk_in_regs),
    .D(_04656_),
    .Q(\inst$top.soc.cpu.sink__payload$18[117] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[118]$_SDFFE_PP0N_  (.CLK(clknet_leaf_378_clk_in_regs),
    .D(_04657_),
    .Q(\inst$top.soc.cpu.sink__payload$18[118] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[119]$_SDFFE_PP0N_  (.CLK(clknet_leaf_349_clk_in_regs),
    .D(_04658_),
    .Q(\inst$top.soc.cpu.sink__payload$18[119] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[11]$_SDFFE_PP0N_  (.CLK(clknet_leaf_613_clk_in_regs),
    .D(_04659_),
    .Q(\inst$top.soc.cpu.sink__payload$18[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[120]$_SDFFE_PP0N_  (.CLK(clknet_leaf_348_clk_in_regs),
    .D(_04660_),
    .Q(\inst$top.soc.cpu.sink__payload$18[120] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[121]$_SDFFE_PP0N_  (.CLK(clknet_6_44__leaf_clk_in_regs),
    .D(_04661_),
    .Q(\inst$top.soc.cpu.sink__payload$18[121] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[122]$_SDFFE_PP0N_  (.CLK(clknet_leaf_578_clk_in_regs),
    .D(_04662_),
    .Q(\inst$top.soc.cpu.sink__payload$18[122] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[123]$_SDFFE_PP0N_  (.CLK(clknet_leaf_359_clk_in_regs),
    .D(_04663_),
    .Q(\inst$top.soc.cpu.sink__payload$18[123] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[124]$_SDFFE_PP0N_  (.CLK(clknet_leaf_350_clk_in_regs),
    .D(_04664_),
    .Q(\inst$top.soc.cpu.sink__payload$18[124] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[125]$_SDFFE_PP0N_  (.CLK(clknet_leaf_577_clk_in_regs),
    .D(_04665_),
    .Q(\inst$top.soc.cpu.sink__payload$18[125] ));
 sky130_fd_sc_hd__dfxtp_2 \inst$top.soc.cpu.sink__payload$18[126]$_SDFFE_PP0N_  (.CLK(clknet_leaf_376_clk_in_regs),
    .D(_04666_),
    .Q(\inst$top.soc.cpu.sink__payload$18[126] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[127]$_SDFFE_PP0N_  (.CLK(clknet_leaf_574_clk_in_regs),
    .D(_04667_),
    .Q(\inst$top.soc.cpu.sink__payload$18[127] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[128]$_SDFFE_PP0N_  (.CLK(clknet_leaf_575_clk_in_regs),
    .D(_04668_),
    .Q(\inst$top.soc.cpu.sink__payload$18[128] ));
 sky130_fd_sc_hd__dfxtp_2 \inst$top.soc.cpu.sink__payload$18[129]$_SDFFE_PP0N_  (.CLK(clknet_leaf_562_clk_in_regs),
    .D(_04669_),
    .Q(\inst$top.soc.cpu.sink__payload$18[129] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[12]$_SDFFE_PP0N_  (.CLK(clknet_leaf_610_clk_in_regs),
    .D(_04670_),
    .Q(\inst$top.soc.cpu.sink__payload$18[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[130]$_SDFFE_PP0N_  (.CLK(clknet_leaf_577_clk_in_regs),
    .D(_04671_),
    .Q(\inst$top.soc.cpu.sink__payload$18[130] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[131]$_SDFFE_PP0N_  (.CLK(clknet_leaf_385_clk_in_regs),
    .D(_04672_),
    .Q(\inst$top.soc.cpu.sink__payload$18[131] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[132]$_SDFFE_PP0N_  (.CLK(clknet_leaf_576_clk_in_regs),
    .D(_04673_),
    .Q(\inst$top.soc.cpu.sink__payload$18[132] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[133]$_SDFFE_PP0N_  (.CLK(clknet_leaf_562_clk_in_regs),
    .D(_04674_),
    .Q(\inst$top.soc.cpu.sink__payload$18[133] ));
 sky130_fd_sc_hd__dfxtp_2 \inst$top.soc.cpu.sink__payload$18[134]$_SDFFE_PP0N_  (.CLK(clknet_leaf_562_clk_in_regs),
    .D(_04675_),
    .Q(\inst$top.soc.cpu.sink__payload$18[134] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[135]$_SDFFE_PP0N_  (.CLK(clknet_leaf_574_clk_in_regs),
    .D(_04676_),
    .Q(\inst$top.soc.cpu.sink__payload$18[135] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[136]$_SDFFE_PP0N_  (.CLK(clknet_leaf_575_clk_in_regs),
    .D(_04677_),
    .Q(\inst$top.soc.cpu.sink__payload$18[136] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[137]$_SDFFE_PP0N_  (.CLK(clknet_leaf_384_clk_in_regs),
    .D(_04678_),
    .Q(\inst$top.soc.cpu.sink__payload$18[137] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[138]$_SDFFE_PP0N_  (.CLK(clknet_leaf_576_clk_in_regs),
    .D(_04679_),
    .Q(\inst$top.soc.cpu.sink__payload$18[138] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[139]$_SDFFE_PP0N_  (.CLK(clknet_leaf_579_clk_in_regs),
    .D(_04680_),
    .Q(\inst$top.soc.cpu.sink__payload$18[139] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[13]$_SDFFE_PP0N_  (.CLK(clknet_leaf_603_clk_in_regs),
    .D(_04681_),
    .Q(\inst$top.soc.cpu.sink__payload$18[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[140]$_SDFFE_PP0N_  (.CLK(clknet_leaf_344_clk_in_regs),
    .D(_04682_),
    .Q(\inst$top.soc.cpu.sink__payload$18[140] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[141]$_SDFFE_PP0N_  (.CLK(clknet_leaf_580_clk_in_regs),
    .D(_04683_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.shift ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[142]$_SDFFE_PP0N_  (.CLK(clknet_leaf_586_clk_in_regs),
    .D(_04684_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.load ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[143]$_SDFFE_PP0N_  (.CLK(clknet_leaf_334_clk_in_regs),
    .D(_04685_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.store ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[14]$_SDFFE_PP0N_  (.CLK(clknet_leaf_595_clk_in_regs),
    .D(_04686_),
    .Q(\inst$top.soc.cpu.sink__payload$18[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[15]$_SDFFE_PP0N_  (.CLK(clknet_leaf_599_clk_in_regs),
    .D(_04687_),
    .Q(\inst$top.soc.cpu.sink__payload$18[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[16]$_SDFFE_PP0N_  (.CLK(clknet_leaf_614_clk_in_regs),
    .D(_04688_),
    .Q(\inst$top.soc.cpu.sink__payload$18[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[176]$_SDFFE_PP0N_  (.CLK(clknet_leaf_573_clk_in_regs),
    .D(_04689_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.compare ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[177]$_SDFFE_PP0N_  (.CLK(clknet_leaf_340_clk_in_regs),
    .D(_04690_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.multiply ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[178]$_SDFFE_PP0N_  (.CLK(clknet_6_31__leaf_clk_in_regs),
    .D(_04691_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.divide ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[179]$_SDFFE_PP0N_  (.CLK(clknet_leaf_579_clk_in_regs),
    .D(_04692_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.condition_met ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[17]$_SDFFE_PP0N_  (.CLK(clknet_leaf_611_clk_in_regs),
    .D(_04693_),
    .Q(\inst$top.soc.cpu.sink__payload$18[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[180]$_SDFFE_PP0N_  (.CLK(clknet_leaf_746_clk_in_regs),
    .D(_04694_),
    .Q(\inst$top.soc.cpu.sink__payload$18[180] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[181]$_SDFFE_PP0N_  (.CLK(clknet_leaf_587_clk_in_regs),
    .D(_04695_),
    .Q(\inst$top.soc.cpu.sink__payload$18[181] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[182]$_SDFFE_PP0N_  (.CLK(clknet_leaf_730_clk_in_regs),
    .D(_04696_),
    .Q(\inst$top.soc.cpu.sink__payload$18[182] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[183]$_SDFFE_PP0N_  (.CLK(clknet_leaf_730_clk_in_regs),
    .D(_04697_),
    .Q(\inst$top.soc.cpu.sink__payload$18[183] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[184]$_SDFFE_PP0N_  (.CLK(clknet_leaf_729_clk_in_regs),
    .D(_04698_),
    .Q(\inst$top.soc.cpu.sink__payload$18[184] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[185]$_SDFFE_PP0N_  (.CLK(clknet_leaf_748_clk_in_regs),
    .D(_04699_),
    .Q(\inst$top.soc.cpu.sink__payload$18[185] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[186]$_SDFFE_PP0N_  (.CLK(clknet_leaf_749_clk_in_regs),
    .D(_04700_),
    .Q(\inst$top.soc.cpu.sink__payload$18[186] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[187]$_SDFFE_PP0N_  (.CLK(clknet_leaf_726_clk_in_regs),
    .D(_04701_),
    .Q(\inst$top.soc.cpu.sink__payload$18[187] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[188]$_SDFFE_PP0N_  (.CLK(clknet_leaf_754_clk_in_regs),
    .D(_04702_),
    .Q(\inst$top.soc.cpu.sink__payload$18[188] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[189]$_SDFFE_PP0N_  (.CLK(clknet_leaf_754_clk_in_regs),
    .D(_04703_),
    .Q(\inst$top.soc.cpu.sink__payload$18[189] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[18]$_SDFFE_PP0N_  (.CLK(clknet_leaf_649_clk_in_regs),
    .D(_04704_),
    .Q(\inst$top.soc.cpu.sink__payload$18[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[190]$_SDFFE_PP0N_  (.CLK(clknet_leaf_594_clk_in_regs),
    .D(_04705_),
    .Q(\inst$top.soc.cpu.sink__payload$18[190] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[191]$_SDFFE_PP0N_  (.CLK(clknet_leaf_749_clk_in_regs),
    .D(_04706_),
    .Q(\inst$top.soc.cpu.sink__payload$18[191] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[192]$_SDFFE_PP0N_  (.CLK(clknet_leaf_744_clk_in_regs),
    .D(_04707_),
    .Q(\inst$top.soc.cpu.sink__payload$18[192] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[193]$_SDFFE_PP0N_  (.CLK(clknet_leaf_595_clk_in_regs),
    .D(_04708_),
    .Q(\inst$top.soc.cpu.sink__payload$18[193] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[194]$_SDFFE_PP0N_  (.CLK(clknet_leaf_596_clk_in_regs),
    .D(_04709_),
    .Q(\inst$top.soc.cpu.sink__payload$18[194] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[195]$_SDFFE_PP0N_  (.CLK(clknet_leaf_593_clk_in_regs),
    .D(_04710_),
    .Q(\inst$top.soc.cpu.sink__payload$18[195] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[196]$_SDFFE_PP0N_  (.CLK(clknet_leaf_743_clk_in_regs),
    .D(_04711_),
    .Q(\inst$top.soc.cpu.sink__payload$18[196] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[197]$_SDFFE_PP0N_  (.CLK(clknet_leaf_754_clk_in_regs),
    .D(_04712_),
    .Q(\inst$top.soc.cpu.sink__payload$18[197] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[198]$_SDFFE_PP0N_  (.CLK(clknet_leaf_744_clk_in_regs),
    .D(_04713_),
    .Q(\inst$top.soc.cpu.sink__payload$18[198] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[199]$_SDFFE_PP0N_  (.CLK(clknet_leaf_751_clk_in_regs),
    .D(_04714_),
    .Q(\inst$top.soc.cpu.sink__payload$18[199] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[19]$_SDFFE_PP0N_  (.CLK(clknet_leaf_614_clk_in_regs),
    .D(_04715_),
    .Q(\inst$top.soc.cpu.sink__payload$18[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[200]$_SDFFE_PP0N_  (.CLK(clknet_leaf_748_clk_in_regs),
    .D(_04716_),
    .Q(\inst$top.soc.cpu.sink__payload$18[200] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[201]$_SDFFE_PP0N_  (.CLK(clknet_leaf_744_clk_in_regs),
    .D(_04717_),
    .Q(\inst$top.soc.cpu.sink__payload$18[201] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[202]$_SDFFE_PP0N_  (.CLK(clknet_leaf_594_clk_in_regs),
    .D(_04718_),
    .Q(\inst$top.soc.cpu.sink__payload$18[202] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[203]$_SDFFE_PP0N_  (.CLK(clknet_leaf_594_clk_in_regs),
    .D(_04719_),
    .Q(\inst$top.soc.cpu.sink__payload$18[203] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[204]$_SDFFE_PP0N_  (.CLK(clknet_leaf_593_clk_in_regs),
    .D(_04720_),
    .Q(\inst$top.soc.cpu.sink__payload$18[204] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[205]$_SDFFE_PP0N_  (.CLK(clknet_leaf_726_clk_in_regs),
    .D(_04721_),
    .Q(\inst$top.soc.cpu.sink__payload$18[205] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[206]$_SDFFE_PP0N_  (.CLK(clknet_leaf_590_clk_in_regs),
    .D(_04722_),
    .Q(\inst$top.soc.cpu.sink__payload$18[206] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[207]$_SDFFE_PP0N_  (.CLK(clknet_leaf_591_clk_in_regs),
    .D(_04723_),
    .Q(\inst$top.soc.cpu.sink__payload$18[207] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[208]$_SDFFE_PP0N_  (.CLK(clknet_leaf_589_clk_in_regs),
    .D(_04724_),
    .Q(\inst$top.soc.cpu.sink__payload$18[208] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[209]$_SDFFE_PP0N_  (.CLK(clknet_leaf_590_clk_in_regs),
    .D(_04725_),
    .Q(\inst$top.soc.cpu.sink__payload$18[209] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[20]$_SDFFE_PP0N_  (.CLK(clknet_leaf_650_clk_in_regs),
    .D(_04726_),
    .Q(\inst$top.soc.cpu.sink__payload$18[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[210]$_SDFFE_PP0N_  (.CLK(clknet_leaf_590_clk_in_regs),
    .D(_04727_),
    .Q(\inst$top.soc.cpu.sink__payload$18[210] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[211]$_SDFFE_PP0N_  (.CLK(clknet_leaf_726_clk_in_regs),
    .D(_04728_),
    .Q(\inst$top.soc.cpu.sink__payload$18[211] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[212]$_SDFFE_PP0N_  (.CLK(clknet_leaf_585_clk_in_regs),
    .D(_04729_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.branch_taken ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[213]$_SDFFE_PP0N_  (.CLK(clknet_leaf_746_clk_in_regs),
    .D(_04730_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.branch_predict_taken ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[214]$_SDFFE_PP0N_  (.CLK(clknet_leaf_757_clk_in_regs),
    .D(_04731_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.csr_we ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[215]$_SDFFE_PP0N_  (.CLK(clknet_leaf_568_clk_in_regs),
    .D(_04732_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[216]$_SDFFE_PP0N_  (.CLK(clknet_leaf_568_clk_in_regs),
    .D(_04733_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[217]$_SDFFE_PP0N_  (.CLK(clknet_leaf_720_clk_in_regs),
    .D(_04734_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[218]$_SDFFE_PP0N_  (.CLK(clknet_leaf_720_clk_in_regs),
    .D(_04735_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[219]$_SDFFE_PP0N_  (.CLK(clknet_leaf_601_clk_in_regs),
    .D(_04736_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[21]$_SDFFE_PP0N_  (.CLK(clknet_leaf_613_clk_in_regs),
    .D(_04737_),
    .Q(\inst$top.soc.cpu.sink__payload$18[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[220]$_SDFFE_PP0N_  (.CLK(clknet_leaf_584_clk_in_regs),
    .D(_04738_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[221]$_SDFFE_PP0N_  (.CLK(clknet_6_31__leaf_clk_in_regs),
    .D(_04739_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[222]$_SDFFE_PP0N_  (.CLK(clknet_leaf_628_clk_in_regs),
    .D(_04740_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[223]$_SDFFE_PP0N_  (.CLK(clknet_leaf_584_clk_in_regs),
    .D(_04741_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[224]$_SDFFE_PP0N_  (.CLK(clknet_leaf_600_clk_in_regs),
    .D(_04742_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[225]$_SDFFE_PP0N_  (.CLK(clknet_leaf_572_clk_in_regs),
    .D(_04743_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[226]$_SDFFE_PP0N_  (.CLK(clknet_leaf_572_clk_in_regs),
    .D(_04744_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[227]$_SDFFE_PP0N_  (.CLK(clknet_leaf_602_clk_in_regs),
    .D(_04745_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[228]$_SDFFE_PP0N_  (.CLK(clknet_6_30__leaf_clk_in_regs),
    .D(_04746_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[229]$_SDFFE_PP0N_  (.CLK(clknet_leaf_602_clk_in_regs),
    .D(_04747_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[22]$_SDFFE_PP0N_  (.CLK(clknet_leaf_619_clk_in_regs),
    .D(_04748_),
    .Q(\inst$top.soc.cpu.sink__payload$18[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[230]$_SDFFE_PP0N_  (.CLK(clknet_leaf_598_clk_in_regs),
    .D(_04749_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[231]$_SDFFE_PP0N_  (.CLK(clknet_leaf_567_clk_in_regs),
    .D(_04750_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[232]$_SDFFE_PP0N_  (.CLK(clknet_leaf_567_clk_in_regs),
    .D(_04751_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[233]$_SDFFE_PP0N_  (.CLK(clknet_leaf_566_clk_in_regs),
    .D(_04752_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[234]$_SDFFE_PP0N_  (.CLK(clknet_leaf_633_clk_in_regs),
    .D(_04753_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[235]$_SDFFE_PP0N_  (.CLK(clknet_leaf_633_clk_in_regs),
    .D(_04754_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[236]$_SDFFE_PP0N_  (.CLK(clknet_6_31__leaf_clk_in_regs),
    .D(_04755_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[237]$_SDFFE_PP0N_  (.CLK(clknet_leaf_565_clk_in_regs),
    .D(_04756_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[238]$_SDFFE_PP0N_  (.CLK(clknet_leaf_566_clk_in_regs),
    .D(_04757_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[239]$_SDFFE_PP0N_  (.CLK(clknet_leaf_570_clk_in_regs),
    .D(_04758_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[23]$_SDFFE_PP0N_  (.CLK(clknet_leaf_622_clk_in_regs),
    .D(_04759_),
    .Q(\inst$top.soc.cpu.sink__payload$18[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[240]$_SDFFE_PP0N_  (.CLK(clknet_leaf_565_clk_in_regs),
    .D(_04760_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[241]$_SDFFE_PP0N_  (.CLK(clknet_leaf_565_clk_in_regs),
    .D(_04761_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[242]$_SDFFE_PP0N_  (.CLK(clknet_leaf_632_clk_in_regs),
    .D(_04762_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[243]$_SDFFE_PP0N_  (.CLK(clknet_leaf_564_clk_in_regs),
    .D(_04763_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[244]$_SDFFE_PP0N_  (.CLK(clknet_leaf_570_clk_in_regs),
    .D(_04764_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[245]$_SDFFE_PP0N_  (.CLK(clknet_leaf_632_clk_in_regs),
    .D(_04765_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[246]$_SDFFE_PP0N_  (.CLK(clknet_leaf_635_clk_in_regs),
    .D(_04766_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__m_wp_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[247]$_SDFFE_PP0N_  (.CLK(clknet_leaf_593_clk_in_regs),
    .D(_04767_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.mret ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[24]$_SDFFE_PP0N_  (.CLK(clknet_leaf_625_clk_in_regs),
    .D(_04768_),
    .Q(\inst$top.soc.cpu.sink__payload$18[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[25]$_SDFFE_PP0N_  (.CLK(clknet_leaf_718_clk_in_regs),
    .D(_04769_),
    .Q(\inst$top.soc.cpu.sink__payload$18[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[26]$_SDFFE_PP0N_  (.CLK(clknet_leaf_626_clk_in_regs),
    .D(_04770_),
    .Q(\inst$top.soc.cpu.sink__payload$18[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[27]$_SDFFE_PP0N_  (.CLK(clknet_leaf_625_clk_in_regs),
    .D(_04771_),
    .Q(\inst$top.soc.cpu.sink__payload$18[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[28]$_SDFFE_PP0N_  (.CLK(clknet_leaf_624_clk_in_regs),
    .D(_04772_),
    .Q(\inst$top.soc.cpu.sink__payload$18[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[29]$_SDFFE_PP0N_  (.CLK(clknet_leaf_623_clk_in_regs),
    .D(_04773_),
    .Q(\inst$top.soc.cpu.sink__payload$18[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_730_clk_in_regs),
    .D(_04774_),
    .Q(\inst$top.soc.cpu.sink__payload$18[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[30]$_SDFFE_PP0N_  (.CLK(clknet_leaf_602_clk_in_regs),
    .D(_04775_),
    .Q(\inst$top.soc.cpu.sink__payload$18[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[31]$_SDFFE_PP0N_  (.CLK(clknet_leaf_732_clk_in_regs),
    .D(_04776_),
    .Q(\inst$top.soc.cpu.sink__payload$18[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[32]$_SDFFE_PP0N_  (.CLK(clknet_leaf_743_clk_in_regs),
    .D(_04777_),
    .Q(\inst$top.soc.cpu.sink__payload$18[32] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[33]$_SDFFE_PP0N_  (.CLK(clknet_leaf_743_clk_in_regs),
    .D(_04778_),
    .Q(\inst$top.soc.cpu.sink__payload$18[33] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[34]$_SDFFE_PP0N_  (.CLK(clknet_leaf_728_clk_in_regs),
    .D(_04779_),
    .Q(\inst$top.soc.cpu.sink__payload$18[34] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[35]$_SDFFE_PP0N_  (.CLK(clknet_leaf_749_clk_in_regs),
    .D(_04780_),
    .Q(\inst$top.soc.cpu.sink__payload$18[35] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[36]$_SDFFE_PP0N_  (.CLK(clknet_leaf_731_clk_in_regs),
    .D(_04781_),
    .Q(\inst$top.soc.cpu.sink__payload$18[36] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[37]$_SDFFE_PP0N_  (.CLK(clknet_leaf_744_clk_in_regs),
    .D(_04782_),
    .Q(\inst$top.soc.cpu.sink__payload$18[37] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[38]$_SDFFE_PP0N_  (.CLK(clknet_leaf_746_clk_in_regs),
    .D(_04783_),
    .Q(\inst$top.soc.cpu.sink__payload$18[38] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_736_clk_in_regs),
    .D(_04784_),
    .Q(\inst$top.soc.cpu.sink__payload$18[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[47]$_SDFFE_PP0N_  (.CLK(clknet_leaf_342_clk_in_regs),
    .D(_04785_),
    .Q(\inst$top.soc.cpu.sink__payload$18[47] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[48]$_SDFFE_PP0N_  (.CLK(clknet_leaf_742_clk_in_regs),
    .D(_04786_),
    .Q(\inst$top.soc.cpu.sink__payload$18[48] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[49]$_SDFFE_PP0N_  (.CLK(clknet_leaf_578_clk_in_regs),
    .D(_04787_),
    .Q(\inst$top.soc.cpu.sink__payload$18[49] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_731_clk_in_regs),
    .D(_04788_),
    .Q(\inst$top.soc.cpu.sink__payload$18[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[50]$_SDFFE_PP0N_  (.CLK(clknet_leaf_578_clk_in_regs),
    .D(_04789_),
    .Q(\inst$top.soc.cpu.sink__payload$18[50] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[51]$_SDFFE_PP0N_  (.CLK(clknet_leaf_578_clk_in_regs),
    .D(_04790_),
    .Q(\inst$top.soc.cpu.sink__payload$18[51] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[52]$_SDFFE_PP0N_  (.CLK(clknet_leaf_651_clk_in_regs),
    .D(_04791_),
    .Q(\inst$top.soc.cpu.sink__payload$18[52] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[53]$_SDFFE_PP0N_  (.CLK(clknet_leaf_586_clk_in_regs),
    .D(_04792_),
    .Q(\inst$top.soc.cpu.sink__payload$18[53] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[54]$_SDFFE_PP0N_  (.CLK(clknet_leaf_624_clk_in_regs),
    .D(_04793_),
    .Q(\inst$top.soc.cpu.sink__payload$18[54] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[55]$_SDFFE_PP0N_  (.CLK(clknet_leaf_623_clk_in_regs),
    .D(_04794_),
    .Q(\inst$top.soc.cpu.sink__payload$18[55] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[56]$_SDFFE_PP0N_  (.CLK(clknet_leaf_624_clk_in_regs),
    .D(_04795_),
    .Q(\inst$top.soc.cpu.sink__payload$18[56] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[57]$_SDFFE_PP0N_  (.CLK(clknet_leaf_725_clk_in_regs),
    .D(_04796_),
    .Q(\inst$top.soc.cpu.sink__payload$18[57] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[58]$_SDFFE_PP0N_  (.CLK(clknet_leaf_587_clk_in_regs),
    .D(_04797_),
    .Q(\inst$top.soc.cpu.sink__payload$18[58] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[59]$_SDFFE_PP0N_  (.CLK(clknet_leaf_591_clk_in_regs),
    .D(_04798_),
    .Q(\inst$top.soc.cpu.sink__payload$18[59] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_745_clk_in_regs),
    .D(_04799_),
    .Q(\inst$top.soc.cpu.sink__payload$18[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[60]$_SDFFE_PP0N_  (.CLK(clknet_leaf_592_clk_in_regs),
    .D(_04800_),
    .Q(\inst$top.soc.cpu.sink__payload$18[60] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[61]$_SDFFE_PP0N_  (.CLK(clknet_leaf_592_clk_in_regs),
    .D(_04801_),
    .Q(\inst$top.soc.cpu.sink__payload$18[61] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[62]$_SDFFE_PP0N_  (.CLK(clknet_leaf_602_clk_in_regs),
    .D(_04802_),
    .Q(\inst$top.soc.cpu.sink__payload$18[62] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[63]$_SDFFE_PP0N_  (.CLK(clknet_leaf_731_clk_in_regs),
    .D(_04803_),
    .Q(\inst$top.soc.cpu.sink__payload$18[63] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[6]$_SDFFE_PP0N_  (.CLK(clknet_leaf_741_clk_in_regs),
    .D(_04804_),
    .Q(\inst$top.soc.cpu.sink__payload$18[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[7]$_SDFFE_PP0N_  (.CLK(clknet_leaf_724_clk_in_regs),
    .D(_04805_),
    .Q(\inst$top.soc.cpu.sink__payload$18[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[8]$_SDFFE_PP0N_  (.CLK(clknet_leaf_754_clk_in_regs),
    .D(_04806_),
    .Q(\inst$top.soc.cpu.sink__payload$18[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[95]$_SDFFE_PP0N_  (.CLK(clknet_leaf_745_clk_in_regs),
    .D(_04807_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.illegal ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[96]$_SDFFE_PP0N_  (.CLK(clknet_leaf_585_clk_in_regs),
    .D(_04808_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.loadstore_misaligned ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[97]$_SDFFE_PP0N_  (.CLK(clknet_leaf_586_clk_in_regs),
    .D(_04809_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.ecall ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[98]$_SDFFE_PP0N_  (.CLK(clknet_leaf_748_clk_in_regs),
    .D(_04810_),
    .Q(\inst$top.soc.cpu.d.sink__payload$6.ebreak ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[99]$_SDFFE_PP0N_  (.CLK(clknet_leaf_321_clk_in_regs),
    .D(_04811_),
    .Q(\inst$top.soc.cpu.sink__payload$18[39] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$18[9]$_SDFFE_PP0N_  (.CLK(clknet_leaf_743_clk_in_regs),
    .D(_04812_),
    .Q(\inst$top.soc.cpu.sink__payload$18[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[100]$_SDFFE_PP0N_  (.CLK(clknet_leaf_309_clk_in_regs),
    .D(_04813_),
    .Q(\inst$top.soc.cpu.sink__payload$24[100] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[101]$_SDFFE_PP0N_  (.CLK(clknet_leaf_317_clk_in_regs),
    .D(_04814_),
    .Q(\inst$top.soc.cpu.sink__payload$24[101] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[102]$_SDFFE_PP0N_  (.CLK(clknet_leaf_316_clk_in_regs),
    .D(_04815_),
    .Q(\inst$top.soc.cpu.sink__payload$24[102] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[103]$_SDFFE_PP0N_  (.CLK(clknet_leaf_276_clk_in_regs),
    .D(_04816_),
    .Q(\inst$top.soc.cpu.sink__payload$24[103] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[104]$_SDFFE_PP0N_  (.CLK(clknet_leaf_308_clk_in_regs),
    .D(_04817_),
    .Q(\inst$top.soc.cpu.sink__payload$24[104] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[105]$_SDFFE_PP0N_  (.CLK(clknet_leaf_314_clk_in_regs),
    .D(_04818_),
    .Q(\inst$top.soc.cpu.sink__payload$24[105] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[106]$_SDFFE_PP0N_  (.CLK(clknet_leaf_757_clk_in_regs),
    .D(_04819_),
    .Q(\inst$top.soc.cpu.d.sink__payload$16.csr_we ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[107]$_SDFFE_PP0N_  (.CLK(clknet_leaf_717_clk_in_regs),
    .D(_04820_),
    .Q(\inst$top.soc.cpu.d.sink__payload$16.csr_rdy ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[108]$_SDFFE_PP0N_  (.CLK(clknet_leaf_564_clk_in_regs),
    .D(_04821_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[109]$_SDFFE_PP0N_  (.CLK(clknet_leaf_662_clk_in_regs),
    .D(_04822_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[10]$_SDFFE_PP0N_  (.CLK(clknet_leaf_606_clk_in_regs),
    .D(_04823_),
    .Q(\inst$top.soc.cpu.sink__payload$24[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[110]$_SDFFE_PP0N_  (.CLK(clknet_leaf_737_clk_in_regs),
    .D(_04824_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[111]$_SDFFE_PP0N_  (.CLK(clknet_leaf_719_clk_in_regs),
    .D(_04825_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[112]$_SDFFE_PP0N_  (.CLK(clknet_leaf_721_clk_in_regs),
    .D(_04826_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[113]$_SDFFE_PP0N_  (.CLK(clknet_leaf_599_clk_in_regs),
    .D(_04827_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[114]$_SDFFE_PP0N_  (.CLK(clknet_leaf_613_clk_in_regs),
    .D(_04828_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[115]$_SDFFE_PP0N_  (.CLK(clknet_leaf_657_clk_in_regs),
    .D(_04829_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[116]$_SDFFE_PP0N_  (.CLK(clknet_leaf_600_clk_in_regs),
    .D(_04830_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[117]$_SDFFE_PP0N_  (.CLK(clknet_leaf_597_clk_in_regs),
    .D(_04831_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[118]$_SDFFE_PP0N_  (.CLK(clknet_leaf_621_clk_in_regs),
    .D(_04832_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[119]$_SDFFE_PP0N_  (.CLK(clknet_leaf_614_clk_in_regs),
    .D(_04833_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[11]$_SDFFE_PP0N_  (.CLK(clknet_leaf_738_clk_in_regs),
    .D(_04834_),
    .Q(\inst$top.soc.cpu.sink__payload$24[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[120]$_SDFFE_PP0N_  (.CLK(clknet_leaf_603_clk_in_regs),
    .D(_04835_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[121]$_SDFFE_PP0N_  (.CLK(clknet_leaf_624_clk_in_regs),
    .D(_04836_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[122]$_SDFFE_PP0N_  (.CLK(clknet_leaf_601_clk_in_regs),
    .D(_04837_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[123]$_SDFFE_PP0N_  (.CLK(clknet_leaf_598_clk_in_regs),
    .D(_04838_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[124]$_SDFFE_PP0N_  (.CLK(clknet_6_29__leaf_clk_in_regs),
    .D(_04839_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[125]$_SDFFE_PP0N_  (.CLK(clknet_leaf_632_clk_in_regs),
    .D(_04840_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[126]$_SDFFE_PP0N_  (.CLK(clknet_leaf_685_clk_in_regs),
    .D(_04841_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[127]$_SDFFE_PP0N_  (.CLK(clknet_leaf_634_clk_in_regs),
    .D(_04842_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[128]$_SDFFE_PP0N_  (.CLK(clknet_leaf_634_clk_in_regs),
    .D(_04843_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[129]$_SDFFE_PP0N_  (.CLK(clknet_leaf_626_clk_in_regs),
    .D(_04844_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[12]$_SDFFE_PP0N_  (.CLK(clknet_leaf_612_clk_in_regs),
    .D(_04845_),
    .Q(\inst$top.soc.cpu.sink__payload$24[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[130]$_SDFFE_PP0N_  (.CLK(clknet_leaf_685_clk_in_regs),
    .D(_04846_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[131]$_SDFFE_PP0N_  (.CLK(clknet_leaf_634_clk_in_regs),
    .D(_04847_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[132]$_SDFFE_PP0N_  (.CLK(clknet_leaf_627_clk_in_regs),
    .D(_04848_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[133]$_SDFFE_PP0N_  (.CLK(clknet_leaf_669_clk_in_regs),
    .D(_04849_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[134]$_SDFFE_PP0N_  (.CLK(clknet_leaf_686_clk_in_regs),
    .D(_04850_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[135]$_SDFFE_PP0N_  (.CLK(clknet_leaf_632_clk_in_regs),
    .D(_04851_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[136]$_SDFFE_PP0N_  (.CLK(clknet_leaf_630_clk_in_regs),
    .D(_04852_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[137]$_SDFFE_PP0N_  (.CLK(clknet_leaf_626_clk_in_regs),
    .D(_04853_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[138]$_SDFFE_PP0N_  (.CLK(clknet_leaf_633_clk_in_regs),
    .D(_04854_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[139]$_SDFFE_PP0N_  (.CLK(clknet_leaf_669_clk_in_regs),
    .D(_04855_),
    .Q(\inst$top.soc.cpu.exception.csr_bank.mcause.port__w_wp_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[13]$_SDFFE_PP0N_  (.CLK(clknet_leaf_603_clk_in_regs),
    .D(_04856_),
    .Q(\inst$top.soc.cpu.sink__payload$24[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[140]$_SDFFE_PP0N_  (.CLK(clknet_leaf_341_clk_in_regs),
    .D(_04857_),
    .Q(\inst$top.soc.cpu.d.sink__payload$16.multiply ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[14]$_SDFFE_PP0N_  (.CLK(clknet_leaf_596_clk_in_regs),
    .D(_04858_),
    .Q(\inst$top.soc.cpu.sink__payload$24[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[15]$_SDFFE_PP0N_  (.CLK(clknet_leaf_595_clk_in_regs),
    .D(_04859_),
    .Q(\inst$top.soc.cpu.sink__payload$24[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[16]$_SDFFE_PP0N_  (.CLK(clknet_leaf_653_clk_in_regs),
    .D(_04860_),
    .Q(\inst$top.soc.cpu.sink__payload$24[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[17]$_SDFFE_PP0N_  (.CLK(clknet_leaf_648_clk_in_regs),
    .D(_04861_),
    .Q(\inst$top.soc.cpu.sink__payload$24[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[18]$_SDFFE_PP0N_  (.CLK(clknet_leaf_649_clk_in_regs),
    .D(_04862_),
    .Q(\inst$top.soc.cpu.sink__payload$24[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[19]$_SDFFE_PP0N_  (.CLK(clknet_leaf_649_clk_in_regs),
    .D(_04863_),
    .Q(\inst$top.soc.cpu.sink__payload$24[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[20]$_SDFFE_PP0N_  (.CLK(clknet_leaf_646_clk_in_regs),
    .D(_04864_),
    .Q(\inst$top.soc.cpu.sink__payload$24[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[21]$_SDFFE_PP0N_  (.CLK(clknet_leaf_613_clk_in_regs),
    .D(_04865_),
    .Q(\inst$top.soc.cpu.sink__payload$24[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[22]$_SDFFE_PP0N_  (.CLK(clknet_leaf_629_clk_in_regs),
    .D(_04866_),
    .Q(\inst$top.soc.cpu.sink__payload$24[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[23]$_SDFFE_PP0N_  (.CLK(clknet_leaf_629_clk_in_regs),
    .D(_04867_),
    .Q(\inst$top.soc.cpu.sink__payload$24[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[24]$_SDFFE_PP0N_  (.CLK(clknet_leaf_625_clk_in_regs),
    .D(_04868_),
    .Q(\inst$top.soc.cpu.sink__payload$24[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[25]$_SDFFE_PP0N_  (.CLK(clknet_leaf_660_clk_in_regs),
    .D(_04869_),
    .Q(\inst$top.soc.cpu.sink__payload$24[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[26]$_SDFFE_PP0N_  (.CLK(clknet_leaf_630_clk_in_regs),
    .D(_04870_),
    .Q(\inst$top.soc.cpu.sink__payload$24[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[27]$_SDFFE_PP0N_  (.CLK(clknet_leaf_627_clk_in_regs),
    .D(_04871_),
    .Q(\inst$top.soc.cpu.sink__payload$24[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[28]$_SDFFE_PP0N_  (.CLK(clknet_leaf_627_clk_in_regs),
    .D(_04872_),
    .Q(\inst$top.soc.cpu.sink__payload$24[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[29]$_SDFFE_PP0N_  (.CLK(clknet_leaf_622_clk_in_regs),
    .D(_04873_),
    .Q(\inst$top.soc.cpu.sink__payload$24[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_730_clk_in_regs),
    .D(_04874_),
    .Q(\inst$top.soc.cpu.sink__payload$24[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[30]$_SDFFE_PP0N_  (.CLK(clknet_leaf_623_clk_in_regs),
    .D(_04875_),
    .Q(\inst$top.soc.cpu.sink__payload$24[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[31]$_SDFFE_PP0N_  (.CLK(clknet_leaf_732_clk_in_regs),
    .D(_04876_),
    .Q(\inst$top.soc.cpu.sink__payload$24[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[32]$_SDFFE_PP0N_  (.CLK(clknet_leaf_296_clk_in_regs),
    .D(_04877_),
    .Q(\inst$top.soc.cpu.sink__payload$24[32] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[33]$_SDFFE_PP0N_  (.CLK(clknet_leaf_296_clk_in_regs),
    .D(_04878_),
    .Q(\inst$top.soc.cpu.sink__payload$24[33] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[34]$_SDFFE_PP0N_  (.CLK(clknet_6_41__leaf_clk_in_regs),
    .D(_04879_),
    .Q(\inst$top.soc.cpu.sink__payload$24[34] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[35]$_SDFFE_PP0N_  (.CLK(clknet_leaf_296_clk_in_regs),
    .D(_04880_),
    .Q(\inst$top.soc.cpu.sink__payload$24[35] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[36]$_SDFFE_PP0N_  (.CLK(clknet_leaf_300_clk_in_regs),
    .D(_04881_),
    .Q(\inst$top.soc.cpu.sink__payload$24[36] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[37]$_SDFFE_PP0N_  (.CLK(clknet_leaf_338_clk_in_regs),
    .D(_04882_),
    .Q(\inst$top.soc.cpu.d.sink__payload$16.rd_we ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[38]$_SDFFE_PP0N_  (.CLK(clknet_leaf_321_clk_in_regs),
    .D(_04883_),
    .Q(\inst$top.soc.cpu.sink__payload$24[38] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[39]$_SDFFE_PP0N_  (.CLK(clknet_leaf_320_clk_in_regs),
    .D(_04884_),
    .Q(\inst$top.soc.cpu.sink__payload$24[39] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_720_clk_in_regs),
    .D(_04885_),
    .Q(\inst$top.soc.cpu.sink__payload$24[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[40]$_SDFFE_PP0N_  (.CLK(clknet_leaf_320_clk_in_regs),
    .D(_04886_),
    .Q(\inst$top.soc.cpu.sink__payload$24[40] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[41]$_SDFFE_PP0N_  (.CLK(clknet_leaf_305_clk_in_regs),
    .D(_04887_),
    .Q(\inst$top.soc.cpu.sink__payload$24[41] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[42]$_SDFFE_PP0N_  (.CLK(clknet_leaf_315_clk_in_regs),
    .D(_04888_),
    .Q(\inst$top.soc.cpu.sink__payload$24[42] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[43]$_SDFFE_PP0N_  (.CLK(clknet_leaf_355_clk_in_regs),
    .D(_04889_),
    .Q(\inst$top.soc.cpu.sink__payload$24[43] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[44]$_SDFFE_PP0N_  (.CLK(clknet_leaf_346_clk_in_regs),
    .D(_04890_),
    .Q(\inst$top.soc.cpu.sink__payload$24[44] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[45]$_SDFFE_PP0N_  (.CLK(clknet_leaf_341_clk_in_regs),
    .D(_04891_),
    .Q(\inst$top.soc.cpu.sink__payload$24[45] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[46]$_SDFFE_PP0N_  (.CLK(clknet_leaf_351_clk_in_regs),
    .D(_04892_),
    .Q(\inst$top.soc.cpu.sink__payload$24[46] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[47]$_SDFFE_PP0N_  (.CLK(clknet_leaf_361_clk_in_regs),
    .D(_04893_),
    .Q(\inst$top.soc.cpu.sink__payload$24[47] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[48]$_SDFFE_PP0N_  (.CLK(clknet_leaf_357_clk_in_regs),
    .D(_04894_),
    .Q(\inst$top.soc.cpu.sink__payload$24[48] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[49]$_SDFFE_PP0N_  (.CLK(clknet_leaf_360_clk_in_regs),
    .D(_04895_),
    .Q(\inst$top.soc.cpu.sink__payload$24[49] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_732_clk_in_regs),
    .D(_04896_),
    .Q(\inst$top.soc.cpu.sink__payload$24[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[50]$_SDFFE_PP0N_  (.CLK(clknet_leaf_361_clk_in_regs),
    .D(_04897_),
    .Q(\inst$top.soc.cpu.sink__payload$24[50] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[51]$_SDFFE_PP0N_  (.CLK(clknet_leaf_355_clk_in_regs),
    .D(_04898_),
    .Q(\inst$top.soc.cpu.sink__payload$24[51] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[52]$_SDFFE_PP0N_  (.CLK(clknet_leaf_350_clk_in_regs),
    .D(_04899_),
    .Q(\inst$top.soc.cpu.sink__payload$24[52] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[53]$_SDFFE_PP0N_  (.CLK(clknet_leaf_369_clk_in_regs),
    .D(_04900_),
    .Q(\inst$top.soc.cpu.sink__payload$24[53] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[54]$_SDFFE_PP0N_  (.CLK(clknet_leaf_352_clk_in_regs),
    .D(_04901_),
    .Q(\inst$top.soc.cpu.sink__payload$24[54] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[55]$_SDFFE_PP0N_  (.CLK(clknet_leaf_358_clk_in_regs),
    .D(_04902_),
    .Q(\inst$top.soc.cpu.sink__payload$24[55] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[56]$_SDFFE_PP0N_  (.CLK(clknet_leaf_354_clk_in_regs),
    .D(_04903_),
    .Q(\inst$top.soc.cpu.sink__payload$24[56] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[57]$_SDFFE_PP0N_  (.CLK(clknet_leaf_379_clk_in_regs),
    .D(_04904_),
    .Q(\inst$top.soc.cpu.sink__payload$24[57] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[58]$_SDFFE_PP0N_  (.CLK(clknet_leaf_367_clk_in_regs),
    .D(_04905_),
    .Q(\inst$top.soc.cpu.sink__payload$24[58] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[59]$_SDFFE_PP0N_  (.CLK(clknet_leaf_303_clk_in_regs),
    .D(_04906_),
    .Q(\inst$top.soc.cpu.sink__payload$24[59] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_745_clk_in_regs),
    .D(_04907_),
    .Q(\inst$top.soc.cpu.sink__payload$24[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[60]$_SDFFE_PP0N_  (.CLK(clknet_leaf_352_clk_in_regs),
    .D(_04908_),
    .Q(\inst$top.soc.cpu.sink__payload$24[60] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[61]$_SDFFE_PP0N_  (.CLK(clknet_leaf_370_clk_in_regs),
    .D(_04909_),
    .Q(\inst$top.soc.cpu.sink__payload$24[61] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[62]$_SDFFE_PP0N_  (.CLK(clknet_leaf_369_clk_in_regs),
    .D(_04910_),
    .Q(\inst$top.soc.cpu.sink__payload$24[62] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[63]$_SDFFE_PP0N_  (.CLK(clknet_leaf_376_clk_in_regs),
    .D(_04911_),
    .Q(\inst$top.soc.cpu.sink__payload$24[63] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[64]$_SDFFE_PP0N_  (.CLK(clknet_leaf_379_clk_in_regs),
    .D(_04912_),
    .Q(\inst$top.soc.cpu.sink__payload$24[64] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[65]$_SDFFE_PP0N_  (.CLK(clknet_leaf_377_clk_in_regs),
    .D(_04913_),
    .Q(\inst$top.soc.cpu.sink__payload$24[65] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[66]$_SDFFE_PP0N_  (.CLK(clknet_leaf_349_clk_in_regs),
    .D(_04914_),
    .Q(\inst$top.soc.cpu.sink__payload$24[66] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[67]$_SDFFE_PP0N_  (.CLK(clknet_leaf_303_clk_in_regs),
    .D(_04915_),
    .Q(\inst$top.soc.cpu.sink__payload$24[67] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[68]$_SDFFE_PP0N_  (.CLK(clknet_leaf_357_clk_in_regs),
    .D(_04916_),
    .Q(\inst$top.soc.cpu.sink__payload$24[68] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[69]$_SDFFE_PP0N_  (.CLK(clknet_leaf_368_clk_in_regs),
    .D(_04917_),
    .Q(\inst$top.soc.cpu.sink__payload$24[69] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[6]$_SDFFE_PP0N_  (.CLK(clknet_leaf_741_clk_in_regs),
    .D(_04918_),
    .Q(\inst$top.soc.cpu.sink__payload$24[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[70]$_SDFFE_PP0N_  (.CLK(clknet_leaf_377_clk_in_regs),
    .D(_04919_),
    .Q(\inst$top.soc.cpu.sink__payload$24[70] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[71]$_SDFFE_PP0N_  (.CLK(clknet_leaf_358_clk_in_regs),
    .D(_04920_),
    .Q(\inst$top.soc.cpu.sink__payload$24[71] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[72]$_SDFFE_PP0N_  (.CLK(clknet_leaf_356_clk_in_regs),
    .D(_04921_),
    .Q(\inst$top.soc.cpu.sink__payload$24[72] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[73]$_SDFFE_PP0N_  (.CLK(clknet_leaf_303_clk_in_regs),
    .D(_04922_),
    .Q(\inst$top.soc.cpu.d.sink__payload$16.load ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[74]$_SDFFE_PP0N_  (.CLK(clknet_leaf_46_clk_in_regs),
    .D(_04923_),
    .Q(\inst$top.soc.cpu.sink__payload$24[74] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[75]$_SDFFE_PP0N_  (.CLK(clknet_leaf_312_clk_in_regs),
    .D(_04924_),
    .Q(\inst$top.soc.cpu.sink__payload$24[75] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[76]$_SDFFE_PP0N_  (.CLK(clknet_leaf_318_clk_in_regs),
    .D(_04925_),
    .Q(\inst$top.soc.cpu.sink__payload$24[76] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[77]$_SDFFE_PP0N_  (.CLK(clknet_leaf_317_clk_in_regs),
    .D(_04926_),
    .Q(\inst$top.soc.cpu.sink__payload$24[77] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[78]$_SDFFE_PP0N_  (.CLK(clknet_leaf_314_clk_in_regs),
    .D(_04927_),
    .Q(\inst$top.soc.cpu.sink__payload$24[78] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[79]$_SDFFE_PP0N_  (.CLK(clknet_leaf_309_clk_in_regs),
    .D(_04928_),
    .Q(\inst$top.soc.cpu.sink__payload$24[79] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[7]$_SDFFE_PP0N_  (.CLK(clknet_leaf_724_clk_in_regs),
    .D(_04929_),
    .Q(\inst$top.soc.cpu.sink__payload$24[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[80]$_SDFFE_PP0N_  (.CLK(clknet_leaf_308_clk_in_regs),
    .D(_04930_),
    .Q(\inst$top.soc.cpu.sink__payload$24[80] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[81]$_SDFFE_PP0N_  (.CLK(clknet_leaf_309_clk_in_regs),
    .D(_04931_),
    .Q(\inst$top.soc.cpu.sink__payload$24[81] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[82]$_SDFFE_PP0N_  (.CLK(clknet_leaf_315_clk_in_regs),
    .D(_04932_),
    .Q(\inst$top.soc.cpu.sink__payload$24[82] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[83]$_SDFFE_PP0N_  (.CLK(clknet_leaf_309_clk_in_regs),
    .D(_04933_),
    .Q(\inst$top.soc.cpu.sink__payload$24[83] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[84]$_SDFFE_PP0N_  (.CLK(clknet_leaf_316_clk_in_regs),
    .D(_04934_),
    .Q(\inst$top.soc.cpu.sink__payload$24[84] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[85]$_SDFFE_PP0N_  (.CLK(clknet_leaf_315_clk_in_regs),
    .D(_04935_),
    .Q(\inst$top.soc.cpu.sink__payload$24[85] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[86]$_SDFFE_PP0N_  (.CLK(clknet_leaf_315_clk_in_regs),
    .D(_04936_),
    .Q(\inst$top.soc.cpu.sink__payload$24[86] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[87]$_SDFFE_PP0N_  (.CLK(clknet_leaf_308_clk_in_regs),
    .D(_04937_),
    .Q(\inst$top.soc.cpu.sink__payload$24[87] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[88]$_SDFFE_PP0N_  (.CLK(clknet_leaf_308_clk_in_regs),
    .D(_04938_),
    .Q(\inst$top.soc.cpu.sink__payload$24[88] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[89]$_SDFFE_PP0N_  (.CLK(clknet_leaf_311_clk_in_regs),
    .D(_04939_),
    .Q(\inst$top.soc.cpu.sink__payload$24[89] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[8]$_SDFFE_PP0N_  (.CLK(clknet_leaf_743_clk_in_regs),
    .D(_04940_),
    .Q(\inst$top.soc.cpu.sink__payload$24[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[90]$_SDFFE_PP0N_  (.CLK(clknet_leaf_274_clk_in_regs),
    .D(_04941_),
    .Q(\inst$top.soc.cpu.sink__payload$24[90] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[91]$_SDFFE_PP0N_  (.CLK(clknet_leaf_275_clk_in_regs),
    .D(_04942_),
    .Q(\inst$top.soc.cpu.sink__payload$24[91] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[92]$_SDFFE_PP0N_  (.CLK(clknet_leaf_272_clk_in_regs),
    .D(_04943_),
    .Q(\inst$top.soc.cpu.sink__payload$24[92] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[93]$_SDFFE_PP0N_  (.CLK(clknet_leaf_276_clk_in_regs),
    .D(_04944_),
    .Q(\inst$top.soc.cpu.sink__payload$24[93] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[94]$_SDFFE_PP0N_  (.CLK(clknet_leaf_310_clk_in_regs),
    .D(_04945_),
    .Q(\inst$top.soc.cpu.sink__payload$24[94] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[95]$_SDFFE_PP0N_  (.CLK(clknet_leaf_273_clk_in_regs),
    .D(_04946_),
    .Q(\inst$top.soc.cpu.sink__payload$24[95] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[96]$_SDFFE_PP0N_  (.CLK(clknet_leaf_273_clk_in_regs),
    .D(_04947_),
    .Q(\inst$top.soc.cpu.sink__payload$24[96] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[97]$_SDFFE_PP0N_  (.CLK(clknet_leaf_310_clk_in_regs),
    .D(_04948_),
    .Q(\inst$top.soc.cpu.sink__payload$24[97] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[98]$_SDFFE_PP0N_  (.CLK(clknet_leaf_273_clk_in_regs),
    .D(_04949_),
    .Q(\inst$top.soc.cpu.sink__payload$24[98] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[99]$_SDFFE_PP0N_  (.CLK(clknet_leaf_309_clk_in_regs),
    .D(_04950_),
    .Q(\inst$top.soc.cpu.sink__payload$24[99] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$24[9]$_SDFFE_PP0N_  (.CLK(clknet_leaf_743_clk_in_regs),
    .D(_04951_),
    .Q(\inst$top.soc.cpu.sink__payload$24[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_756_clk_in_regs),
    .D(_04952_),
    .Q(\inst$top.soc.cpu.sink__payload$6[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_762_clk_in_regs),
    .D(_04953_),
    .Q(\inst$top.soc.cpu.sink__payload$6[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_760_clk_in_regs),
    .D(_04954_),
    .Q(\inst$top.soc.cpu.sink__payload$6[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_760_clk_in_regs),
    .D(_04955_),
    .Q(\inst$top.soc.cpu.sink__payload$6[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_759_clk_in_regs),
    .D(_04956_),
    .Q(\inst$top.soc.cpu.sink__payload$6[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_759_clk_in_regs),
    .D(_04957_),
    .Q(\inst$top.soc.cpu.sink__payload$6[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_768_clk_in_regs),
    .D(_04958_),
    .Q(\inst$top.soc.cpu.sink__payload$6[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_768_clk_in_regs),
    .D(_04959_),
    .Q(\inst$top.soc.cpu.sink__payload$6[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_765_clk_in_regs),
    .D(_04960_),
    .Q(\inst$top.soc.cpu.sink__payload$6[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_767_clk_in_regs),
    .D(_04961_),
    .Q(\inst$top.soc.cpu.sink__payload$6[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_765_clk_in_regs),
    .D(_04962_),
    .Q(\inst$top.soc.cpu.sink__payload$6[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_766_clk_in_regs),
    .D(_04963_),
    .Q(\inst$top.soc.cpu.sink__payload$6[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk_in_regs),
    .D(_04964_),
    .Q(\inst$top.soc.cpu.sink__payload$6[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk_in_regs),
    .D(_04965_),
    .Q(\inst$top.soc.cpu.sink__payload$6[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_19_clk_in_regs),
    .D(_04966_),
    .Q(\inst$top.soc.cpu.sink__payload$6[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk_in_regs),
    .D(_04967_),
    .Q(\inst$top.soc.cpu.sink__payload$6[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk_in_regs),
    .D(_04968_),
    .Q(\inst$top.soc.cpu.sink__payload$6[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk_in_regs),
    .D(_04969_),
    .Q(\inst$top.soc.cpu.sink__payload$6[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk_in_regs),
    .D(_04970_),
    .Q(\inst$top.soc.cpu.sink__payload$6[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk_in_regs),
    .D(_04971_),
    .Q(\inst$top.soc.cpu.sink__payload$6[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_778_clk_in_regs),
    .D(_04972_),
    .Q(\inst$top.soc.cpu.sink__payload$6[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_19_clk_in_regs),
    .D(_04973_),
    .Q(\inst$top.soc.cpu.sink__payload$6[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_776_clk_in_regs),
    .D(_04974_),
    .Q(\inst$top.soc.cpu.sink__payload$6[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[32]$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk_in_regs),
    .D(_04975_),
    .Q(\inst$top.soc.cpu.sink__payload$6[32] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[33]$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk_in_regs),
    .D(_04976_),
    .Q(\inst$top.soc.cpu.sink__payload$6[33] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[34]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk_in_regs),
    .D(_04977_),
    .Q(\inst$top.soc.cpu.sink__payload$6[34] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[35]$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk_in_regs),
    .D(_04978_),
    .Q(\inst$top.soc.cpu.sink__payload$6[35] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[36]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk_in_regs),
    .D(_04979_),
    .Q(\inst$top.soc.cpu.sink__payload$6[36] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[37]$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk_in_regs),
    .D(_04980_),
    .Q(\inst$top.soc.cpu.sink__payload$6[37] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[38]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk_in_regs),
    .D(_04981_),
    .Q(\inst$top.soc.cpu.sink__payload$6[38] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[39]$_SDFFE_PP0P_  (.CLK(clknet_leaf_315_clk_in_regs),
    .D(_04982_),
    .Q(\inst$top.soc.cpu.sink__payload$6[39] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_778_clk_in_regs),
    .D(_04983_),
    .Q(\inst$top.soc.cpu.sink__payload$6[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[40]$_SDFFE_PP0P_  (.CLK(clknet_leaf_316_clk_in_regs),
    .D(_04984_),
    .Q(\inst$top.soc.cpu.sink__payload$6[40] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[41]$_SDFFE_PP0P_  (.CLK(clknet_leaf_319_clk_in_regs),
    .D(_04985_),
    .Q(\inst$top.soc.cpu.sink__payload$6[41] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[42]$_SDFFE_PP0P_  (.CLK(clknet_leaf_318_clk_in_regs),
    .D(_04986_),
    .Q(\inst$top.soc.cpu.sink__payload$6[42] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[43]$_SDFFE_PP0P_  (.CLK(clknet_leaf_320_clk_in_regs),
    .D(_04987_),
    .Q(\inst$top.soc.cpu.sink__payload$6[43] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[44]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk_in_regs),
    .D(_04988_),
    .Q(\inst$top.soc.cpu.sink__payload$6[44] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[45]$_SDFFE_PP0P_  (.CLK(clknet_leaf_318_clk_in_regs),
    .D(_04989_),
    .Q(\inst$top.soc.cpu.sink__payload$6[45] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[46]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk_in_regs),
    .D(_04990_),
    .Q(\inst$top.soc.cpu.csr_fmt_i ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[47]$_SDFFE_PP0P_  (.CLK(clknet_leaf_311_clk_in_regs),
    .D(_04991_),
    .Q(\inst$top.soc.cpu.sink__payload$6[47] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[48]$_SDFFE_PP0P_  (.CLK(clknet_leaf_274_clk_in_regs),
    .D(_04992_),
    .Q(\inst$top.soc.cpu.sink__payload$6[48] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[49]$_SDFFE_PP0P_  (.CLK(clknet_leaf_274_clk_in_regs),
    .D(_04993_),
    .Q(\inst$top.soc.cpu.sink__payload$6[49] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_779_clk_in_regs),
    .D(_04994_),
    .Q(\inst$top.soc.cpu.sink__payload$6[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[50]$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk_in_regs),
    .D(_04995_),
    .Q(\inst$top.soc.cpu.sink__payload$6[50] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[51]$_SDFFE_PP0P_  (.CLK(clknet_leaf_312_clk_in_regs),
    .D(_04996_),
    .Q(\inst$top.soc.cpu.sink__payload$6[51] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[52]$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk_in_regs),
    .D(_04997_),
    .Q(\inst$top.soc.cpu.sink__payload$6[52] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[53]$_SDFFE_PP0P_  (.CLK(clknet_leaf_311_clk_in_regs),
    .D(_04998_),
    .Q(\inst$top.soc.cpu.sink__payload$6[53] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[54]$_SDFFE_PP0P_  (.CLK(clknet_leaf_273_clk_in_regs),
    .D(_04999_),
    .Q(\inst$top.soc.cpu.sink__payload$6[54] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[55]$_SDFFE_PP0P_  (.CLK(clknet_leaf_38_clk_in_regs),
    .D(_05000_),
    .Q(\inst$top.soc.cpu.sink__payload$6[55] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[56]$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk_in_regs),
    .D(_05001_),
    .Q(\inst$top.soc.cpu.sink__payload$6[56] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[57]$_SDFFE_PP0P_  (.CLK(clknet_leaf_31_clk_in_regs),
    .D(_05002_),
    .Q(\inst$top.soc.cpu.sink__payload$6[57] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[58]$_SDFFE_PP0P_  (.CLK(clknet_leaf_31_clk_in_regs),
    .D(_05003_),
    .Q(\inst$top.soc.cpu.sink__payload$6[58] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[59]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk_in_regs),
    .D(_05004_),
    .Q(\inst$top.soc.cpu.sink__payload$6[59] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_763_clk_in_regs),
    .D(_05005_),
    .Q(\inst$top.soc.cpu.sink__payload$6[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[60]$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk_in_regs),
    .D(_05006_),
    .Q(\inst$top.soc.cpu.sink__payload$6[60] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[61]$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk_in_regs),
    .D(_05007_),
    .Q(\inst$top.soc.cpu.sink__payload$6[61] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[62]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk_in_regs),
    .D(_05008_),
    .Q(\inst$top.soc.cpu.sink__payload$6[62] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[63]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk_in_regs),
    .D(_05009_),
    .Q(\inst$top.soc.cpu.sink__payload$6[63] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_763_clk_in_regs),
    .D(_05010_),
    .Q(\inst$top.soc.cpu.sink__payload$6[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_750_clk_in_regs),
    .D(_05011_),
    .Q(\inst$top.soc.cpu.sink__payload$6[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_752_clk_in_regs),
    .D(_05012_),
    .Q(\inst$top.soc.cpu.sink__payload$6[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload$6[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_752_clk_in_regs),
    .D(_05013_),
    .Q(\inst$top.soc.cpu.sink__payload$6[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[10]$_SDFFE_PP1P_  (.CLK(clknet_leaf_761_clk_in_regs),
    .D(_05014_),
    .Q(\inst$top.soc.cpu.sink__payload[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[11]$_SDFFE_PP1P_  (.CLK(clknet_leaf_764_clk_in_regs),
    .D(_05015_),
    .Q(\inst$top.soc.cpu.sink__payload[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[12]$_SDFFE_PP1P_  (.CLK(clknet_leaf_760_clk_in_regs),
    .D(_05016_),
    .Q(\inst$top.soc.cpu.sink__payload[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[13]$_SDFFE_PP1P_  (.CLK(clknet_leaf_759_clk_in_regs),
    .D(_05017_),
    .Q(\inst$top.soc.cpu.sink__payload[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[14]$_SDFFE_PP1P_  (.CLK(clknet_leaf_759_clk_in_regs),
    .D(_05018_),
    .Q(\inst$top.soc.cpu.sink__payload[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[15]$_SDFFE_PP1P_  (.CLK(clknet_leaf_22_clk_in_regs),
    .D(_05019_),
    .Q(\inst$top.soc.cpu.sink__payload[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[16]$_SDFFE_PP1P_  (.CLK(clknet_leaf_768_clk_in_regs),
    .D(_05020_),
    .Q(\inst$top.soc.cpu.sink__payload[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[17]$_SDFFE_PP1P_  (.CLK(clknet_leaf_768_clk_in_regs),
    .D(_05021_),
    .Q(\inst$top.soc.cpu.sink__payload[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[18]$_SDFFE_PP1P_  (.CLK(clknet_leaf_766_clk_in_regs),
    .D(_05022_),
    .Q(\inst$top.soc.cpu.sink__payload[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[19]$_SDFFE_PP1P_  (.CLK(clknet_leaf_767_clk_in_regs),
    .D(_05023_),
    .Q(\inst$top.soc.cpu.sink__payload[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_770_clk_in_regs),
    .D(_05024_),
    .Q(\inst$top.soc.cpu.sink__payload[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_769_clk_in_regs),
    .D(_05025_),
    .Q(\inst$top.soc.cpu.sink__payload[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_21_clk_in_regs),
    .D(_05026_),
    .Q(\inst$top.soc.cpu.sink__payload[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_21_clk_in_regs),
    .D(_05027_),
    .Q(\inst$top.soc.cpu.sink__payload[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_21_clk_in_regs),
    .D(_05028_),
    .Q(\inst$top.soc.cpu.sink__payload[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk_in_regs),
    .D(_05029_),
    .Q(\inst$top.soc.cpu.sink__payload[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk_in_regs),
    .D(_05030_),
    .Q(\inst$top.soc.cpu.sink__payload[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk_in_regs),
    .D(_05031_),
    .Q(\inst$top.soc.cpu.sink__payload[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk_in_regs),
    .D(_05032_),
    .Q(\inst$top.soc.cpu.sink__payload[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_19_clk_in_regs),
    .D(_05033_),
    .Q(\inst$top.soc.cpu.sink__payload[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[2]$_SDFFE_PP1P_  (.CLK(clknet_leaf_778_clk_in_regs),
    .D(_05034_),
    .Q(\inst$top.soc.cpu.sink__payload[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_19_clk_in_regs),
    .D(_05035_),
    .Q(\inst$top.soc.cpu.sink__payload[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_774_clk_in_regs),
    .D(_05036_),
    .Q(\inst$top.soc.cpu.sink__payload[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[3]$_SDFFE_PP1P_  (.CLK(clknet_leaf_777_clk_in_regs),
    .D(_05037_),
    .Q(\inst$top.soc.cpu.sink__payload[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[4]$_SDFFE_PP1P_  (.CLK(clknet_leaf_779_clk_in_regs),
    .D(_05038_),
    .Q(\inst$top.soc.cpu.sink__payload[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[5]$_SDFFE_PP1P_  (.CLK(clknet_leaf_764_clk_in_regs),
    .D(_05039_),
    .Q(\inst$top.soc.cpu.sink__payload[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[6]$_SDFFE_PP1P_  (.CLK(clknet_leaf_764_clk_in_regs),
    .D(_05040_),
    .Q(\inst$top.soc.cpu.sink__payload[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[7]$_SDFFE_PP1P_  (.CLK(clknet_leaf_764_clk_in_regs),
    .D(_05041_),
    .Q(\inst$top.soc.cpu.sink__payload[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[8]$_SDFFE_PP1P_  (.CLK(clknet_leaf_761_clk_in_regs),
    .D(_05042_),
    .Q(\inst$top.soc.cpu.sink__payload[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.sink__payload[9]$_SDFFE_PP1P_  (.CLK(clknet_leaf_761_clk_in_regs),
    .D(_05043_),
    .Q(\inst$top.soc.cpu.sink__payload[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.cpu.x.source__valid$_SDFFE_PP0N_  (.CLK(clknet_leaf_338_clk_in_regs),
    .D(_05044_),
    .Q(\inst$top.soc.cpu.x.source__valid ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__0._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_239_clk_in_regs),
    .D(_05045_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__0._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__0._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_239_clk_in_regs),
    .D(_05046_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__0._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__1._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_239_clk_in_regs),
    .D(_05047_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__1._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__1._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_239_clk_in_regs),
    .D(_05048_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__1._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__2._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_265_clk_in_regs),
    .D(_05049_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__2._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__2._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_265_clk_in_regs),
    .D(_05050_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__2._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__3._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_239_clk_in_regs),
    .D(_05051_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__3._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__3._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_239_clk_in_regs),
    .D(_05052_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__3._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__4._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_236_clk_in_regs),
    .D(_05053_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__4._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__4._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_237_clk_in_regs),
    .D(_05054_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__4._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__5._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_265_clk_in_regs),
    .D(_05055_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__5._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__5._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_263_clk_in_regs),
    .D(_05056_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__5._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__6._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_237_clk_in_regs),
    .D(_05057_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__6._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__6._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_237_clk_in_regs),
    .D(_05058_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__6._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__7._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_238_clk_in_regs),
    .D(_05059_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__7._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Mode.pin__7._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_238_clk_in_regs),
    .D(_05060_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Mode.pin__7._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Output.pin__0._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_238_clk_in_regs),
    .D(_05061_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__0._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Output.pin__1._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_239_clk_in_regs),
    .D(_05062_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__1._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Output.pin__2._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_265_clk_in_regs),
    .D(_05063_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__2._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Output.pin__3._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_240_clk_in_regs),
    .D(_05064_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__3._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Output.pin__4._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_237_clk_in_regs),
    .D(_05065_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__4._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Output.pin__5._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_264_clk_in_regs),
    .D(_05066_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__5._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Output.pin__6._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_237_clk_in_regs),
    .D(_05067_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__6._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.Output.pin__7._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_238_clk_in_regs),
    .D(_05068_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__7._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb$20$_SDFF_PP0_  (.CLK(clknet_leaf_271_clk_in_regs),
    .D(_05069_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb$20 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb$21$_SDFF_PP0_  (.CLK(clknet_leaf_270_clk_in_regs),
    .D(_05070_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb$21 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb$_SDFF_PP0_  (.CLK(clknet_leaf_271_clk_in_regs),
    .D(_05071_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_263_clk_in_regs),
    .D(_05072_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_263_clk_in_regs),
    .D(_05073_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_283_clk_in_regs),
    .D(_05074_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_264_clk_in_regs),
    .D(_05075_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_266_clk_in_regs),
    .D(_05076_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_282_clk_in_regs),
    .D(_05077_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_282_clk_in_regs),
    .D(_05078_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_263_clk_in_regs),
    .D(_05079_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_266_clk_in_regs),
    .D(_05080_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__0__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_265_clk_in_regs),
    .D(_05081_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_262_clk_in_regs),
    .D(_05082_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_265_clk_in_regs),
    .D(_05083_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_262_clk_in_regs),
    .D(_05084_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_266_clk_in_regs),
    .D(_05085_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_262_clk_in_regs),
    .D(_05086_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_267_clk_in_regs),
    .D(_05087_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_262_clk_in_regs),
    .D(_05088_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_270_clk_in_regs),
    .D(_05089_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.mux.r_shadow__1__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__0__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_240_clk_in_regs),
    .D(_05090_),
    .Q(\inst$top.soc.gpio_0._gpio.w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__0__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_241_clk_in_regs),
    .D(_05091_),
    .Q(\inst$top.soc.gpio_0._gpio.w_data$16 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__0__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_240_clk_in_regs),
    .D(_05092_),
    .Q(\inst$top.soc.gpio_0._gpio.w_data$26 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__0__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_241_clk_in_regs),
    .D(_05093_),
    .Q(\inst$top.soc.gpio_0._gpio.w_data$29 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__0__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_267_clk_in_regs),
    .D(_05094_),
    .Q(\inst$top.soc.gpio_0._gpio.w_data$38 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__0__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_267_clk_in_regs),
    .D(_05095_),
    .Q(\inst$top.soc.gpio_0._gpio.w_data$41 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__0__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_241_clk_in_regs),
    .D(_05096_),
    .Q(\inst$top.soc.gpio_0._gpio.w_data$50 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__0__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_241_clk_in_regs),
    .D(_05097_),
    .Q(\inst$top.soc.gpio_0._gpio.w_data$53 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__1__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_236_clk_in_regs),
    .D(_05098_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__0.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__1__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_241_clk_in_regs),
    .D(_05099_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__1.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__1__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_262_clk_in_regs),
    .D(_05100_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__2.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__1__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_261_clk_in_regs),
    .D(_05101_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__3.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__1__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_236_clk_in_regs),
    .D(_05102_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__4.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__1__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_261_clk_in_regs),
    .D(_05103_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__5.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__1__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_244_clk_in_regs),
    .D(_05104_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__6.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.bridge.mux.w_shadow__1__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_241_clk_in_regs),
    .D(_05105_),
    .Q(\inst$top.soc.gpio_0._gpio.bridge.Output.pin__7.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.pin_0_i_sync_ff_0$_DFF_P_  (.CLK(clknet_leaf_147_clk_in_regs),
    .D(net3017),
    .Q(\inst$top.soc.gpio_0._gpio.pin_0_i_sync_ff_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.pin_1_i_sync_ff_0$_DFF_P_  (.CLK(clknet_leaf_237_clk_in_regs),
    .D(net3016),
    .Q(\inst$top.soc.gpio_0._gpio.pin_1_i_sync_ff_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.pin_2_i_sync_ff_0$_DFF_P_  (.CLK(clknet_leaf_143_clk_in_regs),
    .D(net3029),
    .Q(\inst$top.soc.gpio_0._gpio.pin_2_i_sync_ff_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.pin_3_i_sync_ff_0$_DFF_P_  (.CLK(clknet_leaf_144_clk_in_regs),
    .D(net3028),
    .Q(\inst$top.soc.gpio_0._gpio.pin_3_i_sync_ff_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.pin_4_i_sync_ff_0$_DFF_P_  (.CLK(clknet_6_56__leaf_clk_in_regs),
    .D(net3027),
    .Q(\inst$top.soc.gpio_0._gpio.pin_4_i_sync_ff_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.pin_5_i_sync_ff_0$_DFF_P_  (.CLK(clknet_leaf_231_clk_in_regs),
    .D(net3026),
    .Q(\inst$top.soc.gpio_0._gpio.pin_5_i_sync_ff_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.pin_6_i_sync_ff_0$_DFF_P_  (.CLK(clknet_leaf_144_clk_in_regs),
    .D(net3025),
    .Q(\inst$top.soc.gpio_0._gpio.pin_6_i_sync_ff_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.pin_7_i_sync_ff_0$_DFF_P_  (.CLK(clknet_leaf_233_clk_in_regs),
    .D(net3024),
    .Q(\inst$top.soc.gpio_0._gpio.pin_7_i_sync_ff_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.r_data$23$_DFF_P_  (.CLK(clknet_leaf_225_clk_in_regs),
    .D(\inst$top.soc.gpio_0._gpio.pin_1_i_sync_ff_0 ),
    .Q(\inst$top.soc.gpio_0._gpio.r_data$23 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.r_data$35$_DFF_P_  (.CLK(clknet_leaf_147_clk_in_regs),
    .D(\inst$top.soc.gpio_0._gpio.pin_2_i_sync_ff_0 ),
    .Q(\inst$top.soc.gpio_0._gpio.r_data$35 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.r_data$47$_DFF_P_  (.CLK(clknet_leaf_144_clk_in_regs),
    .D(\inst$top.soc.gpio_0._gpio.pin_3_i_sync_ff_0 ),
    .Q(\inst$top.soc.gpio_0._gpio.r_data$47 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.r_data$59$_DFF_P_  (.CLK(clknet_leaf_189_clk_in_regs),
    .D(\inst$top.soc.gpio_0._gpio.pin_4_i_sync_ff_0 ),
    .Q(\inst$top.soc.gpio_0._gpio.r_data$59 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.r_data$71$_DFF_P_  (.CLK(clknet_6_50__leaf_clk_in_regs),
    .D(\inst$top.soc.gpio_0._gpio.pin_5_i_sync_ff_0 ),
    .Q(\inst$top.soc.gpio_0._gpio.r_data$71 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.r_data$83$_DFF_P_  (.CLK(clknet_leaf_144_clk_in_regs),
    .D(\inst$top.soc.gpio_0._gpio.pin_6_i_sync_ff_0 ),
    .Q(\inst$top.soc.gpio_0._gpio.r_data$83 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.r_data$95$_DFF_P_  (.CLK(clknet_6_56__leaf_clk_in_regs),
    .D(\inst$top.soc.gpio_0._gpio.pin_7_i_sync_ff_0 ),
    .Q(\inst$top.soc.gpio_0._gpio.r_data$95 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_0._gpio.r_data$_DFF_P_  (.CLK(clknet_leaf_143_clk_in_regs),
    .D(\inst$top.soc.gpio_0._gpio.pin_0_i_sync_ff_0 ),
    .Q(\inst$top.soc.gpio_0._gpio.r_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__0._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_246_clk_in_regs),
    .D(_05106_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__0._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__0._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_245_clk_in_regs),
    .D(_05107_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__0._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__1._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_245_clk_in_regs),
    .D(_05108_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__1._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__1._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_245_clk_in_regs),
    .D(_05109_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__1._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__2._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_236_clk_in_regs),
    .D(_05110_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__2._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__2._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_244_clk_in_regs),
    .D(_05111_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__2._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__3._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_245_clk_in_regs),
    .D(_05112_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__3._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__3._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_245_clk_in_regs),
    .D(_05113_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Mode.pin__3._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__0._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_246_clk_in_regs),
    .D(_05114_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__0._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__1._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_246_clk_in_regs),
    .D(_05115_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__1._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__2._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_244_clk_in_regs),
    .D(_05116_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__2._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__3._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_243_clk_in_regs),
    .D(_05117_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__3._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$14$_SDFF_PP0_  (.CLK(clknet_leaf_242_clk_in_regs),
    .D(_05118_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$14 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$15$_SDFF_PP0_  (.CLK(clknet_leaf_242_clk_in_regs),
    .D(_05119_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$15 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb$_SDFF_PP0_  (.CLK(clknet_leaf_238_clk_in_regs),
    .D(_05120_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_242_clk_in_regs),
    .D(_05121_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_243_clk_in_regs),
    .D(_05122_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_242_clk_in_regs),
    .D(_05123_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_247_clk_in_regs),
    .D(_05124_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_260_clk_in_regs),
    .D(_05125_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_260_clk_in_regs),
    .D(_05126_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_260_clk_in_regs),
    .D(_05127_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_261_clk_in_regs),
    .D(_05128_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_261_clk_in_regs),
    .D(_05129_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.r_shadow__0__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.w_shadow__0__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_249_clk_in_regs),
    .D(_05130_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__0.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.w_shadow__0__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_246_clk_in_regs),
    .D(_05131_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__1.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.w_shadow__0__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_247_clk_in_regs),
    .D(_05132_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__2.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.w_shadow__0__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_249_clk_in_regs),
    .D(_05133_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.bridge.Output.pin__3.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.w_shadow__0__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_243_clk_in_regs),
    .D(_05134_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.w_data$38 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.w_shadow__0__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_244_clk_in_regs),
    .D(_05135_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.w_data$41 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.w_shadow__0__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_247_clk_in_regs),
    .D(_05136_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.w_data$50 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.bridge.mux.w_shadow__0__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_243_clk_in_regs),
    .D(_05137_),
    .Q(\inst$top.soc.gpio_open_drain._gpio.w_data$53 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.pin_0_i_sync_ff_0$_DFF_P_  (.CLK(clknet_6_56__leaf_clk_in_regs),
    .D(net3023),
    .Q(\inst$top.soc.gpio_open_drain._gpio.pin_0_i_sync_ff_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.pin_1_i_sync_ff_0$_DFF_P_  (.CLK(clknet_leaf_140_clk_in_regs),
    .D(net3022),
    .Q(\inst$top.soc.gpio_open_drain._gpio.pin_1_i_sync_ff_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.pin_2_i_sync_ff_0$_DFF_P_  (.CLK(clknet_leaf_140_clk_in_regs),
    .D(net3021),
    .Q(\inst$top.soc.gpio_open_drain._gpio.pin_2_i_sync_ff_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.pin_3_i_sync_ff_0$_DFF_P_  (.CLK(clknet_leaf_135_clk_in_regs),
    .D(net3020),
    .Q(\inst$top.soc.gpio_open_drain._gpio.pin_3_i_sync_ff_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.r_data$23$_DFF_P_  (.CLK(clknet_6_50__leaf_clk_in_regs),
    .D(\inst$top.soc.gpio_open_drain._gpio.pin_1_i_sync_ff_0 ),
    .Q(\inst$top.soc.gpio_open_drain._gpio.r_data$23 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.r_data$35$_DFF_P_  (.CLK(clknet_leaf_246_clk_in_regs),
    .D(\inst$top.soc.gpio_open_drain._gpio.pin_2_i_sync_ff_0 ),
    .Q(\inst$top.soc.gpio_open_drain._gpio.r_data$35 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.r_data$47$_DFF_P_  (.CLK(clknet_6_50__leaf_clk_in_regs),
    .D(\inst$top.soc.gpio_open_drain._gpio.pin_3_i_sync_ff_0 ),
    .Q(\inst$top.soc.gpio_open_drain._gpio.r_data$47 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.gpio_open_drain._gpio.r_data$_DFF_P_  (.CLK(clknet_leaf_135_clk_in_regs),
    .D(\inst$top.soc.gpio_open_drain._gpio.pin_0_i_sync_ff_0 ),
    .Q(\inst$top.soc.gpio_open_drain._gpio.r_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_85_clk_in_regs),
    .D(_05138_),
    .Q(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.soc_id.bridge.mux.r_shadow__0__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_86_clk_in_regs),
    .D(_05139_),
    .Q(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.soc_id.bridge.mux.r_shadow__1__r_en$_SDFF_PP0_  (.CLK(clknet_6_33__leaf_clk_in_regs),
    .D(_05140_),
    .Q(\inst$top.soc.soc_id.bridge.mux.r_shadow__1__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.soc_id.bridge.mux.r_shadow__2__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_87_clk_in_regs),
    .D(_05141_),
    .Q(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.soc_id.bridge.mux.r_shadow__2__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_85_clk_in_regs),
    .D(_05142_),
    .Q(\inst$top.soc.soc_id.bridge.mux.r_shadow__0__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.soc_id.bridge.mux.r_shadow__2__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_85_clk_in_regs),
    .D(_05143_),
    .Q(\inst$top.soc.soc_id.bridge.mux.r_shadow__2__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.soc_id.bridge.mux.r_shadow__3__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_84_clk_in_regs),
    .D(_05144_),
    .Q(\inst$top.soc.soc_id.bridge.mux.r_shadow__3__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_55_clk_in_regs),
    .D(_05145_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk_in_regs),
    .D(_05146_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.dummy_bytes._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.Config.raw_enable._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk_in_regs),
    .D(_05147_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.raw_enable._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_54_clk_in_regs),
    .D(_05148_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_55_clk_in_regs),
    .D(_05149_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.width._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk_in_regs),
    .D(_05150_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_55_clk_in_regs),
    .D(_05151_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_56_clk_in_regs),
    .D(_05152_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_50_clk_in_regs),
    .D(_05153_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk_in_regs),
    .D(_05154_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_86_clk_in_regs),
    .D(_05155_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_51_clk_in_regs),
    .D(_05156_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_86_clk_in_regs),
    .D(_05157_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12._storage[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12.w_stb$_SDFF_PP0_  (.CLK(clknet_leaf_58_clk_in_regs),
    .D(_05158_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.RawTxData.data$12.w_stb ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb$16$_SDFF_PP0_  (.CLK(clknet_leaf_83_clk_in_regs),
    .D(_05159_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb$16 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb$17$_SDFF_PP0_  (.CLK(clknet_leaf_83_clk_in_regs),
    .D(_05160_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb$17 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb$_SDFF_PP0_  (.CLK(clknet_leaf_86_clk_in_regs),
    .D(_05161_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk_in_regs),
    .D(_05162_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_54_clk_in_regs),
    .D(_05163_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_54_clk_in_regs),
    .D(_05164_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_51_clk_in_regs),
    .D(_05165_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk_in_regs),
    .D(_05166_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_83_clk_in_regs),
    .D(_05167_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_82_clk_in_regs),
    .D(_05168_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_51_clk_in_regs),
    .D(_05169_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk_in_regs),
    .D(_05170_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.r_shadow__0__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk_in_regs),
    .D(_05171_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.Config.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_53_clk_in_regs),
    .D(_05172_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.RawControl.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_54_clk_in_regs),
    .D(_05173_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_53_clk_in_regs),
    .D(_05174_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_51_clk_in_regs),
    .D(_05175_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_85_clk_in_regs),
    .D(_05176_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_51_clk_in_regs),
    .D(_05177_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_86_clk_in_regs),
    .D(_05178_),
    .Q(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.w_shadow__0__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.fsm_state[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_58_clk_in_regs),
    .D(_05179_),
    .Q(\inst$top.soc.spiflash.ctrl.fsm_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.fsm_state[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_58_clk_in_regs),
    .D(_05180_),
    .Q(\inst$top.soc.spiflash.ctrl.fsm_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.fsm_state[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk_in_regs),
    .D(_05181_),
    .Q(\inst$top.soc.spiflash.ctrl.fsm_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.fsm_state[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk_in_regs),
    .D(_05182_),
    .Q(\inst$top.soc.spiflash.ctrl.fsm_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.i_data_count[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_785_clk_in_regs),
    .D(_05183_),
    .Q(\inst$top.soc.spiflash.ctrl.i_data_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.i_data_count[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_785_clk_in_regs),
    .D(_05184_),
    .Q(\inst$top.soc.spiflash.ctrl.i_data_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.i_data_count[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_785_clk_in_regs),
    .D(_05185_),
    .Q(\inst$top.soc.spiflash.ctrl.i_data_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.o_addr_count[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk_in_regs),
    .D(_05186_),
    .Q(\inst$top.soc.spiflash.ctrl.o_addr_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.o_addr_count[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk_in_regs),
    .D(_05187_),
    .Q(\inst$top.soc.spiflash.ctrl.o_addr_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.o_data_count[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_789_clk_in_regs),
    .D(_05188_),
    .Q(\inst$top.soc.spiflash.ctrl.o_data_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.o_data_count[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_789_clk_in_regs),
    .D(_05189_),
    .Q(\inst$top.soc.spiflash.ctrl.o_data_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.o_data_count[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_6_clk_in_regs),
    .D(_05190_),
    .Q(\inst$top.soc.spiflash.ctrl.o_data_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.o_dummy_count[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_16_clk_in_regs),
    .D(_05191_),
    .Q(\inst$top.soc.spiflash.ctrl.o_dummy_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.o_dummy_count[1]$_SDFFE_PP0P_  (.CLK(clknet_6_25__leaf_clk_in_regs),
    .D(_05192_),
    .Q(\inst$top.soc.spiflash.ctrl.o_dummy_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.r_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_52_clk_in_regs),
    .D(_05193_),
    .Q(\inst$top.soc.spiflash.ctrl.r_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.r_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_53_clk_in_regs),
    .D(_05194_),
    .Q(\inst$top.soc.spiflash.ctrl.r_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.r_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_60_clk_in_regs),
    .D(_05195_),
    .Q(\inst$top.soc.spiflash.ctrl.r_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.r_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_52_clk_in_regs),
    .D(_05196_),
    .Q(\inst$top.soc.spiflash.ctrl.r_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.r_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_52_clk_in_regs),
    .D(_05197_),
    .Q(\inst$top.soc.spiflash.ctrl.r_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.r_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_52_clk_in_regs),
    .D(_05198_),
    .Q(\inst$top.soc.spiflash.ctrl.r_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.r_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_81_clk_in_regs),
    .D(_05199_),
    .Q(\inst$top.soc.spiflash.ctrl.r_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.r_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_81_clk_in_regs),
    .D(_05200_),
    .Q(\inst$top.soc.spiflash.ctrl.r_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.raw_tx_data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_56_clk_in_regs),
    .D(_05201_),
    .Q(\inst$top.soc.spiflash.ctrl.raw_tx_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.raw_tx_data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk_in_regs),
    .D(_05202_),
    .Q(\inst$top.soc.spiflash.ctrl.raw_tx_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.raw_tx_data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_57_clk_in_regs),
    .D(_05203_),
    .Q(\inst$top.soc.spiflash.ctrl.raw_tx_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.raw_tx_data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_56_clk_in_regs),
    .D(_05204_),
    .Q(\inst$top.soc.spiflash.ctrl.raw_tx_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.raw_tx_data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_57_clk_in_regs),
    .D(_05205_),
    .Q(\inst$top.soc.spiflash.ctrl.raw_tx_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.raw_tx_data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_57_clk_in_regs),
    .D(_05206_),
    .Q(\inst$top.soc.spiflash.ctrl.raw_tx_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.raw_tx_data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_56_clk_in_regs),
    .D(_05207_),
    .Q(\inst$top.soc.spiflash.ctrl.raw_tx_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.raw_tx_data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_57_clk_in_regs),
    .D(_05208_),
    .Q(\inst$top.soc.spiflash.ctrl.raw_tx_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__ack$_SDFFE_PP0P_  (.CLK(clknet_leaf_58_clk_in_regs),
    .D(_05209_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__ack ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_787_clk_in_regs),
    .D(_05210_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_68_clk_in_regs),
    .D(_05211_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_68_clk_in_regs),
    .D(_05212_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_62_clk_in_regs),
    .D(_05213_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_61_clk_in_regs),
    .D(_05214_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_67_clk_in_regs),
    .D(_05215_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_66_clk_in_regs),
    .D(_05216_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_81_clk_in_regs),
    .D(_05217_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_69_clk_in_regs),
    .D(_05218_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_69_clk_in_regs),
    .D(_05219_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_71_clk_in_regs),
    .D(_05220_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk_in_regs),
    .D(_05221_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_70_clk_in_regs),
    .D(_05222_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_70_clk_in_regs),
    .D(_05223_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_71_clk_in_regs),
    .D(_05224_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_69_clk_in_regs),
    .D(_05225_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_58_clk_in_regs),
    .D(_05226_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_58_clk_in_regs),
    .D(_05227_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_64_clk_in_regs),
    .D(_05228_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_63_clk_in_regs),
    .D(_05229_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_58_clk_in_regs),
    .D(_05230_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_59_clk_in_regs),
    .D(_05231_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_66_clk_in_regs),
    .D(_05232_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_63_clk_in_regs),
    .D(_05233_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_63_clk_in_regs),
    .D(_05234_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_65_clk_in_regs),
    .D(_05235_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_64_clk_in_regs),
    .D(_05236_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_63_clk_in_regs),
    .D(_05237_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_65_clk_in_regs),
    .D(_05238_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_66_clk_in_regs),
    .D(_05239_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_60_clk_in_regs),
    .D(_05240_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.ctrl.wb_bus__dat_r[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_60_clk_in_regs),
    .D(_05241_),
    .Q(\inst$top.soc.spiflash.ctrl.wb_bus__dat_r[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.deframer.cycle[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_788_clk_in_regs),
    .D(_05242_),
    .Q(\inst$top.soc.spiflash.phy.deframer.cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.deframer.cycle[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_788_clk_in_regs),
    .D(_05243_),
    .Q(\inst$top.soc.spiflash.phy.deframer.cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.deframer.cycle[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_788_clk_in_regs),
    .D(_05244_),
    .Q(\inst$top.soc.spiflash.phy.deframer.cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.deframer.data_reg[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_787_clk_in_regs),
    .D(_05245_),
    .Q(\inst$top.soc.spiflash.phy.deframer.data_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.deframer.data_reg[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_787_clk_in_regs),
    .D(_05246_),
    .Q(\inst$top.soc.spiflash.phy.deframer.data_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.deframer.data_reg[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_787_clk_in_regs),
    .D(_05247_),
    .Q(\inst$top.soc.spiflash.phy.deframer.data_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.deframer.data_reg[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_786_clk_in_regs),
    .D(_05248_),
    .Q(\inst$top.soc.spiflash.phy.deframer.data_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.deframer.data_reg[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_786_clk_in_regs),
    .D(_05249_),
    .Q(\inst$top.soc.spiflash.phy.deframer.data_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.deframer.data_reg[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_786_clk_in_regs),
    .D(_05250_),
    .Q(\inst$top.soc.spiflash.phy.deframer.data_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.deframer.data_reg[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_786_clk_in_regs),
    .D(_05251_),
    .Q(\inst$top.soc.spiflash.phy.deframer.data_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.enframer.cycle[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_4_clk_in_regs),
    .D(_05252_),
    .Q(\inst$top.soc.spiflash.phy.enframer.cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.enframer.cycle[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_5_clk_in_regs),
    .D(_05253_),
    .Q(\inst$top.soc.spiflash.phy.enframer.cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.enframer.cycle[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_5_clk_in_regs),
    .D(_05254_),
    .Q(\inst$top.soc.spiflash.phy.enframer.cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.fsm_state$_SDFFE_PP0N_  (.CLK(clknet_leaf_6_clk_in_regs),
    .D(_05255_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.fsm_state ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[0]$_SDFFE_PP0P_  (.CLK(clknet_6_10__leaf_clk_in_regs),
    .D(_05256_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_784_clk_in_regs),
    .D(_05257_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_783_clk_in_regs),
    .D(_05258_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_783_clk_in_regs),
    .D(_05259_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_783_clk_in_regs),
    .D(_05260_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_784_clk_in_regs),
    .D(_05261_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_784_clk_in_regs),
    .D(_05262_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_781_clk_in_regs),
    .D(_05263_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_781_clk_in_regs),
    .D(_05264_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_9_clk_in_regs),
    .D(_05265_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_8_clk_in_regs),
    .D(_05266_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_9_clk_in_regs),
    .D(_05267_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_9_clk_in_regs),
    .D(_05268_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_781_clk_in_regs),
    .D(_05269_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_784_clk_in_regs),
    .D(_05270_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_clocker.timer[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_784_clk_in_regs),
    .D(_05271_),
    .Q(\inst$top.soc.spiflash.phy.io_clocker.timer[9] ));
 sky130_fd_sc_hd__dfxtp_4 \inst$top.soc.spiflash.phy.io_streamer.buffer_cs.o_ff$_DFF_P_  (.CLK(clknet_leaf_10_clk_in_regs),
    .D(\inst$top.soc.spiflash.phy.io_streamer.buffer_cs.o ),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.buffer_cs.o_ff ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.buffer_io0.i_ff$_DFF_P_  (.CLK(clknet_6_8__leaf_clk_in_regs),
    .D(net542),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.buffer_io0.i_ff ));
 sky130_fd_sc_hd__dfxtp_4 \inst$top.soc.spiflash.phy.io_streamer.buffer_io0.o_ff$_DFF_P_  (.CLK(clknet_leaf_749_clk_in_regs),
    .D(\inst$top.soc.spiflash.phy.io_streamer.buffer_io0.o ),
    .Q(net594));
 sky130_fd_sc_hd__dfxtp_4 \inst$top.soc.spiflash.phy.io_streamer.buffer_io0.oe_ff$_DFF_P_  (.CLK(clknet_leaf_773_clk_in_regs),
    .D(\inst$top.soc.spiflash.phy.io_streamer.buffer_io0.oe ),
    .Q(net560));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.buffer_io1.i_ff$_DFF_P_  (.CLK(clknet_leaf_789_clk_in_regs),
    .D(net543),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.buffer_io1.i_ff ));
 sky130_fd_sc_hd__dfxtp_4 \inst$top.soc.spiflash.phy.io_streamer.buffer_io1.o_ff$_DFF_P_  (.CLK(clknet_leaf_4_clk_in_regs),
    .D(\inst$top.soc.spiflash.phy.io_streamer.buffer_io1.o ),
    .Q(net595));
 sky130_fd_sc_hd__dfxtp_4 \inst$top.soc.spiflash.phy.io_streamer.buffer_io1.oe_ff$_DFF_P_  (.CLK(clknet_leaf_10_clk_in_regs),
    .D(\inst$top.soc.spiflash.phy.io_streamer.buffer_io1.oe ),
    .Q(net561));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.buffer_io2.i_ff$_DFF_P_  (.CLK(clknet_leaf_54_clk_in_regs),
    .D(net3019),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.buffer_io2.i_ff ));
 sky130_fd_sc_hd__dfxtp_4 \inst$top.soc.spiflash.phy.io_streamer.buffer_io2.o_ff$_DFF_P_  (.CLK(clknet_leaf_33_clk_in_regs),
    .D(\inst$top.soc.spiflash.phy.io_streamer.buffer_io2.o ),
    .Q(net596));
 sky130_fd_sc_hd__dfxtp_4 \inst$top.soc.spiflash.phy.io_streamer.buffer_io2.oe_ff$_DFF_P_  (.CLK(clknet_leaf_681_clk_in_regs),
    .D(\inst$top.soc.spiflash.phy.io_streamer.buffer_io2.oe ),
    .Q(net562));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.buffer_io3.i_ff$_DFF_P_  (.CLK(clknet_leaf_34_clk_in_regs),
    .D(net3018),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.buffer_io3.i_ff ));
 sky130_fd_sc_hd__dfxtp_4 \inst$top.soc.spiflash.phy.io_streamer.buffer_io3.o_ff$_DFF_P_  (.CLK(clknet_leaf_633_clk_in_regs),
    .D(\inst$top.soc.spiflash.phy.io_streamer.buffer_io3.o ),
    .Q(net597));
 sky130_fd_sc_hd__dfxtp_4 \inst$top.soc.spiflash.phy.io_streamer.buffer_io3.oe_ff$_DFF_P_  (.CLK(clknet_leaf_675_clk_in_regs),
    .D(\inst$top.soc.spiflash.phy.io_streamer.buffer_io3.oe ),
    .Q(net563));
 sky130_fd_sc_hd__dfxtp_4 \inst$top.soc.spiflash.phy.io_streamer.buffer_sck.o_ff$_DFF_P_  (.CLK(clknet_6_0__leaf_clk_in_regs),
    .D(\inst$top.soc.spiflash.phy.io_streamer.buffer_sck.o ),
    .Q(net582));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.i_en_0$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk_in_regs),
    .D(_05272_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.i_en_0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.meta_0[0]$_SDFF_PP0_  (.CLK(clknet_leaf_790_clk_in_regs),
    .D(_05273_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.meta_0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.meta_0[1]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk_in_regs),
    .D(_05274_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.meta_0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.meta_0[2]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk_in_regs),
    .D(_05275_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.meta_0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.o_latch[0]$_SDFF_PP1_  (.CLK(clknet_leaf_8_clk_in_regs),
    .D(_05276_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.o_latch.sck.o ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.o_latch[10]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk_in_regs),
    .D(_05277_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.o_latch.cs.o ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.o_latch[2]$_SDFF_PP0_  (.CLK(clknet_leaf_756_clk_in_regs),
    .D(_05278_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io0.o ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.o_latch[3]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk_in_regs),
    .D(_05279_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io0.oe ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.o_latch[4]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk_in_regs),
    .D(_05280_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io1.o ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.o_latch[5]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk_in_regs),
    .D(_05281_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io1.oe ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.o_latch[6]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk_in_regs),
    .D(_05282_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io2.o ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.o_latch[7]$_SDFF_PP0_  (.CLK(clknet_leaf_678_clk_in_regs),
    .D(_05283_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io2.oe ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.o_latch[8]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk_in_regs),
    .D(_05284_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io3.o ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.o_latch[9]$_SDFF_PP0_  (.CLK(clknet_leaf_679_clk_in_regs),
    .D(_05285_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.o_latch.io3.oe ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.skid_1[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk_in_regs),
    .D(_05286_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io0 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.skid_1[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_789_clk_in_regs),
    .D(_05287_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io1 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.skid_1[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk_in_regs),
    .D(_05288_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io2 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.skid_1[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk_in_regs),
    .D(_05289_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.skid_1.port.io3 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.skid_1[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_789_clk_in_regs),
    .D(_05290_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.skid_1.meta[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.skid_1[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk_in_regs),
    .D(_05291_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.skid_1.meta[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.skid_1[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk_in_regs),
    .D(_05292_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.skid_1.meta[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.spiflash.phy.io_streamer.skid_at$_SDFFE_PP0P_  (.CLK(clknet_leaf_790_clk_in_regs),
    .D(_05293_),
    .Q(\inst$top.soc.spiflash.phy.io_streamer.skid_at ));
 CF_SRAM_1024x32 \inst$top.soc.sram.mem.0.0  (.WLBI(net433),
    .CLKin(clknet_1_0__leaf_clk_in),
    .EN(net529),
    .R_WB(_00161_),
    .SM(net434),
    .TM(net435),
    .ScanInDR(net436),
    .ScanInDL(net437),
    .ScanInCC(net440),
    .vpwrpc(net530),
    .vpwrac(net531),
    .AD({net439,
    net438,
    net1833,
    \inst$top.soc.bus__adr[6] ,
    net1834,
    \inst$top.soc.bus__adr[4] ,
    \inst$top.soc.bus__adr[3] ,
    \inst$top.soc.bus__adr[2] ,
    \inst$top.soc.bus__addr[3] ,
    \inst$top.soc.bus__addr[2] }),
    .BEN({net758,
    net758,
    net758,
    net758,
    net758,
    net758,
    net758,
    net758,
    net756,
    net756,
    net756,
    net756,
    net756,
    net756,
    net756,
    net756,
    net762,
    net761,
    net761,
    net761,
    net761,
    net761,
    net761,
    net761,
    net760,
    net760,
    net760,
    net760,
    net760,
    net760,
    net760,
    net760}),
    .DI({\inst$top.soc.bus__dat_w[31] ,
    \inst$top.soc.bus__dat_w[30] ,
    \inst$top.soc.bus__dat_w[29] ,
    \inst$top.soc.bus__dat_w[28] ,
    \inst$top.soc.bus__dat_w[27] ,
    \inst$top.soc.bus__dat_w[26] ,
    \inst$top.soc.bus__dat_w[25] ,
    \inst$top.soc.bus__dat_w[24] ,
    \inst$top.soc.bus__dat_w[23] ,
    \inst$top.soc.bus__dat_w[22] ,
    \inst$top.soc.bus__dat_w[21] ,
    \inst$top.soc.bus__dat_w[20] ,
    \inst$top.soc.bus__dat_w[19] ,
    \inst$top.soc.bus__dat_w[18] ,
    \inst$top.soc.bus__dat_w[17] ,
    \inst$top.soc.bus__dat_w[16] ,
    \inst$top.soc.bus__dat_w[15] ,
    \inst$top.soc.bus__dat_w[14] ,
    \inst$top.soc.bus__dat_w[13] ,
    \inst$top.soc.bus__dat_w[12] ,
    \inst$top.soc.bus__dat_w[11] ,
    \inst$top.soc.bus__dat_w[10] ,
    \inst$top.soc.bus__dat_w[9] ,
    \inst$top.soc.bus__dat_w[8] ,
    \inst$top.soc.bus__dat_w[7] ,
    \inst$top.soc.bus__dat_w[6] ,
    \inst$top.soc.bus__dat_w[5] ,
    \inst$top.soc.bus__dat_w[4] ,
    \inst$top.soc.bus__dat_w[3] ,
    \inst$top.soc.bus__dat_w[2] ,
    \inst$top.soc.bus__dat_w[1] ,
    \inst$top.soc.bus__dat_w[0] }),
    .DO({_00088_,
    _00087_,
    _00085_,
    _00084_,
    _00083_,
    _00082_,
    _00081_,
    _00080_,
    _00079_,
    _00078_,
    _00077_,
    _00076_,
    _00074_,
    _00073_,
    _00072_,
    _00071_,
    _00070_,
    _00069_,
    _00068_,
    _00067_,
    _00066_,
    _00065_,
    _00095_,
    _00094_,
    _00093_,
    _00092_,
    _00091_,
    _00090_,
    _00089_,
    _00086_,
    _00075_,
    _00064_}));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.sram.wb_bus__ack$_SDFF_PP0_  (.CLK(clknet_leaf_56_clk_in_regs),
    .D(_05294_),
    .Q(\inst$top.soc.sram.wb_bus__ack ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.bitno[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_134_clk_in_regs),
    .D(_05295_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.bitno[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.bitno[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_134_clk_in_regs),
    .D(_05296_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.bitno[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.bitno[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_138_clk_in_regs),
    .D(_05297_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.bitno[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.bitno[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_134_clk_in_regs),
    .D(_05298_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.bitno[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_260_clk_in_regs),
    .D(_05299_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_259_clk_in_regs),
    .D(_05300_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_254_clk_in_regs),
    .D(_05301_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_252_clk_in_regs),
    .D(_05302_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_252_clk_in_regs),
    .D(_05303_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_252_clk_in_regs),
    .D(_05304_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_254_clk_in_regs),
    .D(_05305_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_259_clk_in_regs),
    .D(_05306_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.err[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_260_clk_in_regs),
    .D(_05307_),
    .Q(\inst$top.soc.uart_0._phy.rx.err.frame ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.fsm_state[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_250_clk_in_regs),
    .D(_05308_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.fsm_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.fsm_state[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_250_clk_in_regs),
    .D(_05309_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.fsm_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.rdy$_SDFF_PP0_  (.CLK(clknet_leaf_258_clk_in_regs),
    .D(_05310_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.rdy ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.shreg[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_248_clk_in_regs),
    .D(_05311_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.shreg.start ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.shreg[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_248_clk_in_regs),
    .D(_05312_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.shreg[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.shreg[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_254_clk_in_regs),
    .D(_05313_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.shreg[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.shreg[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_253_clk_in_regs),
    .D(_05314_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.shreg[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.shreg[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_252_clk_in_regs),
    .D(_05315_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.shreg[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.shreg[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_253_clk_in_regs),
    .D(_05316_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.shreg[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.shreg[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_253_clk_in_regs),
    .D(_05317_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.shreg[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.shreg[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_254_clk_in_regs),
    .D(_05318_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.shreg[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.shreg[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_254_clk_in_regs),
    .D(_05319_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.shreg[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.shreg[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_248_clk_in_regs),
    .D(_05320_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.shreg.stop ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_104_clk_in_regs),
    .D(_05321_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_110_clk_in_regs),
    .D(_05322_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_110_clk_in_regs),
    .D(_05323_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_252_clk_in_regs),
    .D(_05324_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_255_clk_in_regs),
    .D(_05325_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_252_clk_in_regs),
    .D(_05326_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_255_clk_in_regs),
    .D(_05327_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_111_clk_in_regs),
    .D(_05328_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_109_clk_in_regs),
    .D(_05329_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_108_clk_in_regs),
    .D(_05330_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_108_clk_in_regs),
    .D(_05331_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_103_clk_in_regs),
    .D(_05332_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_108_clk_in_regs),
    .D(_05333_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_107_clk_in_regs),
    .D(_05334_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_109_clk_in_regs),
    .D(_05335_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_109_clk_in_regs),
    .D(_05336_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_103_clk_in_regs),
    .D(_05337_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[3]$_SDFFE_PP1P_  (.CLK(clknet_leaf_114_clk_in_regs),
    .D(_05338_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[4]$_SDFFE_PP1P_  (.CLK(clknet_leaf_114_clk_in_regs),
    .D(_05339_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_103_clk_in_regs),
    .D(_05340_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[6]$_SDFFE_PP1P_  (.CLK(clknet_leaf_114_clk_in_regs),
    .D(_05341_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[7]$_SDFFE_PP1P_  (.CLK(clknet_6_34__leaf_clk_in_regs),
    .D(_05342_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[8]$_SDFFE_PP0P_  (.CLK(clknet_6_42__leaf_clk_in_regs),
    .D(_05343_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.lower.timer[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_111_clk_in_regs),
    .D(_05344_),
    .Q(\inst$top.soc.uart_0._phy.rx.lower.timer[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.overflow$_SDFF_PP0_  (.CLK(clknet_leaf_267_clk_in_regs),
    .D(_05345_),
    .Q(\inst$top.soc.uart_0._phy.rx.overflow ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.symbols__payload[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_258_clk_in_regs),
    .D(_05346_),
    .Q(\inst$top.soc.uart_0._phy.rx.symbols__payload[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.symbols__payload[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_259_clk_in_regs),
    .D(_05347_),
    .Q(\inst$top.soc.uart_0._phy.rx.symbols__payload[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.symbols__payload[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_254_clk_in_regs),
    .D(_05348_),
    .Q(\inst$top.soc.uart_0._phy.rx.symbols__payload[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.symbols__payload[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_256_clk_in_regs),
    .D(_05349_),
    .Q(\inst$top.soc.uart_0._phy.rx.symbols__payload[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.symbols__payload[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_255_clk_in_regs),
    .D(_05350_),
    .Q(\inst$top.soc.uart_0._phy.rx.symbols__payload[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.symbols__payload[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_255_clk_in_regs),
    .D(_05351_),
    .Q(\inst$top.soc.uart_0._phy.rx.symbols__payload[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.symbols__payload[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_259_clk_in_regs),
    .D(_05352_),
    .Q(\inst$top.soc.uart_0._phy.rx.symbols__payload[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.symbols__payload[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_259_clk_in_regs),
    .D(_05353_),
    .Q(\inst$top.soc.uart_0._phy.rx.symbols__payload[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.rx.symbols__valid$_SDFFE_PP0P_  (.CLK(clknet_leaf_267_clk_in_regs),
    .D(_05354_),
    .Q(\inst$top.soc.uart_0._phy.rx.symbols__valid ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.bitno[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_115_clk_in_regs),
    .D(_05355_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.bitno[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.bitno[1]$_SDFFE_PP0P_  (.CLK(clknet_6_34__leaf_clk_in_regs),
    .D(_05356_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.bitno[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.bitno[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_113_clk_in_regs),
    .D(_05357_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.bitno[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.bitno[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_118_clk_in_regs),
    .D(_05358_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.bitno[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.fsm_state$_SDFF_PP0_  (.CLK(clknet_leaf_116_clk_in_regs),
    .D(_05359_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.fsm_state ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.o$_SDFFE_PP1P_  (.CLK(clknet_leaf_115_clk_in_regs),
    .D(_05360_),
    .Q(net598));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.shreg[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_113_clk_in_regs),
    .D(_05361_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.shreg.start ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.shreg[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_115_clk_in_regs),
    .D(_05362_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.shreg[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.shreg[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_102_clk_in_regs),
    .D(_05363_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.shreg[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.shreg[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_116_clk_in_regs),
    .D(_05364_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.shreg[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.shreg[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_100_clk_in_regs),
    .D(_05365_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.shreg[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.shreg[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_117_clk_in_regs),
    .D(_05366_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.shreg[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.shreg[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_117_clk_in_regs),
    .D(_05367_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.shreg[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.shreg[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_117_clk_in_regs),
    .D(_05368_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.shreg[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.shreg[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_117_clk_in_regs),
    .D(_05369_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.shreg[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.shreg[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_116_clk_in_regs),
    .D(_05370_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.shreg.stop ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_118_clk_in_regs),
    .D(_05371_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_123_clk_in_regs),
    .D(_05372_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_121_clk_in_regs),
    .D(_05373_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_123_clk_in_regs),
    .D(_05374_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_121_clk_in_regs),
    .D(_05375_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_121_clk_in_regs),
    .D(_05376_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_121_clk_in_regs),
    .D(_05377_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[16]$_SDFFE_PP0P_  (.CLK(clknet_6_33__leaf_clk_in_regs),
    .D(_05378_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_124_clk_in_regs),
    .D(_05379_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_124_clk_in_regs),
    .D(_05380_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_75_clk_in_regs),
    .D(_05381_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_119_clk_in_regs),
    .D(_05382_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk_in_regs),
    .D(_05383_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk_in_regs),
    .D(_05384_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_124_clk_in_regs),
    .D(_05385_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_123_clk_in_regs),
    .D(_05386_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_118_clk_in_regs),
    .D(_05387_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[3]$_SDFFE_PP1P_  (.CLK(clknet_leaf_117_clk_in_regs),
    .D(_05388_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[4]$_SDFFE_PP1P_  (.CLK(clknet_leaf_123_clk_in_regs),
    .D(_05389_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_99_clk_in_regs),
    .D(_05390_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[6]$_SDFFE_PP1P_  (.CLK(clknet_leaf_119_clk_in_regs),
    .D(_05391_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[7]$_SDFFE_PP1P_  (.CLK(clknet_leaf_119_clk_in_regs),
    .D(_05392_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_121_clk_in_regs),
    .D(_05393_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._phy.tx.lower.timer[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_121_clk_in_regs),
    .D(_05394_),
    .Q(\inst$top.soc.uart_0._phy.tx.lower.timer[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.Config.enable._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_269_clk_in_regs),
    .D(_05395_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.Config.enable._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_268_clk_in_regs),
    .D(_05396_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_249_clk_in_regs),
    .D(_05397_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_110_clk_in_regs),
    .D(_05398_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_110_clk_in_regs),
    .D(_05399_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_249_clk_in_regs),
    .D(_05400_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_255_clk_in_regs),
    .D(_05401_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_138_clk_in_regs),
    .D(_05402_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_258_clk_in_regs),
    .D(_05403_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_115_clk_in_regs),
    .D(_05404_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_104_clk_in_regs),
    .D(_05405_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_256_clk_in_regs),
    .D(_05406_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_93_clk_in_regs),
    .D(_05407_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_107_clk_in_regs),
    .D(_05408_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_104_clk_in_regs),
    .D(_05409_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_104_clk_in_regs),
    .D(_05410_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_103_clk_in_regs),
    .D(_05411_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_93_clk_in_regs),
    .D(_05412_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[3]$_SDFFE_PP1P_  (.CLK(clknet_leaf_107_clk_in_regs),
    .D(_05413_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[4]$_SDFFE_PP1P_  (.CLK(clknet_leaf_268_clk_in_regs),
    .D(_05414_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_106_clk_in_regs),
    .D(_05415_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[6]$_SDFFE_PP1P_  (.CLK(clknet_leaf_106_clk_in_regs),
    .D(_05416_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[7]$_SDFFE_PP1P_  (.CLK(clknet_leaf_257_clk_in_regs),
    .D(_05417_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_110_clk_in_regs),
    .D(_05418_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_110_clk_in_regs),
    .D(_05419_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.PhyConfig.U$0._storage[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.Status.error._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_268_clk_in_regs),
    .D(_05420_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.Status.error._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.Status.overflow._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_270_clk_in_regs),
    .D(_05421_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.Status.overflow._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb$25$_SDFF_PP0_  (.CLK(clknet_leaf_268_clk_in_regs),
    .D(_05422_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb$25 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb$34$_SDFF_PP0_  (.CLK(clknet_leaf_92_clk_in_regs),
    .D(_05423_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb$34 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb$_SDFF_PP0_  (.CLK(clknet_leaf_269_clk_in_regs),
    .D(_05424_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.element__w_stb ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_92_clk_in_regs),
    .D(_05425_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_92_clk_in_regs),
    .D(_05426_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_91_clk_in_regs),
    .D(_05427_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_268_clk_in_regs),
    .D(_05428_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_267_clk_in_regs),
    .D(_05429_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_93_clk_in_regs),
    .D(_05430_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_93_clk_in_regs),
    .D(_05431_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_268_clk_in_regs),
    .D(_05432_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_269_clk_in_regs),
    .D(_05433_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__0__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_258_clk_in_regs),
    .D(_05434_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_268_clk_in_regs),
    .D(_05435_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_93_clk_in_regs),
    .D(_05436_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_256_clk_in_regs),
    .D(_05437_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_256_clk_in_regs),
    .D(_05438_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_93_clk_in_regs),
    .D(_05439_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_267_clk_in_regs),
    .D(_05440_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_257_clk_in_regs),
    .D(_05441_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_91_clk_in_regs),
    .D(_05442_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__1__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_257_clk_in_regs),
    .D(_05443_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_93_clk_in_regs),
    .D(_05444_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_94_clk_in_regs),
    .D(_05445_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_256_clk_in_regs),
    .D(_05446_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_256_clk_in_regs),
    .D(_05447_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_105_clk_in_regs),
    .D(_05448_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_94_clk_in_regs),
    .D(_05449_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_107_clk_in_regs),
    .D(_05450_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_91_clk_in_regs),
    .D(_05451_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.r_shadow__2__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_269_clk_in_regs),
    .D(_05452_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.Config.enable.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_270_clk_in_regs),
    .D(_05453_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.Status.overflow.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_268_clk_in_regs),
    .D(_05454_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.Status.error.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_106_clk_in_regs),
    .D(_05455_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_268_clk_in_regs),
    .D(_05456_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_106_clk_in_regs),
    .D(_05457_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_106_clk_in_regs),
    .D(_05458_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_107_clk_in_regs),
    .D(_05459_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__0__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_251_clk_in_regs),
    .D(_05460_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_110_clk_in_regs),
    .D(_05461_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_250_clk_in_regs),
    .D(_05462_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_138_clk_in_regs),
    .D(_05463_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_251_clk_in_regs),
    .D(_05464_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[5]$_SDFFE_PP0P_  (.CLK(clknet_6_50__leaf_clk_in_regs),
    .D(_05465_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_255_clk_in_regs),
    .D(_05466_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_138_clk_in_regs),
    .D(_05467_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__1__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_256_clk_in_regs),
    .D(_05468_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_115_clk_in_regs),
    .D(_05469_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_102_clk_in_regs),
    .D(_05470_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_255_clk_in_regs),
    .D(_05471_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_107_clk_in_regs),
    .D(_05472_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_104_clk_in_regs),
    .D(_05473_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_102_clk_in_regs),
    .D(_05474_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_102_clk_in_regs),
    .D(_05475_),
    .Q(\inst$top.soc.uart_0._uart.rx.bridge.mux.w_shadow__2__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.Config.enable._storage$_SDFFE_PP0P_  (.CLK(clknet_leaf_90_clk_in_regs),
    .D(_05476_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.Config.enable._storage ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_96_clk_in_regs),
    .D(_05477_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_76_clk_in_regs),
    .D(_05478_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_75_clk_in_regs),
    .D(_05479_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_75_clk_in_regs),
    .D(_05480_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_76_clk_in_regs),
    .D(_05481_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_75_clk_in_regs),
    .D(_05482_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_75_clk_in_regs),
    .D(_05483_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_76_clk_in_regs),
    .D(_05484_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_78_clk_in_regs),
    .D(_05485_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_79_clk_in_regs),
    .D(_05486_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_74_clk_in_regs),
    .D(_05487_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_98_clk_in_regs),
    .D(_05488_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_74_clk_in_regs),
    .D(_05489_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_80_clk_in_regs),
    .D(_05490_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_79_clk_in_regs),
    .D(_05491_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_80_clk_in_regs),
    .D(_05492_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_97_clk_in_regs),
    .D(_05493_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[3]$_SDFFE_PP1P_  (.CLK(clknet_leaf_96_clk_in_regs),
    .D(_05494_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[4]$_SDFFE_PP1P_  (.CLK(clknet_leaf_94_clk_in_regs),
    .D(_05495_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_100_clk_in_regs),
    .D(_05496_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[6]$_SDFFE_PP1P_  (.CLK(clknet_6_34__leaf_clk_in_regs),
    .D(_05497_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[7]$_SDFFE_PP1P_  (.CLK(clknet_leaf_94_clk_in_regs),
    .D(_05498_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_99_clk_in_regs),
    .D(_05499_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_76_clk_in_regs),
    .D(_05500_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.PhyConfig.U$0._storage[9] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb$27$_SDFF_PP0_  (.CLK(clknet_leaf_91_clk_in_regs),
    .D(_05501_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb$27 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb$32$_SDFF_PP0_  (.CLK(clknet_leaf_90_clk_in_regs),
    .D(_05502_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb$32 ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb$_SDFF_PP0_  (.CLK(clknet_leaf_89_clk_in_regs),
    .D(_05503_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.element__w_stb ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_90_clk_in_regs),
    .D(_05504_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_90_clk_in_regs),
    .D(_05505_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_95_clk_in_regs),
    .D(_05506_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_96_clk_in_regs),
    .D(_05507_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_96_clk_in_regs),
    .D(_05508_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_95_clk_in_regs),
    .D(_05509_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_96_clk_in_regs),
    .D(_05510_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_96_clk_in_regs),
    .D(_05511_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_95_clk_in_regs),
    .D(_05512_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__0__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_97_clk_in_regs),
    .D(_05513_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_77_clk_in_regs),
    .D(_05514_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_77_clk_in_regs),
    .D(_05515_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_77_clk_in_regs),
    .D(_05516_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_77_clk_in_regs),
    .D(_05517_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_77_clk_in_regs),
    .D(_05518_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_78_clk_in_regs),
    .D(_05519_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_78_clk_in_regs),
    .D(_05520_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_87_clk_in_regs),
    .D(_05521_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__1__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_79_clk_in_regs),
    .D(_05522_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_84_clk_in_regs),
    .D(_05523_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_79_clk_in_regs),
    .D(_05524_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_79_clk_in_regs),
    .D(_05525_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_84_clk_in_regs),
    .D(_05526_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_78_clk_in_regs),
    .D(_05527_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_77_clk_in_regs),
    .D(_05528_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_78_clk_in_regs),
    .D(_05529_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__r_en$_SDFF_PP0_  (.CLK(clknet_leaf_89_clk_in_regs),
    .D(_05530_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.r_shadow__2__r_en ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_95_clk_in_regs),
    .D(_05531_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.Config.enable.port__w_data ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_100_clk_in_regs),
    .D(_05532_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_98_clk_in_regs),
    .D(_05533_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_97_clk_in_regs),
    .D(_05534_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_94_clk_in_regs),
    .D(_05535_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_105_clk_in_regs),
    .D(_05536_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_94_clk_in_regs),
    .D(_05537_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_95_clk_in_regs),
    .D(_05538_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__0__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_102_clk_in_regs),
    .D(_05539_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_102_clk_in_regs),
    .D(_05540_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_100_clk_in_regs),
    .D(_05541_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_100_clk_in_regs),
    .D(_05542_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_100_clk_in_regs),
    .D(_05543_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_99_clk_in_regs),
    .D(_05544_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_99_clk_in_regs),
    .D(_05545_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_99_clk_in_regs),
    .D(_05546_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__1__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_76_clk_in_regs),
    .D(_05547_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_78_clk_in_regs),
    .D(_05548_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_74_clk_in_regs),
    .D(_05549_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_71_clk_in_regs),
    .D(_05550_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk_in_regs),
    .D(_05551_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_80_clk_in_regs),
    .D(_05552_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_71_clk_in_regs),
    .D(_05553_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_82_clk_in_regs),
    .D(_05554_),
    .Q(\inst$top.soc.uart_0._uart.tx.bridge.mux.w_shadow__2__data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_arbiter.grant$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk_in_regs),
    .D(_05555_),
    .Q(\inst$top.soc.wb_arbiter.grant ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.cycle[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_82_clk_in_regs),
    .D(_05556_),
    .Q(\inst$top.soc.wb_to_csr.cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.cycle[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_82_clk_in_regs),
    .D(_19668_),
    .Q(\inst$top.soc.wb_to_csr.cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.cycle[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_52_clk_in_regs),
    .D(_05558_),
    .Q(\inst$top.soc.wb_to_csr.cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__ack$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk_in_regs),
    .D(_05559_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__ack ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_64_clk_in_regs),
    .D(_05560_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[0] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_69_clk_in_regs),
    .D(_05561_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[10] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_62_clk_in_regs),
    .D(_05562_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[11] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_62_clk_in_regs),
    .D(_05563_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[12] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_61_clk_in_regs),
    .D(_05564_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[13] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_67_clk_in_regs),
    .D(_05565_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[14] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_68_clk_in_regs),
    .D(_05566_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[15] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_81_clk_in_regs),
    .D(_05567_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[16] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_70_clk_in_regs),
    .D(_05568_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[17] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_69_clk_in_regs),
    .D(_05569_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[18] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_70_clk_in_regs),
    .D(_05570_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[19] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_59_clk_in_regs),
    .D(_05571_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[1] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_81_clk_in_regs),
    .D(_05572_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[20] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_52_clk_in_regs),
    .D(_05573_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[21] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_71_clk_in_regs),
    .D(_05574_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[22] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_61_clk_in_regs),
    .D(_05575_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[23] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_59_clk_in_regs),
    .D(_05576_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[24] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_59_clk_in_regs),
    .D(_05577_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[25] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_64_clk_in_regs),
    .D(_05578_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[26] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[27]$_SDFFE_PP0P_  (.CLK(clknet_leaf_63_clk_in_regs),
    .D(_05579_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[27] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_59_clk_in_regs),
    .D(_05580_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[28] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[29]$_SDFFE_PP0P_  (.CLK(clknet_leaf_59_clk_in_regs),
    .D(_05581_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[29] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_65_clk_in_regs),
    .D(_05582_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[2] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_63_clk_in_regs),
    .D(_05583_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[30] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_62_clk_in_regs),
    .D(_05584_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[31] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_65_clk_in_regs),
    .D(_05585_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[3] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_65_clk_in_regs),
    .D(_05586_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[4] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_62_clk_in_regs),
    .D(_05587_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[5] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_65_clk_in_regs),
    .D(_05588_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[6] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_65_clk_in_regs),
    .D(_05589_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[7] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_60_clk_in_regs),
    .D(_05590_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[8] ));
 sky130_fd_sc_hd__dfxtp_1 \inst$top.soc.wb_to_csr.wb_bus__dat_r[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_53_clk_in_regs),
    .D(_05591_),
    .Q(\inst$top.soc.wb_to_csr.wb_bus__dat_r[9] ));
 sky130_fd_sc_hd__conb_1 _43885__1 (.LO(gpio_analog_en[0]));
 sky130_fd_sc_hd__conb_1 _43886__2 (.LO(gpio_analog_en[1]));
 sky130_fd_sc_hd__conb_1 _43887__3 (.LO(gpio_analog_en[2]));
 sky130_fd_sc_hd__conb_1 _43888__4 (.LO(gpio_analog_en[3]));
 sky130_fd_sc_hd__conb_1 _43889__5 (.LO(gpio_analog_en[4]));
 sky130_fd_sc_hd__conb_1 _43890__6 (.LO(gpio_analog_en[5]));
 sky130_fd_sc_hd__conb_1 _43891__7 (.LO(gpio_analog_en[6]));
 sky130_fd_sc_hd__conb_1 _43892__8 (.LO(gpio_analog_en[7]));
 sky130_fd_sc_hd__conb_1 _43893__9 (.LO(gpio_analog_en[8]));
 sky130_fd_sc_hd__conb_1 _43894__10 (.LO(gpio_analog_en[9]));
 sky130_fd_sc_hd__conb_1 _43895__11 (.LO(gpio_analog_en[10]));
 sky130_fd_sc_hd__conb_1 _43896__12 (.LO(gpio_analog_en[11]));
 sky130_fd_sc_hd__conb_1 _43897__13 (.LO(gpio_analog_en[12]));
 sky130_fd_sc_hd__conb_1 _43898__14 (.LO(gpio_analog_en[13]));
 sky130_fd_sc_hd__conb_1 _43899__15 (.LO(gpio_analog_en[14]));
 sky130_fd_sc_hd__conb_1 _43900__16 (.LO(gpio_analog_en[15]));
 sky130_fd_sc_hd__conb_1 _43901__17 (.LO(gpio_analog_en[16]));
 sky130_fd_sc_hd__conb_1 _43902__18 (.LO(gpio_analog_en[17]));
 sky130_fd_sc_hd__conb_1 _43903__19 (.LO(gpio_analog_en[18]));
 sky130_fd_sc_hd__conb_1 _43904__20 (.LO(gpio_analog_en[19]));
 sky130_fd_sc_hd__conb_1 _43905__21 (.LO(gpio_analog_en[20]));
 sky130_fd_sc_hd__conb_1 _43906__22 (.LO(gpio_analog_en[21]));
 sky130_fd_sc_hd__conb_1 _43907__23 (.LO(gpio_analog_en[22]));
 sky130_fd_sc_hd__conb_1 _43908__24 (.LO(gpio_analog_en[23]));
 sky130_fd_sc_hd__conb_1 _43909__25 (.LO(gpio_analog_en[24]));
 sky130_fd_sc_hd__conb_1 _43910__26 (.LO(gpio_analog_en[25]));
 sky130_fd_sc_hd__conb_1 _43911__27 (.LO(gpio_analog_en[26]));
 sky130_fd_sc_hd__conb_1 _43912__28 (.LO(gpio_analog_en[27]));
 sky130_fd_sc_hd__conb_1 _43913__29 (.LO(gpio_analog_en[28]));
 sky130_fd_sc_hd__conb_1 _43914__30 (.LO(gpio_analog_en[29]));
 sky130_fd_sc_hd__conb_1 _43915__31 (.LO(gpio_analog_en[30]));
 sky130_fd_sc_hd__conb_1 _43916__32 (.LO(gpio_analog_en[31]));
 sky130_fd_sc_hd__conb_1 _43917__33 (.LO(gpio_analog_en[32]));
 sky130_fd_sc_hd__conb_1 _43918__34 (.LO(gpio_analog_en[33]));
 sky130_fd_sc_hd__conb_1 _43919__35 (.LO(gpio_analog_en[34]));
 sky130_fd_sc_hd__conb_1 _43920__36 (.LO(gpio_analog_en[35]));
 sky130_fd_sc_hd__conb_1 _43921__37 (.LO(gpio_analog_en[36]));
 sky130_fd_sc_hd__conb_1 _43922__38 (.LO(gpio_analog_en[37]));
 sky130_fd_sc_hd__conb_1 _43923__39 (.LO(gpio_analog_en[38]));
 sky130_fd_sc_hd__conb_1 _43924__40 (.LO(gpio_analog_en[39]));
 sky130_fd_sc_hd__conb_1 _43925__41 (.LO(gpio_analog_en[40]));
 sky130_fd_sc_hd__conb_1 _43926__42 (.LO(gpio_analog_en[41]));
 sky130_fd_sc_hd__conb_1 _43927__43 (.LO(gpio_analog_en[42]));
 sky130_fd_sc_hd__conb_1 _43928__44 (.LO(gpio_analog_en[43]));
 sky130_fd_sc_hd__conb_1 _43929__45 (.LO(gpio_analog_pol[0]));
 sky130_fd_sc_hd__conb_1 _43930__46 (.LO(gpio_analog_pol[1]));
 sky130_fd_sc_hd__conb_1 _43931__47 (.LO(gpio_analog_pol[2]));
 sky130_fd_sc_hd__conb_1 _43932__48 (.LO(gpio_analog_pol[3]));
 sky130_fd_sc_hd__conb_1 _43933__49 (.LO(gpio_analog_pol[4]));
 sky130_fd_sc_hd__conb_1 _43934__50 (.LO(gpio_analog_pol[5]));
 sky130_fd_sc_hd__conb_1 _43935__51 (.LO(gpio_analog_pol[6]));
 sky130_fd_sc_hd__conb_1 _43936__52 (.LO(gpio_analog_pol[7]));
 sky130_fd_sc_hd__conb_1 _43937__53 (.LO(gpio_analog_pol[8]));
 sky130_fd_sc_hd__conb_1 _43938__54 (.LO(gpio_analog_pol[9]));
 sky130_fd_sc_hd__conb_1 _43939__55 (.LO(gpio_analog_pol[10]));
 sky130_fd_sc_hd__conb_1 _43940__56 (.LO(gpio_analog_pol[11]));
 sky130_fd_sc_hd__conb_1 _43941__57 (.LO(gpio_analog_pol[12]));
 sky130_fd_sc_hd__conb_1 _43942__58 (.LO(gpio_analog_pol[13]));
 sky130_fd_sc_hd__conb_1 _43943__59 (.LO(gpio_analog_pol[14]));
 sky130_fd_sc_hd__conb_1 _43944__60 (.LO(gpio_analog_pol[15]));
 sky130_fd_sc_hd__conb_1 _43945__61 (.LO(gpio_analog_pol[16]));
 sky130_fd_sc_hd__conb_1 _43946__62 (.LO(gpio_analog_pol[17]));
 sky130_fd_sc_hd__conb_1 _43947__63 (.LO(gpio_analog_pol[18]));
 sky130_fd_sc_hd__conb_1 _43948__64 (.LO(gpio_analog_pol[19]));
 sky130_fd_sc_hd__conb_1 _43949__65 (.LO(gpio_analog_pol[20]));
 sky130_fd_sc_hd__conb_1 _43950__66 (.LO(gpio_analog_pol[21]));
 sky130_fd_sc_hd__conb_1 _43951__67 (.LO(gpio_analog_pol[22]));
 sky130_fd_sc_hd__conb_1 _43952__68 (.LO(gpio_analog_pol[23]));
 sky130_fd_sc_hd__conb_1 _43953__69 (.LO(gpio_analog_pol[24]));
 sky130_fd_sc_hd__conb_1 _43954__70 (.LO(gpio_analog_pol[25]));
 sky130_fd_sc_hd__conb_1 _43955__71 (.LO(gpio_analog_pol[26]));
 sky130_fd_sc_hd__conb_1 _43956__72 (.LO(gpio_analog_pol[27]));
 sky130_fd_sc_hd__conb_1 _43957__73 (.LO(gpio_analog_pol[28]));
 sky130_fd_sc_hd__conb_1 _43958__74 (.LO(gpio_analog_pol[29]));
 sky130_fd_sc_hd__conb_1 _43959__75 (.LO(gpio_analog_pol[30]));
 sky130_fd_sc_hd__conb_1 _43960__76 (.LO(gpio_analog_pol[31]));
 sky130_fd_sc_hd__conb_1 _43961__77 (.LO(gpio_analog_pol[32]));
 sky130_fd_sc_hd__conb_1 _43962__78 (.LO(gpio_analog_pol[33]));
 sky130_fd_sc_hd__conb_1 _43963__79 (.LO(gpio_analog_pol[34]));
 sky130_fd_sc_hd__conb_1 _43964__80 (.LO(gpio_analog_pol[35]));
 sky130_fd_sc_hd__conb_1 _43965__81 (.LO(gpio_analog_pol[36]));
 sky130_fd_sc_hd__conb_1 _43966__82 (.LO(gpio_analog_pol[37]));
 sky130_fd_sc_hd__conb_1 _43967__83 (.LO(gpio_analog_pol[38]));
 sky130_fd_sc_hd__conb_1 _43968__84 (.LO(gpio_analog_pol[39]));
 sky130_fd_sc_hd__conb_1 _43969__85 (.LO(gpio_analog_pol[40]));
 sky130_fd_sc_hd__conb_1 _43970__86 (.LO(gpio_analog_pol[41]));
 sky130_fd_sc_hd__conb_1 _43971__87 (.LO(gpio_analog_pol[42]));
 sky130_fd_sc_hd__conb_1 _43972__88 (.LO(gpio_analog_pol[43]));
 sky130_fd_sc_hd__conb_1 _43973__89 (.LO(gpio_analog_sel[0]));
 sky130_fd_sc_hd__conb_1 _43974__90 (.LO(gpio_analog_sel[1]));
 sky130_fd_sc_hd__conb_1 _43975__91 (.LO(gpio_analog_sel[2]));
 sky130_fd_sc_hd__conb_1 _43976__92 (.LO(gpio_analog_sel[3]));
 sky130_fd_sc_hd__conb_1 _43977__93 (.LO(gpio_analog_sel[4]));
 sky130_fd_sc_hd__conb_1 _43978__94 (.LO(gpio_analog_sel[5]));
 sky130_fd_sc_hd__conb_1 _43979__95 (.LO(gpio_analog_sel[6]));
 sky130_fd_sc_hd__conb_1 _43980__96 (.LO(gpio_analog_sel[7]));
 sky130_fd_sc_hd__conb_1 _43981__97 (.LO(gpio_analog_sel[8]));
 sky130_fd_sc_hd__conb_1 _43982__98 (.LO(gpio_analog_sel[9]));
 sky130_fd_sc_hd__conb_1 _43983__99 (.LO(gpio_analog_sel[10]));
 sky130_fd_sc_hd__conb_1 _43984__100 (.LO(gpio_analog_sel[11]));
 sky130_fd_sc_hd__conb_1 _43985__101 (.LO(gpio_analog_sel[12]));
 sky130_fd_sc_hd__conb_1 _43986__102 (.LO(gpio_analog_sel[13]));
 sky130_fd_sc_hd__conb_1 _43987__103 (.LO(gpio_analog_sel[14]));
 sky130_fd_sc_hd__conb_1 _43988__104 (.LO(gpio_analog_sel[15]));
 sky130_fd_sc_hd__conb_1 _43989__105 (.LO(gpio_analog_sel[16]));
 sky130_fd_sc_hd__conb_1 _43990__106 (.LO(gpio_analog_sel[17]));
 sky130_fd_sc_hd__conb_1 _43991__107 (.LO(gpio_analog_sel[18]));
 sky130_fd_sc_hd__conb_1 _43992__108 (.LO(gpio_analog_sel[19]));
 sky130_fd_sc_hd__conb_1 _43993__109 (.LO(gpio_analog_sel[20]));
 sky130_fd_sc_hd__conb_1 _43994__110 (.LO(gpio_analog_sel[21]));
 sky130_fd_sc_hd__conb_1 _43995__111 (.LO(gpio_analog_sel[22]));
 sky130_fd_sc_hd__conb_1 _43996__112 (.LO(gpio_analog_sel[23]));
 sky130_fd_sc_hd__conb_1 _43997__113 (.LO(gpio_analog_sel[24]));
 sky130_fd_sc_hd__conb_1 _43998__114 (.LO(gpio_analog_sel[25]));
 sky130_fd_sc_hd__conb_1 _43999__115 (.LO(gpio_analog_sel[26]));
 sky130_fd_sc_hd__conb_1 _44000__116 (.LO(gpio_analog_sel[27]));
 sky130_fd_sc_hd__conb_1 _44001__117 (.LO(gpio_analog_sel[28]));
 sky130_fd_sc_hd__conb_1 _44002__118 (.LO(gpio_analog_sel[29]));
 sky130_fd_sc_hd__conb_1 _44003__119 (.LO(gpio_analog_sel[30]));
 sky130_fd_sc_hd__conb_1 _44004__120 (.LO(gpio_analog_sel[31]));
 sky130_fd_sc_hd__conb_1 _44005__121 (.LO(gpio_analog_sel[32]));
 sky130_fd_sc_hd__conb_1 _44006__122 (.LO(gpio_analog_sel[33]));
 sky130_fd_sc_hd__conb_1 _44007__123 (.LO(gpio_analog_sel[34]));
 sky130_fd_sc_hd__conb_1 _44008__124 (.LO(gpio_analog_sel[35]));
 sky130_fd_sc_hd__conb_1 _44009__125 (.LO(gpio_analog_sel[36]));
 sky130_fd_sc_hd__conb_1 _44010__126 (.LO(gpio_analog_sel[37]));
 sky130_fd_sc_hd__conb_1 _44011__127 (.LO(gpio_analog_sel[38]));
 sky130_fd_sc_hd__conb_1 _44012__128 (.LO(gpio_analog_sel[39]));
 sky130_fd_sc_hd__conb_1 _44013__129 (.LO(gpio_analog_sel[40]));
 sky130_fd_sc_hd__conb_1 _44014__130 (.LO(gpio_analog_sel[41]));
 sky130_fd_sc_hd__conb_1 _44015__131 (.LO(gpio_analog_sel[42]));
 sky130_fd_sc_hd__conb_1 _44016__132 (.LO(gpio_analog_sel[43]));
 sky130_fd_sc_hd__conb_1 _44024__133 (.LO(gpio_dm0[7]));
 sky130_fd_sc_hd__conb_1 _44033__134 (.LO(gpio_dm0[16]));
 sky130_fd_sc_hd__conb_1 _44034__135 (.LO(gpio_dm0[17]));
 sky130_fd_sc_hd__conb_1 _44035__136 (.LO(gpio_dm0[18]));
 sky130_fd_sc_hd__conb_1 _44036__137 (.LO(gpio_dm0[19]));
 sky130_fd_sc_hd__conb_1 _44037__138 (.LO(gpio_dm0[20]));
 sky130_fd_sc_hd__conb_1 _44038__139 (.LO(gpio_dm0[21]));
 sky130_fd_sc_hd__conb_1 _44039__140 (.LO(gpio_dm0[22]));
 sky130_fd_sc_hd__conb_1 _44040__141 (.LO(gpio_dm0[23]));
 sky130_fd_sc_hd__conb_1 _44041__142 (.LO(gpio_dm0[24]));
 sky130_fd_sc_hd__conb_1 _44046__143 (.LO(gpio_dm0[29]));
 sky130_fd_sc_hd__conb_1 _44047__144 (.LO(gpio_dm0[30]));
 sky130_fd_sc_hd__conb_1 _44048__145 (.LO(gpio_dm0[31]));
 sky130_fd_sc_hd__conb_1 _44049__146 (.LO(gpio_dm0[32]));
 sky130_fd_sc_hd__conb_1 _44050__147 (.LO(gpio_dm0[33]));
 sky130_fd_sc_hd__conb_1 _44051__148 (.LO(gpio_dm0[34]));
 sky130_fd_sc_hd__conb_1 _44052__149 (.LO(gpio_dm0[35]));
 sky130_fd_sc_hd__conb_1 _44053__150 (.LO(gpio_dm0[36]));
 sky130_fd_sc_hd__conb_1 _44054__151 (.LO(gpio_dm0[37]));
 sky130_fd_sc_hd__conb_1 _44055__152 (.LO(gpio_dm0[38]));
 sky130_fd_sc_hd__conb_1 _44056__153 (.LO(gpio_dm0[39]));
 sky130_fd_sc_hd__conb_1 _44057__154 (.LO(gpio_dm0[40]));
 sky130_fd_sc_hd__conb_1 _44058__155 (.LO(gpio_dm0[41]));
 sky130_fd_sc_hd__conb_1 _44059__156 (.LO(gpio_dm0[42]));
 sky130_fd_sc_hd__conb_1 _44060__157 (.LO(gpio_dm0[43]));
 sky130_fd_sc_hd__conb_1 _44068__158 (.LO(gpio_dm1[7]));
 sky130_fd_sc_hd__conb_1 _44077__159 (.LO(gpio_dm1[16]));
 sky130_fd_sc_hd__conb_1 _44078__160 (.LO(gpio_dm1[17]));
 sky130_fd_sc_hd__conb_1 _44079__161 (.LO(gpio_dm1[18]));
 sky130_fd_sc_hd__conb_1 _44080__162 (.LO(gpio_dm1[19]));
 sky130_fd_sc_hd__conb_1 _44081__163 (.LO(gpio_dm1[20]));
 sky130_fd_sc_hd__conb_1 _44082__164 (.LO(gpio_dm1[21]));
 sky130_fd_sc_hd__conb_1 _44083__165 (.LO(gpio_dm1[22]));
 sky130_fd_sc_hd__conb_1 _44084__166 (.LO(gpio_dm1[23]));
 sky130_fd_sc_hd__conb_1 _44085__167 (.LO(gpio_dm1[24]));
 sky130_fd_sc_hd__conb_1 _44090__168 (.LO(gpio_dm1[29]));
 sky130_fd_sc_hd__conb_1 _44091__169 (.LO(gpio_dm1[30]));
 sky130_fd_sc_hd__conb_1 _44092__170 (.LO(gpio_dm1[31]));
 sky130_fd_sc_hd__conb_1 _44093__171 (.LO(gpio_dm1[32]));
 sky130_fd_sc_hd__conb_1 _44094__172 (.LO(gpio_dm1[33]));
 sky130_fd_sc_hd__conb_1 _44095__173 (.LO(gpio_dm1[34]));
 sky130_fd_sc_hd__conb_1 _44096__174 (.LO(gpio_dm1[35]));
 sky130_fd_sc_hd__conb_1 _44097__175 (.LO(gpio_dm1[36]));
 sky130_fd_sc_hd__conb_1 _44098__176 (.LO(gpio_dm1[37]));
 sky130_fd_sc_hd__conb_1 _44099__177 (.LO(gpio_dm1[38]));
 sky130_fd_sc_hd__conb_1 _44100__178 (.LO(gpio_dm1[39]));
 sky130_fd_sc_hd__conb_1 _44101__179 (.LO(gpio_dm1[40]));
 sky130_fd_sc_hd__conb_1 _44102__180 (.LO(gpio_dm1[41]));
 sky130_fd_sc_hd__conb_1 _44103__181 (.LO(gpio_dm1[42]));
 sky130_fd_sc_hd__conb_1 _44104__182 (.LO(gpio_dm1[43]));
 sky130_fd_sc_hd__conb_1 _44105__183 (.LO(gpio_dm2[0]));
 sky130_fd_sc_hd__conb_1 _44106__184 (.LO(gpio_dm2[1]));
 sky130_fd_sc_hd__conb_1 _44107__185 (.LO(gpio_dm2[2]));
 sky130_fd_sc_hd__conb_1 _44108__186 (.LO(gpio_dm2[3]));
 sky130_fd_sc_hd__conb_1 _44109__187 (.LO(gpio_dm2[4]));
 sky130_fd_sc_hd__conb_1 _44110__188 (.LO(gpio_dm2[5]));
 sky130_fd_sc_hd__conb_1 _44111__189 (.LO(gpio_dm2[6]));
 sky130_fd_sc_hd__conb_1 _44112__190 (.LO(gpio_dm2[7]));
 sky130_fd_sc_hd__conb_1 _44113__191 (.LO(gpio_dm2[8]));
 sky130_fd_sc_hd__conb_1 _44114__192 (.LO(gpio_dm2[9]));
 sky130_fd_sc_hd__conb_1 _44115__193 (.LO(gpio_dm2[10]));
 sky130_fd_sc_hd__conb_1 _44116__194 (.LO(gpio_dm2[11]));
 sky130_fd_sc_hd__conb_1 _44117__195 (.LO(gpio_dm2[12]));
 sky130_fd_sc_hd__conb_1 _44118__196 (.LO(gpio_dm2[13]));
 sky130_fd_sc_hd__conb_1 _44119__197 (.LO(gpio_dm2[14]));
 sky130_fd_sc_hd__conb_1 _44120__198 (.LO(gpio_dm2[15]));
 sky130_fd_sc_hd__conb_1 _44121__199 (.LO(gpio_dm2[16]));
 sky130_fd_sc_hd__conb_1 _44122__200 (.LO(gpio_dm2[17]));
 sky130_fd_sc_hd__conb_1 _44123__201 (.LO(gpio_dm2[18]));
 sky130_fd_sc_hd__conb_1 _44124__202 (.LO(gpio_dm2[19]));
 sky130_fd_sc_hd__conb_1 _44125__203 (.LO(gpio_dm2[20]));
 sky130_fd_sc_hd__conb_1 _44126__204 (.LO(gpio_dm2[21]));
 sky130_fd_sc_hd__conb_1 _44127__205 (.LO(gpio_dm2[22]));
 sky130_fd_sc_hd__conb_1 _44128__206 (.LO(gpio_dm2[23]));
 sky130_fd_sc_hd__conb_1 _44129__207 (.LO(gpio_dm2[24]));
 sky130_fd_sc_hd__conb_1 _44130__208 (.LO(gpio_dm2[25]));
 sky130_fd_sc_hd__conb_1 _44131__209 (.LO(gpio_dm2[26]));
 sky130_fd_sc_hd__conb_1 _44132__210 (.LO(gpio_dm2[27]));
 sky130_fd_sc_hd__conb_1 _44133__211 (.LO(gpio_dm2[28]));
 sky130_fd_sc_hd__conb_1 _44134__212 (.LO(gpio_dm2[29]));
 sky130_fd_sc_hd__conb_1 _44135__213 (.LO(gpio_dm2[30]));
 sky130_fd_sc_hd__conb_1 _44136__214 (.LO(gpio_dm2[31]));
 sky130_fd_sc_hd__conb_1 _44137__215 (.LO(gpio_dm2[32]));
 sky130_fd_sc_hd__conb_1 _44138__216 (.LO(gpio_dm2[33]));
 sky130_fd_sc_hd__conb_1 _44139__217 (.LO(gpio_dm2[34]));
 sky130_fd_sc_hd__conb_1 _44140__218 (.LO(gpio_dm2[35]));
 sky130_fd_sc_hd__conb_1 _44141__219 (.LO(gpio_dm2[36]));
 sky130_fd_sc_hd__conb_1 _44142__220 (.LO(gpio_dm2[37]));
 sky130_fd_sc_hd__conb_1 _44143__221 (.LO(gpio_dm2[38]));
 sky130_fd_sc_hd__conb_1 _44144__222 (.LO(gpio_dm2[39]));
 sky130_fd_sc_hd__conb_1 _44145__223 (.LO(gpio_dm2[40]));
 sky130_fd_sc_hd__conb_1 _44146__224 (.LO(gpio_dm2[41]));
 sky130_fd_sc_hd__conb_1 _44147__225 (.LO(gpio_dm2[42]));
 sky130_fd_sc_hd__conb_1 _44148__226 (.LO(gpio_dm2[43]));
 sky130_fd_sc_hd__conb_1 _44149__227 (.LO(gpio_holdover[0]));
 sky130_fd_sc_hd__conb_1 _44150__228 (.LO(gpio_holdover[1]));
 sky130_fd_sc_hd__conb_1 _44151__229 (.LO(gpio_holdover[2]));
 sky130_fd_sc_hd__conb_1 _44152__230 (.LO(gpio_holdover[3]));
 sky130_fd_sc_hd__conb_1 _44153__231 (.LO(gpio_holdover[4]));
 sky130_fd_sc_hd__conb_1 _44154__232 (.LO(gpio_holdover[5]));
 sky130_fd_sc_hd__conb_1 _44155__233 (.LO(gpio_holdover[6]));
 sky130_fd_sc_hd__conb_1 _44156__234 (.LO(gpio_holdover[7]));
 sky130_fd_sc_hd__conb_1 _44157__235 (.LO(gpio_holdover[8]));
 sky130_fd_sc_hd__conb_1 _44158__236 (.LO(gpio_holdover[9]));
 sky130_fd_sc_hd__conb_1 _44159__237 (.LO(gpio_holdover[10]));
 sky130_fd_sc_hd__conb_1 _44160__238 (.LO(gpio_holdover[11]));
 sky130_fd_sc_hd__conb_1 _44161__239 (.LO(gpio_holdover[12]));
 sky130_fd_sc_hd__conb_1 _44162__240 (.LO(gpio_holdover[13]));
 sky130_fd_sc_hd__conb_1 _44163__241 (.LO(gpio_holdover[14]));
 sky130_fd_sc_hd__conb_1 _44164__242 (.LO(gpio_holdover[15]));
 sky130_fd_sc_hd__conb_1 _44165__243 (.LO(gpio_holdover[16]));
 sky130_fd_sc_hd__conb_1 _44166__244 (.LO(gpio_holdover[17]));
 sky130_fd_sc_hd__conb_1 _44167__245 (.LO(gpio_holdover[18]));
 sky130_fd_sc_hd__conb_1 _44168__246 (.LO(gpio_holdover[19]));
 sky130_fd_sc_hd__conb_1 _44169__247 (.LO(gpio_holdover[20]));
 sky130_fd_sc_hd__conb_1 _44170__248 (.LO(gpio_holdover[21]));
 sky130_fd_sc_hd__conb_1 _44171__249 (.LO(gpio_holdover[22]));
 sky130_fd_sc_hd__conb_1 _44172__250 (.LO(gpio_holdover[23]));
 sky130_fd_sc_hd__conb_1 _44173__251 (.LO(gpio_holdover[24]));
 sky130_fd_sc_hd__conb_1 _44174__252 (.LO(gpio_holdover[25]));
 sky130_fd_sc_hd__conb_1 _44175__253 (.LO(gpio_holdover[26]));
 sky130_fd_sc_hd__conb_1 _44176__254 (.LO(gpio_holdover[27]));
 sky130_fd_sc_hd__conb_1 _44177__255 (.LO(gpio_holdover[28]));
 sky130_fd_sc_hd__conb_1 _44178__256 (.LO(gpio_holdover[29]));
 sky130_fd_sc_hd__conb_1 _44179__257 (.LO(gpio_holdover[30]));
 sky130_fd_sc_hd__conb_1 _44180__258 (.LO(gpio_holdover[31]));
 sky130_fd_sc_hd__conb_1 _44181__259 (.LO(gpio_holdover[32]));
 sky130_fd_sc_hd__conb_1 _44182__260 (.LO(gpio_holdover[33]));
 sky130_fd_sc_hd__conb_1 _44183__261 (.LO(gpio_holdover[34]));
 sky130_fd_sc_hd__conb_1 _44184__262 (.LO(gpio_holdover[35]));
 sky130_fd_sc_hd__conb_1 _44185__263 (.LO(gpio_holdover[36]));
 sky130_fd_sc_hd__conb_1 _44186__264 (.LO(gpio_holdover[37]));
 sky130_fd_sc_hd__conb_1 _44187__265 (.LO(gpio_holdover[38]));
 sky130_fd_sc_hd__conb_1 _44188__266 (.LO(gpio_holdover[39]));
 sky130_fd_sc_hd__conb_1 _44189__267 (.LO(gpio_holdover[40]));
 sky130_fd_sc_hd__conb_1 _44190__268 (.LO(gpio_holdover[41]));
 sky130_fd_sc_hd__conb_1 _44191__269 (.LO(gpio_holdover[42]));
 sky130_fd_sc_hd__conb_1 _44192__270 (.LO(gpio_holdover[43]));
 sky130_fd_sc_hd__conb_1 _44193__271 (.LO(gpio_ib_mode_sel[0]));
 sky130_fd_sc_hd__conb_1 _44194__272 (.LO(gpio_ib_mode_sel[1]));
 sky130_fd_sc_hd__conb_1 _44195__273 (.LO(gpio_ib_mode_sel[2]));
 sky130_fd_sc_hd__conb_1 _44196__274 (.LO(gpio_ib_mode_sel[3]));
 sky130_fd_sc_hd__conb_1 _44197__275 (.LO(gpio_ib_mode_sel[4]));
 sky130_fd_sc_hd__conb_1 _44198__276 (.LO(gpio_ib_mode_sel[5]));
 sky130_fd_sc_hd__conb_1 _44199__277 (.LO(gpio_ib_mode_sel[6]));
 sky130_fd_sc_hd__conb_1 _44200__278 (.LO(gpio_ib_mode_sel[7]));
 sky130_fd_sc_hd__conb_1 _44201__279 (.LO(gpio_ib_mode_sel[8]));
 sky130_fd_sc_hd__conb_1 _44202__280 (.LO(gpio_ib_mode_sel[9]));
 sky130_fd_sc_hd__conb_1 _44203__281 (.LO(gpio_ib_mode_sel[10]));
 sky130_fd_sc_hd__conb_1 _44204__282 (.LO(gpio_ib_mode_sel[11]));
 sky130_fd_sc_hd__conb_1 _44205__283 (.LO(gpio_ib_mode_sel[12]));
 sky130_fd_sc_hd__conb_1 _44206__284 (.LO(gpio_ib_mode_sel[13]));
 sky130_fd_sc_hd__conb_1 _44207__285 (.LO(gpio_ib_mode_sel[14]));
 sky130_fd_sc_hd__conb_1 _44208__286 (.LO(gpio_ib_mode_sel[15]));
 sky130_fd_sc_hd__conb_1 _44209__287 (.LO(gpio_ib_mode_sel[16]));
 sky130_fd_sc_hd__conb_1 _44210__288 (.LO(gpio_ib_mode_sel[17]));
 sky130_fd_sc_hd__conb_1 _44211__289 (.LO(gpio_ib_mode_sel[18]));
 sky130_fd_sc_hd__conb_1 _44212__290 (.LO(gpio_ib_mode_sel[19]));
 sky130_fd_sc_hd__conb_1 _44213__291 (.LO(gpio_ib_mode_sel[20]));
 sky130_fd_sc_hd__conb_1 _44214__292 (.LO(gpio_ib_mode_sel[21]));
 sky130_fd_sc_hd__conb_1 _44215__293 (.LO(gpio_ib_mode_sel[22]));
 sky130_fd_sc_hd__conb_1 _44216__294 (.LO(gpio_ib_mode_sel[23]));
 sky130_fd_sc_hd__conb_1 _44217__295 (.LO(gpio_ib_mode_sel[24]));
 sky130_fd_sc_hd__conb_1 _44218__296 (.LO(gpio_ib_mode_sel[25]));
 sky130_fd_sc_hd__conb_1 _44219__297 (.LO(gpio_ib_mode_sel[26]));
 sky130_fd_sc_hd__conb_1 _44220__298 (.LO(gpio_ib_mode_sel[27]));
 sky130_fd_sc_hd__conb_1 _44221__299 (.LO(gpio_ib_mode_sel[28]));
 sky130_fd_sc_hd__conb_1 _44222__300 (.LO(gpio_ib_mode_sel[29]));
 sky130_fd_sc_hd__conb_1 _44223__301 (.LO(gpio_ib_mode_sel[30]));
 sky130_fd_sc_hd__conb_1 _44224__302 (.LO(gpio_ib_mode_sel[31]));
 sky130_fd_sc_hd__conb_1 _44225__303 (.LO(gpio_ib_mode_sel[32]));
 sky130_fd_sc_hd__conb_1 _44226__304 (.LO(gpio_ib_mode_sel[33]));
 sky130_fd_sc_hd__conb_1 _44227__305 (.LO(gpio_ib_mode_sel[34]));
 sky130_fd_sc_hd__conb_1 _44228__306 (.LO(gpio_ib_mode_sel[35]));
 sky130_fd_sc_hd__conb_1 _44229__307 (.LO(gpio_ib_mode_sel[36]));
 sky130_fd_sc_hd__conb_1 _44230__308 (.LO(gpio_ib_mode_sel[37]));
 sky130_fd_sc_hd__conb_1 _44231__309 (.LO(gpio_ib_mode_sel[38]));
 sky130_fd_sc_hd__conb_1 _44232__310 (.LO(gpio_ib_mode_sel[39]));
 sky130_fd_sc_hd__conb_1 _44233__311 (.LO(gpio_ib_mode_sel[40]));
 sky130_fd_sc_hd__conb_1 _44234__312 (.LO(gpio_ib_mode_sel[41]));
 sky130_fd_sc_hd__conb_1 _44235__313 (.LO(gpio_ib_mode_sel[42]));
 sky130_fd_sc_hd__conb_1 _44236__314 (.LO(gpio_ib_mode_sel[43]));
 sky130_fd_sc_hd__conb_1 _44244__315 (.LO(gpio_inp_dis[7]));
 sky130_fd_sc_hd__conb_1 _44275__316 (.LO(gpio_inp_dis[38]));
 sky130_fd_sc_hd__conb_1 _44277__317 (.LO(gpio_inp_dis[40]));
 sky130_fd_sc_hd__conb_1 _44281__318 (.LO(gpio_oeb[0]));
 sky130_fd_sc_hd__conb_1 _44282__319 (.LO(gpio_oeb[1]));
 sky130_fd_sc_hd__conb_1 _44287__320 (.LO(gpio_oeb[6]));
 sky130_fd_sc_hd__conb_1 _44332__321 (.LO(gpio_out[7]));
 sky130_fd_sc_hd__conb_1 _44341__322 (.LO(gpio_out[16]));
 sky130_fd_sc_hd__conb_1 _44342__323 (.LO(gpio_out[17]));
 sky130_fd_sc_hd__conb_1 _44343__324 (.LO(gpio_out[18]));
 sky130_fd_sc_hd__conb_1 _44344__325 (.LO(gpio_out[19]));
 sky130_fd_sc_hd__conb_1 _44345__326 (.LO(gpio_out[20]));
 sky130_fd_sc_hd__conb_1 _44346__327 (.LO(gpio_out[21]));
 sky130_fd_sc_hd__conb_1 _44347__328 (.LO(gpio_out[22]));
 sky130_fd_sc_hd__conb_1 _44348__329 (.LO(gpio_out[23]));
 sky130_fd_sc_hd__conb_1 _44349__330 (.LO(gpio_out[24]));
 sky130_fd_sc_hd__conb_1 _44354__331 (.LO(gpio_out[29]));
 sky130_fd_sc_hd__conb_1 _44355__332 (.LO(gpio_out[30]));
 sky130_fd_sc_hd__conb_1 _44356__333 (.LO(gpio_out[31]));
 sky130_fd_sc_hd__conb_1 _44357__334 (.LO(gpio_out[32]));
 sky130_fd_sc_hd__conb_1 _44358__335 (.LO(gpio_out[33]));
 sky130_fd_sc_hd__conb_1 _44359__336 (.LO(gpio_out[34]));
 sky130_fd_sc_hd__conb_1 _44360__337 (.LO(gpio_out[35]));
 sky130_fd_sc_hd__conb_1 _44361__338 (.LO(gpio_out[36]));
 sky130_fd_sc_hd__conb_1 _44362__339 (.LO(gpio_out[37]));
 sky130_fd_sc_hd__conb_1 _44363__340 (.LO(gpio_out[38]));
 sky130_fd_sc_hd__conb_1 _44364__341 (.LO(gpio_out[39]));
 sky130_fd_sc_hd__conb_1 _44365__342 (.LO(gpio_out[40]));
 sky130_fd_sc_hd__conb_1 _44366__343 (.LO(gpio_out[41]));
 sky130_fd_sc_hd__conb_1 _44367__344 (.LO(gpio_out[42]));
 sky130_fd_sc_hd__conb_1 _44368__345 (.LO(gpio_out[43]));
 sky130_fd_sc_hd__conb_1 _44369__346 (.LO(gpio_slow_sel[0]));
 sky130_fd_sc_hd__conb_1 _44370__347 (.LO(gpio_slow_sel[1]));
 sky130_fd_sc_hd__conb_1 _44371__348 (.LO(gpio_slow_sel[2]));
 sky130_fd_sc_hd__conb_1 _44372__349 (.LO(gpio_slow_sel[3]));
 sky130_fd_sc_hd__conb_1 _44373__350 (.LO(gpio_slow_sel[4]));
 sky130_fd_sc_hd__conb_1 _44374__351 (.LO(gpio_slow_sel[5]));
 sky130_fd_sc_hd__conb_1 _44375__352 (.LO(gpio_slow_sel[6]));
 sky130_fd_sc_hd__conb_1 _44376__353 (.LO(gpio_slow_sel[7]));
 sky130_fd_sc_hd__conb_1 _44377__354 (.LO(gpio_slow_sel[8]));
 sky130_fd_sc_hd__conb_1 _44378__355 (.LO(gpio_slow_sel[9]));
 sky130_fd_sc_hd__conb_1 _44379__356 (.LO(gpio_slow_sel[10]));
 sky130_fd_sc_hd__conb_1 _44380__357 (.LO(gpio_slow_sel[11]));
 sky130_fd_sc_hd__conb_1 _44381__358 (.LO(gpio_slow_sel[12]));
 sky130_fd_sc_hd__conb_1 _44382__359 (.LO(gpio_slow_sel[13]));
 sky130_fd_sc_hd__conb_1 _44383__360 (.LO(gpio_slow_sel[14]));
 sky130_fd_sc_hd__conb_1 _44384__361 (.LO(gpio_slow_sel[15]));
 sky130_fd_sc_hd__conb_1 _44385__362 (.LO(gpio_slow_sel[16]));
 sky130_fd_sc_hd__conb_1 _44386__363 (.LO(gpio_slow_sel[17]));
 sky130_fd_sc_hd__conb_1 _44387__364 (.LO(gpio_slow_sel[18]));
 sky130_fd_sc_hd__conb_1 _44388__365 (.LO(gpio_slow_sel[19]));
 sky130_fd_sc_hd__conb_1 _44389__366 (.LO(gpio_slow_sel[20]));
 sky130_fd_sc_hd__conb_1 _44390__367 (.LO(gpio_slow_sel[21]));
 sky130_fd_sc_hd__conb_1 _44391__368 (.LO(gpio_slow_sel[22]));
 sky130_fd_sc_hd__conb_1 _44392__369 (.LO(gpio_slow_sel[23]));
 sky130_fd_sc_hd__conb_1 _44393__370 (.LO(gpio_slow_sel[24]));
 sky130_fd_sc_hd__conb_1 _44394__371 (.LO(gpio_slow_sel[25]));
 sky130_fd_sc_hd__conb_1 _44395__372 (.LO(gpio_slow_sel[26]));
 sky130_fd_sc_hd__conb_1 _44396__373 (.LO(gpio_slow_sel[27]));
 sky130_fd_sc_hd__conb_1 _44397__374 (.LO(gpio_slow_sel[28]));
 sky130_fd_sc_hd__conb_1 _44398__375 (.LO(gpio_slow_sel[29]));
 sky130_fd_sc_hd__conb_1 _44399__376 (.LO(gpio_slow_sel[30]));
 sky130_fd_sc_hd__conb_1 _44400__377 (.LO(gpio_slow_sel[31]));
 sky130_fd_sc_hd__conb_1 _44401__378 (.LO(gpio_slow_sel[32]));
 sky130_fd_sc_hd__conb_1 _44402__379 (.LO(gpio_slow_sel[33]));
 sky130_fd_sc_hd__conb_1 _44403__380 (.LO(gpio_slow_sel[34]));
 sky130_fd_sc_hd__conb_1 _44404__381 (.LO(gpio_slow_sel[35]));
 sky130_fd_sc_hd__conb_1 _44405__382 (.LO(gpio_slow_sel[36]));
 sky130_fd_sc_hd__conb_1 _44406__383 (.LO(gpio_slow_sel[37]));
 sky130_fd_sc_hd__conb_1 _44407__384 (.LO(gpio_slow_sel[38]));
 sky130_fd_sc_hd__conb_1 _44408__385 (.LO(gpio_slow_sel[39]));
 sky130_fd_sc_hd__conb_1 _44409__386 (.LO(gpio_slow_sel[40]));
 sky130_fd_sc_hd__conb_1 _44410__387 (.LO(gpio_slow_sel[41]));
 sky130_fd_sc_hd__conb_1 _44411__388 (.LO(gpio_slow_sel[42]));
 sky130_fd_sc_hd__conb_1 _44412__389 (.LO(gpio_slow_sel[43]));
 sky130_fd_sc_hd__conb_1 _44413__390 (.LO(gpio_vtrip_sel[0]));
 sky130_fd_sc_hd__conb_1 _44414__391 (.LO(gpio_vtrip_sel[1]));
 sky130_fd_sc_hd__conb_1 _44415__392 (.LO(gpio_vtrip_sel[2]));
 sky130_fd_sc_hd__conb_1 _44416__393 (.LO(gpio_vtrip_sel[3]));
 sky130_fd_sc_hd__conb_1 _44417__394 (.LO(gpio_vtrip_sel[4]));
 sky130_fd_sc_hd__conb_1 _44418__395 (.LO(gpio_vtrip_sel[5]));
 sky130_fd_sc_hd__conb_1 _44419__396 (.LO(gpio_vtrip_sel[6]));
 sky130_fd_sc_hd__conb_1 _44420__397 (.LO(gpio_vtrip_sel[7]));
 sky130_fd_sc_hd__conb_1 _44421__398 (.LO(gpio_vtrip_sel[8]));
 sky130_fd_sc_hd__conb_1 _44422__399 (.LO(gpio_vtrip_sel[9]));
 sky130_fd_sc_hd__conb_1 _44423__400 (.LO(gpio_vtrip_sel[10]));
 sky130_fd_sc_hd__conb_1 _44424__401 (.LO(gpio_vtrip_sel[11]));
 sky130_fd_sc_hd__conb_1 _44425__402 (.LO(gpio_vtrip_sel[12]));
 sky130_fd_sc_hd__conb_1 _44426__403 (.LO(gpio_vtrip_sel[13]));
 sky130_fd_sc_hd__conb_1 _44427__404 (.LO(gpio_vtrip_sel[14]));
 sky130_fd_sc_hd__conb_1 _44428__405 (.LO(gpio_vtrip_sel[15]));
 sky130_fd_sc_hd__conb_1 _44429__406 (.LO(gpio_vtrip_sel[16]));
 sky130_fd_sc_hd__conb_1 _44430__407 (.LO(gpio_vtrip_sel[17]));
 sky130_fd_sc_hd__conb_1 _44431__408 (.LO(gpio_vtrip_sel[18]));
 sky130_fd_sc_hd__conb_1 _44432__409 (.LO(gpio_vtrip_sel[19]));
 sky130_fd_sc_hd__conb_1 _44433__410 (.LO(gpio_vtrip_sel[20]));
 sky130_fd_sc_hd__conb_1 _44434__411 (.LO(gpio_vtrip_sel[21]));
 sky130_fd_sc_hd__conb_1 _44435__412 (.LO(gpio_vtrip_sel[22]));
 sky130_fd_sc_hd__conb_1 _44436__413 (.LO(gpio_vtrip_sel[23]));
 sky130_fd_sc_hd__conb_1 _44437__414 (.LO(gpio_vtrip_sel[24]));
 sky130_fd_sc_hd__conb_1 _44438__415 (.LO(gpio_vtrip_sel[25]));
 sky130_fd_sc_hd__conb_1 _44439__416 (.LO(gpio_vtrip_sel[26]));
 sky130_fd_sc_hd__conb_1 _44440__417 (.LO(gpio_vtrip_sel[27]));
 sky130_fd_sc_hd__conb_1 _44441__418 (.LO(gpio_vtrip_sel[28]));
 sky130_fd_sc_hd__conb_1 _44442__419 (.LO(gpio_vtrip_sel[29]));
 sky130_fd_sc_hd__conb_1 _44443__420 (.LO(gpio_vtrip_sel[30]));
 sky130_fd_sc_hd__conb_1 _44444__421 (.LO(gpio_vtrip_sel[31]));
 sky130_fd_sc_hd__conb_1 _44445__422 (.LO(gpio_vtrip_sel[32]));
 sky130_fd_sc_hd__conb_1 _44446__423 (.LO(gpio_vtrip_sel[33]));
 sky130_fd_sc_hd__conb_1 _44447__424 (.LO(gpio_vtrip_sel[34]));
 sky130_fd_sc_hd__conb_1 _44448__425 (.LO(gpio_vtrip_sel[35]));
 sky130_fd_sc_hd__conb_1 _44449__426 (.LO(gpio_vtrip_sel[36]));
 sky130_fd_sc_hd__conb_1 _44450__427 (.LO(gpio_vtrip_sel[37]));
 sky130_fd_sc_hd__conb_1 _44451__428 (.LO(gpio_vtrip_sel[38]));
 sky130_fd_sc_hd__conb_1 _44452__429 (.LO(gpio_vtrip_sel[39]));
 sky130_fd_sc_hd__conb_1 _44453__430 (.LO(gpio_vtrip_sel[40]));
 sky130_fd_sc_hd__conb_1 _44454__431 (.LO(gpio_vtrip_sel[41]));
 sky130_fd_sc_hd__conb_1 _44455__432 (.LO(gpio_vtrip_sel[42]));
 sky130_fd_sc_hd__conb_1 _44456__433 (.LO(gpio_vtrip_sel[43]));
 sky130_fd_sc_hd__conb_1 \inst$top.soc.sram.mem.0.0_434  (.LO(net433));
 sky130_fd_sc_hd__conb_1 \inst$top.soc.sram.mem.0.0_435  (.LO(net434));
 sky130_fd_sc_hd__conb_1 \inst$top.soc.sram.mem.0.0_436  (.LO(net435));
 sky130_fd_sc_hd__conb_1 \inst$top.soc.sram.mem.0.0_437  (.LO(net436));
 sky130_fd_sc_hd__conb_1 \inst$top.soc.sram.mem.0.0_438  (.LO(net437));
 sky130_fd_sc_hd__conb_1 \inst$top.soc.sram.mem.0.0_439  (.LO(net438));
 sky130_fd_sc_hd__conb_1 \inst$top.soc.sram.mem.0.0_440  (.LO(net439));
 sky130_fd_sc_hd__conb_1 \inst$top.soc.sram.mem.0.0_441  (.LO(net440));
 sky130_fd_sc_hd__conb_1 _44018__443 (.HI(gpio_dm0[1]));
 sky130_fd_sc_hd__conb_1 _44019__444 (.HI(gpio_dm0[2]));
 sky130_fd_sc_hd__conb_1 _44020__445 (.HI(gpio_dm0[3]));
 sky130_fd_sc_hd__conb_1 _44021__446 (.HI(gpio_dm0[4]));
 sky130_fd_sc_hd__conb_1 _44022__447 (.HI(gpio_dm0[5]));
 sky130_fd_sc_hd__conb_1 _44023__448 (.HI(gpio_dm0[6]));
 sky130_fd_sc_hd__conb_1 _44025__449 (.HI(gpio_dm0[8]));
 sky130_fd_sc_hd__conb_1 _44026__450 (.HI(gpio_dm0[9]));
 sky130_fd_sc_hd__conb_1 _44027__451 (.HI(gpio_dm0[10]));
 sky130_fd_sc_hd__conb_1 _44028__452 (.HI(gpio_dm0[11]));
 sky130_fd_sc_hd__conb_1 _44029__453 (.HI(gpio_dm0[12]));
 sky130_fd_sc_hd__conb_1 _44030__454 (.HI(gpio_dm0[13]));
 sky130_fd_sc_hd__conb_1 _44031__455 (.HI(gpio_dm0[14]));
 sky130_fd_sc_hd__conb_1 _44032__456 (.HI(gpio_dm0[15]));
 sky130_fd_sc_hd__conb_1 _44042__457 (.HI(gpio_dm0[25]));
 sky130_fd_sc_hd__conb_1 _44043__458 (.HI(gpio_dm0[26]));
 sky130_fd_sc_hd__conb_1 _44044__459 (.HI(gpio_dm0[27]));
 sky130_fd_sc_hd__conb_1 _44045__460 (.HI(gpio_dm0[28]));
 sky130_fd_sc_hd__conb_1 _44061__461 (.HI(gpio_dm1[0]));
 sky130_fd_sc_hd__conb_1 _44062__462 (.HI(gpio_dm1[1]));
 sky130_fd_sc_hd__conb_1 _44063__463 (.HI(gpio_dm1[2]));
 sky130_fd_sc_hd__conb_1 _44064__464 (.HI(gpio_dm1[3]));
 sky130_fd_sc_hd__conb_1 _44065__465 (.HI(gpio_dm1[4]));
 sky130_fd_sc_hd__conb_1 _44066__466 (.HI(gpio_dm1[5]));
 sky130_fd_sc_hd__conb_1 _44067__467 (.HI(gpio_dm1[6]));
 sky130_fd_sc_hd__conb_1 _44069__468 (.HI(gpio_dm1[8]));
 sky130_fd_sc_hd__conb_1 _44070__469 (.HI(gpio_dm1[9]));
 sky130_fd_sc_hd__conb_1 _44071__470 (.HI(gpio_dm1[10]));
 sky130_fd_sc_hd__conb_1 _44072__471 (.HI(gpio_dm1[11]));
 sky130_fd_sc_hd__conb_1 _44073__472 (.HI(gpio_dm1[12]));
 sky130_fd_sc_hd__conb_1 _44074__473 (.HI(gpio_dm1[13]));
 sky130_fd_sc_hd__conb_1 _44075__474 (.HI(gpio_dm1[14]));
 sky130_fd_sc_hd__conb_1 _44076__475 (.HI(gpio_dm1[15]));
 sky130_fd_sc_hd__conb_1 _44086__476 (.HI(gpio_dm1[25]));
 sky130_fd_sc_hd__conb_1 _44087__477 (.HI(gpio_dm1[26]));
 sky130_fd_sc_hd__conb_1 _44088__478 (.HI(gpio_dm1[27]));
 sky130_fd_sc_hd__conb_1 _44089__479 (.HI(gpio_dm1[28]));
 sky130_fd_sc_hd__conb_1 _44237__480 (.HI(gpio_inp_dis[0]));
 sky130_fd_sc_hd__conb_1 _44238__481 (.HI(gpio_inp_dis[1]));
 sky130_fd_sc_hd__conb_1 _44243__482 (.HI(gpio_inp_dis[6]));
 sky130_fd_sc_hd__conb_1 _44253__483 (.HI(gpio_inp_dis[16]));
 sky130_fd_sc_hd__conb_1 _44254__484 (.HI(gpio_inp_dis[17]));
 sky130_fd_sc_hd__conb_1 _44255__485 (.HI(gpio_inp_dis[18]));
 sky130_fd_sc_hd__conb_1 _44256__486 (.HI(gpio_inp_dis[19]));
 sky130_fd_sc_hd__conb_1 _44257__487 (.HI(gpio_inp_dis[20]));
 sky130_fd_sc_hd__conb_1 _44258__488 (.HI(gpio_inp_dis[21]));
 sky130_fd_sc_hd__conb_1 _44259__489 (.HI(gpio_inp_dis[22]));
 sky130_fd_sc_hd__conb_1 _44260__490 (.HI(gpio_inp_dis[23]));
 sky130_fd_sc_hd__conb_1 _44261__491 (.HI(gpio_inp_dis[24]));
 sky130_fd_sc_hd__conb_1 _44266__492 (.HI(gpio_inp_dis[29]));
 sky130_fd_sc_hd__conb_1 _44267__493 (.HI(gpio_inp_dis[30]));
 sky130_fd_sc_hd__conb_1 _44268__494 (.HI(gpio_inp_dis[31]));
 sky130_fd_sc_hd__conb_1 _44269__495 (.HI(gpio_inp_dis[32]));
 sky130_fd_sc_hd__conb_1 _44270__496 (.HI(gpio_inp_dis[33]));
 sky130_fd_sc_hd__conb_1 _44271__497 (.HI(gpio_inp_dis[34]));
 sky130_fd_sc_hd__conb_1 _44272__498 (.HI(gpio_inp_dis[35]));
 sky130_fd_sc_hd__conb_1 _44273__499 (.HI(gpio_inp_dis[36]));
 sky130_fd_sc_hd__conb_1 _44274__500 (.HI(gpio_inp_dis[37]));
 sky130_fd_sc_hd__conb_1 _44276__501 (.HI(gpio_inp_dis[39]));
 sky130_fd_sc_hd__conb_1 _44278__502 (.HI(gpio_inp_dis[41]));
 sky130_fd_sc_hd__conb_1 _44279__503 (.HI(gpio_inp_dis[42]));
 sky130_fd_sc_hd__conb_1 _44280__504 (.HI(gpio_inp_dis[43]));
 sky130_fd_sc_hd__conb_1 _44288__505 (.HI(gpio_oeb[7]));
 sky130_fd_sc_hd__conb_1 _44297__506 (.HI(gpio_oeb[16]));
 sky130_fd_sc_hd__conb_1 _44298__507 (.HI(gpio_oeb[17]));
 sky130_fd_sc_hd__conb_1 _44299__508 (.HI(gpio_oeb[18]));
 sky130_fd_sc_hd__conb_1 _44300__509 (.HI(gpio_oeb[19]));
 sky130_fd_sc_hd__conb_1 _44301__510 (.HI(gpio_oeb[20]));
 sky130_fd_sc_hd__conb_1 _44302__511 (.HI(gpio_oeb[21]));
 sky130_fd_sc_hd__conb_1 _44303__512 (.HI(gpio_oeb[22]));
 sky130_fd_sc_hd__conb_1 _44304__513 (.HI(gpio_oeb[23]));
 sky130_fd_sc_hd__conb_1 _44305__514 (.HI(gpio_oeb[24]));
 sky130_fd_sc_hd__conb_1 _44310__515 (.HI(gpio_oeb[29]));
 sky130_fd_sc_hd__conb_1 _44311__516 (.HI(gpio_oeb[30]));
 sky130_fd_sc_hd__conb_1 _44312__517 (.HI(gpio_oeb[31]));
 sky130_fd_sc_hd__conb_1 _44313__518 (.HI(gpio_oeb[32]));
 sky130_fd_sc_hd__conb_1 _44314__519 (.HI(gpio_oeb[33]));
 sky130_fd_sc_hd__conb_1 _44315__520 (.HI(gpio_oeb[34]));
 sky130_fd_sc_hd__conb_1 _44316__521 (.HI(gpio_oeb[35]));
 sky130_fd_sc_hd__conb_1 _44317__522 (.HI(gpio_oeb[36]));
 sky130_fd_sc_hd__conb_1 _44318__523 (.HI(gpio_oeb[37]));
 sky130_fd_sc_hd__conb_1 _44319__524 (.HI(gpio_oeb[38]));
 sky130_fd_sc_hd__conb_1 _44320__525 (.HI(gpio_oeb[39]));
 sky130_fd_sc_hd__conb_1 _44321__526 (.HI(gpio_oeb[40]));
 sky130_fd_sc_hd__conb_1 _44322__527 (.HI(gpio_oeb[41]));
 sky130_fd_sc_hd__conb_1 _44323__528 (.HI(gpio_oeb[42]));
 sky130_fd_sc_hd__conb_1 _44324__529 (.HI(gpio_oeb[43]));
 sky130_fd_sc_hd__conb_1 \inst$top.soc.sram.mem.0.0_530  (.HI(net529));
 sky130_fd_sc_hd__conb_1 \inst$top.soc.sram.mem.0.0_531  (.HI(net530));
 sky130_fd_sc_hd__conb_1 \inst$top.soc.sram.mem.0.0_532  (.HI(net531));
 sky130_fd_sc_hd__buf_6 input533 (.A(gpio_in[10]),
    .X(net532));
 sky130_fd_sc_hd__buf_6 input534 (.A(gpio_in[11]),
    .X(net533));
 sky130_fd_sc_hd__buf_8 input535 (.A(gpio_in[12]),
    .X(net534));
 sky130_fd_sc_hd__buf_4 input536 (.A(gpio_in[13]),
    .X(net535));
 sky130_fd_sc_hd__buf_4 input537 (.A(gpio_in[14]),
    .X(net536));
 sky130_fd_sc_hd__buf_4 input538 (.A(gpio_in[15]),
    .X(net537));
 sky130_fd_sc_hd__buf_4 input539 (.A(gpio_in[25]),
    .X(net538));
 sky130_fd_sc_hd__buf_4 input540 (.A(gpio_in[26]),
    .X(net539));
 sky130_fd_sc_hd__buf_2 input541 (.A(gpio_in[27]),
    .X(net540));
 sky130_fd_sc_hd__buf_2 input542 (.A(gpio_in[28]),
    .X(net541));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input543 (.A(gpio_in[2]),
    .X(net542));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input544 (.A(gpio_in[3]),
    .X(net543));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input545 (.A(gpio_in[40]),
    .X(net544));
 sky130_fd_sc_hd__buf_4 input546 (.A(gpio_in[4]),
    .X(net545));
 sky130_fd_sc_hd__buf_4 input547 (.A(gpio_in[5]),
    .X(net546));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input548 (.A(net3034),
    .X(net547));
 sky130_fd_sc_hd__buf_6 input549 (.A(gpio_in[8]),
    .X(net548));
 sky130_fd_sc_hd__buf_6 input550 (.A(gpio_in[9]),
    .X(net549));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output551 (.A(net1622),
    .X(gpio_inp_dis[10]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output552 (.A(net1619),
    .X(gpio_inp_dis[11]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output553 (.A(net1615),
    .X(gpio_inp_dis[12]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output554 (.A(net1611),
    .X(gpio_inp_dis[13]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output555 (.A(net1606),
    .X(gpio_inp_dis[14]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output556 (.A(net1602),
    .X(gpio_inp_dis[15]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output557 (.A(net1632),
    .X(gpio_inp_dis[25]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output558 (.A(net1631),
    .X(gpio_inp_dis[26]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output559 (.A(net1610),
    .X(gpio_inp_dis[27]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output560 (.A(net1601),
    .X(gpio_inp_dis[28]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output561 (.A(net2575),
    .X(gpio_inp_dis[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output562 (.A(net2573),
    .X(gpio_inp_dis[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output563 (.A(net2571),
    .X(gpio_inp_dis[4]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output564 (.A(net2569),
    .X(gpio_inp_dis[5]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output565 (.A(net1628),
    .X(gpio_inp_dis[8]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output566 (.A(net1625),
    .X(gpio_inp_dis[9]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output567 (.A(net566),
    .X(gpio_oeb[10]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output568 (.A(net567),
    .X(gpio_oeb[11]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output569 (.A(net568),
    .X(gpio_oeb[12]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output570 (.A(net569),
    .X(gpio_oeb[13]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output571 (.A(net570),
    .X(gpio_oeb[14]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output572 (.A(net571),
    .X(gpio_oeb[15]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output573 (.A(net572),
    .X(gpio_oeb[25]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output574 (.A(net573),
    .X(gpio_oeb[26]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output575 (.A(net574),
    .X(gpio_oeb[27]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output576 (.A(net575),
    .X(gpio_oeb[28]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output577 (.A(net576),
    .X(gpio_oeb[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output578 (.A(net577),
    .X(gpio_oeb[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output579 (.A(net578),
    .X(gpio_oeb[4]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output580 (.A(net579),
    .X(gpio_oeb[5]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output581 (.A(net580),
    .X(gpio_oeb[8]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output582 (.A(net581),
    .X(gpio_oeb[9]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output583 (.A(net2568),
    .X(gpio_out[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output584 (.A(net1750),
    .X(gpio_out[10]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output585 (.A(net1747),
    .X(gpio_out[11]));
 sky130_fd_sc_hd__buf_6 output586 (.A(net1746),
    .X(gpio_out[12]));
 sky130_fd_sc_hd__buf_8 output587 (.A(net586),
    .X(gpio_out[13]));
 sky130_fd_sc_hd__buf_8 output588 (.A(net587),
    .X(gpio_out[14]));
 sky130_fd_sc_hd__buf_4 output589 (.A(net1745),
    .X(gpio_out[15]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output590 (.A(net589),
    .X(gpio_out[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output591 (.A(net1744),
    .X(gpio_out[25]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output592 (.A(net1743),
    .X(gpio_out[26]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output593 (.A(net1742),
    .X(gpio_out[27]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output594 (.A(net1741),
    .X(gpio_out[28]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output595 (.A(net2576),
    .X(gpio_out[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output596 (.A(net2574),
    .X(gpio_out[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output597 (.A(net2572),
    .X(gpio_out[4]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output598 (.A(net2570),
    .X(gpio_out[5]));
 sky130_fd_sc_hd__buf_4 output599 (.A(net598),
    .X(gpio_out[6]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output600 (.A(net1756),
    .X(gpio_out[8]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output601 (.A(net1753),
    .X(gpio_out[9]));
 sky130_fd_sc_hd__buf_6 wire602 (.A(_15152_),
    .X(net601));
 sky130_fd_sc_hd__buf_6 wire603 (.A(_13295_),
    .X(net602));
 sky130_fd_sc_hd__buf_6 wire604 (.A(_13858_),
    .X(net603));
 sky130_fd_sc_hd__buf_6 wire605 (.A(_13338_),
    .X(net604));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout606 (.A(net608),
    .X(net605));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout607 (.A(net607),
    .X(net606));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout608 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout609 (.A(_10303_),
    .X(net608));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout610 (.A(_10024_),
    .X(net609));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout611 (.A(_10024_),
    .X(net610));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout612 (.A(net613),
    .X(net611));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout613 (.A(net613),
    .X(net612));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout614 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout615 (.A(_09841_),
    .X(net614));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout616 (.A(net618),
    .X(net615));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout617 (.A(net617),
    .X(net616));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout618 (.A(net618),
    .X(net617));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout619 (.A(net619),
    .X(net618));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout620 (.A(_09841_),
    .X(net619));
 sky130_fd_sc_hd__buf_4 wire621 (.A(_14492_),
    .X(net620));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout622 (.A(net632),
    .X(net621));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout623 (.A(net632),
    .X(net622));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout624 (.A(net625),
    .X(net623));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout625 (.A(net625),
    .X(net624));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout626 (.A(net632),
    .X(net625));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout627 (.A(net631),
    .X(net626));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout628 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout629 (.A(net631),
    .X(net628));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout630 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout631 (.A(net631),
    .X(net630));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout632 (.A(net632),
    .X(net631));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout633 (.A(net634),
    .X(net632));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout634 (.A(net634),
    .X(net633));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout635 (.A(net661),
    .X(net634));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout636 (.A(net636),
    .X(net635));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout637 (.A(net637),
    .X(net636));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout638 (.A(net646),
    .X(net637));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout639 (.A(net640),
    .X(net638));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout640 (.A(net640),
    .X(net639));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout641 (.A(net646),
    .X(net640));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout642 (.A(net642),
    .X(net641));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout643 (.A(net643),
    .X(net642));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout644 (.A(net646),
    .X(net643));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout645 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout646 (.A(net646),
    .X(net645));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout647 (.A(net661),
    .X(net646));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout648 (.A(net648),
    .X(net647));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout649 (.A(net649),
    .X(net648));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout650 (.A(net652),
    .X(net649));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout651 (.A(net652),
    .X(net650));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout652 (.A(net652),
    .X(net651));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout653 (.A(net661),
    .X(net652));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout654 (.A(net655),
    .X(net653));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout655 (.A(net655),
    .X(net654));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout656 (.A(net661),
    .X(net655));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout657 (.A(net660),
    .X(net656));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout658 (.A(net660),
    .X(net657));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout659 (.A(net659),
    .X(net658));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout660 (.A(net660),
    .X(net659));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout661 (.A(net661),
    .X(net660));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout662 (.A(_09415_),
    .X(net661));
 sky130_fd_sc_hd__buf_16 wire663 (.A(_14550_),
    .X(net662));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout664 (.A(net664),
    .X(net663));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout665 (.A(net665),
    .X(net664));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout666 (.A(_09413_),
    .X(net665));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout667 (.A(net674),
    .X(net666));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout668 (.A(net674),
    .X(net667));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout669 (.A(net670),
    .X(net668));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout670 (.A(net670),
    .X(net669));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout671 (.A(net674),
    .X(net670));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout672 (.A(net673),
    .X(net671));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout673 (.A(net673),
    .X(net672));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout674 (.A(net674),
    .X(net673));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout675 (.A(net721),
    .X(net674));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout676 (.A(net676),
    .X(net675));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout677 (.A(net678),
    .X(net676));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout678 (.A(net678),
    .X(net677));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout679 (.A(net681),
    .X(net678));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout680 (.A(net680),
    .X(net679));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout681 (.A(net681),
    .X(net680));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout682 (.A(net721),
    .X(net681));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout683 (.A(net685),
    .X(net682));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout684 (.A(net684),
    .X(net683));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout685 (.A(net685),
    .X(net684));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout686 (.A(net703),
    .X(net685));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout687 (.A(net689),
    .X(net686));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout688 (.A(net689),
    .X(net687));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout689 (.A(net689),
    .X(net688));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout690 (.A(net703),
    .X(net689));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout691 (.A(net691),
    .X(net690));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout692 (.A(net692),
    .X(net691));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout693 (.A(net703),
    .X(net692));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout694 (.A(net694),
    .X(net693));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout695 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout696 (.A(net698),
    .X(net695));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout697 (.A(net697),
    .X(net696));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout698 (.A(net698),
    .X(net697));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout699 (.A(net703),
    .X(net698));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout700 (.A(net703),
    .X(net699));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout701 (.A(net702),
    .X(net700));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout702 (.A(net702),
    .X(net701));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout703 (.A(net703),
    .X(net702));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout704 (.A(net721),
    .X(net703));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout705 (.A(net705),
    .X(net704));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout706 (.A(net708),
    .X(net705));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout707 (.A(net708),
    .X(net706));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout708 (.A(net708),
    .X(net707));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout709 (.A(net711),
    .X(net708));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout710 (.A(net710),
    .X(net709));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout711 (.A(net711),
    .X(net710));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout712 (.A(net722),
    .X(net711));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout713 (.A(net713),
    .X(net712));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout714 (.A(net714),
    .X(net713));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout715 (.A(net722),
    .X(net714));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout716 (.A(net716),
    .X(net715));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout717 (.A(net722),
    .X(net716));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout718 (.A(net720),
    .X(net717));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout719 (.A(net720),
    .X(net718));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout720 (.A(net720),
    .X(net719));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout721 (.A(net722),
    .X(net720));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout722 (.A(_20370_),
    .X(net721));
 sky130_fd_sc_hd__buf_12 wire723 (.A(net721),
    .X(net722));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout724 (.A(_10023_),
    .X(net723));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout725 (.A(_10023_),
    .X(net724));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout726 (.A(_10023_),
    .X(net725));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout727 (.A(_10023_),
    .X(net726));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout728 (.A(net728),
    .X(net727));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout729 (.A(_14814_),
    .X(net728));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout730 (.A(_14600_),
    .X(net729));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout731 (.A(_14589_),
    .X(net730));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout732 (.A(_14587_),
    .X(net731));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout733 (.A(_14584_),
    .X(net732));
 sky130_fd_sc_hd__buf_4 load_slew734 (.A(_14584_),
    .X(net733));
 sky130_fd_sc_hd__buf_16 wire735 (.A(_14519_),
    .X(net734));
 sky130_fd_sc_hd__buf_8 wire736 (.A(_14464_),
    .X(net735));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout737 (.A(_12960_),
    .X(net736));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout738 (.A(net738),
    .X(net737));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout739 (.A(net739),
    .X(net738));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout740 (.A(_12957_),
    .X(net739));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout741 (.A(_11915_),
    .X(net740));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout742 (.A(_11915_),
    .X(net741));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout743 (.A(_11915_),
    .X(net742));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout744 (.A(_11915_),
    .X(net743));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout745 (.A(net746),
    .X(net744));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout746 (.A(net746),
    .X(net745));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout747 (.A(net752),
    .X(net746));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout748 (.A(net748),
    .X(net747));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout749 (.A(net752),
    .X(net748));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout750 (.A(net752),
    .X(net749));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout751 (.A(net752),
    .X(net750));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout752 (.A(net752),
    .X(net751));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout753 (.A(_09927_),
    .X(net752));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout754 (.A(net754),
    .X(net753));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout755 (.A(net755),
    .X(net754));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout756 (.A(_09414_),
    .X(net755));
 sky130_fd_sc_hd__buf_12 wire757 (.A(net757),
    .X(net756));
 sky130_fd_sc_hd__buf_12 wire758 (.A(\inst$top.soc.sram.write_port__en[2] ),
    .X(net757));
 sky130_fd_sc_hd__buf_12 wire759 (.A(net759),
    .X(net758));
 sky130_fd_sc_hd__buf_12 wire760 (.A(\inst$top.soc.sram.write_port__en[3] ),
    .X(net759));
 sky130_fd_sc_hd__buf_16 wire761 (.A(\inst$top.soc.sram.write_port__en[0] ),
    .X(net760));
 sky130_fd_sc_hd__buf_12 load_slew762 (.A(net762),
    .X(net761));
 sky130_fd_sc_hd__buf_12 wire763 (.A(\inst$top.soc.sram.write_port__en[1] ),
    .X(net762));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout764 (.A(net764),
    .X(net763));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout765 (.A(net778),
    .X(net764));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout766 (.A(net766),
    .X(net765));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout767 (.A(net778),
    .X(net766));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout768 (.A(net778),
    .X(net767));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout769 (.A(net778),
    .X(net768));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout770 (.A(net770),
    .X(net769));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout771 (.A(net778),
    .X(net770));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout772 (.A(net776),
    .X(net771));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout773 (.A(net776),
    .X(net772));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout774 (.A(net775),
    .X(net773));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout775 (.A(net775),
    .X(net774));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout776 (.A(net776),
    .X(net775));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout777 (.A(net778),
    .X(net776));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout778 (.A(net778),
    .X(net777));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout779 (.A(_14813_),
    .X(net778));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout780 (.A(net780),
    .X(net779));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout781 (.A(_14588_),
    .X(net780));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout782 (.A(_14586_),
    .X(net781));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout783 (.A(_14586_),
    .X(net782));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout784 (.A(net784),
    .X(net783));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout785 (.A(net785),
    .X(net784));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout786 (.A(_12983_),
    .X(net785));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout787 (.A(net787),
    .X(net786));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout788 (.A(_12959_),
    .X(net787));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout789 (.A(_02205_),
    .X(net788));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout790 (.A(_02178_),
    .X(net789));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout791 (.A(_20363_),
    .X(net790));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout792 (.A(_20363_),
    .X(net791));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout793 (.A(_20363_),
    .X(net792));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout794 (.A(_20363_),
    .X(net793));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout795 (.A(net795),
    .X(net794));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout796 (.A(_19652_),
    .X(net795));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout797 (.A(net798),
    .X(net796));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout798 (.A(net798),
    .X(net797));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout799 (.A(_19591_),
    .X(net798));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout800 (.A(_19591_),
    .X(net799));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout801 (.A(_19529_),
    .X(net800));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout802 (.A(_19529_),
    .X(net801));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout803 (.A(_19505_),
    .X(net802));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout804 (.A(_19505_),
    .X(net803));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout805 (.A(_19439_),
    .X(net804));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout806 (.A(_19439_),
    .X(net805));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout807 (.A(_18628_),
    .X(net806));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout808 (.A(_18179_),
    .X(net807));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout809 (.A(_18147_),
    .X(net808));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout810 (.A(_18147_),
    .X(net809));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout811 (.A(_14919_),
    .X(net810));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout812 (.A(_14919_),
    .X(net811));
 sky130_fd_sc_hd__buf_16 wire813 (.A(_14402_),
    .X(net812));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout814 (.A(net815),
    .X(net813));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout815 (.A(net815),
    .X(net814));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout816 (.A(_11907_),
    .X(net815));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout817 (.A(_11907_),
    .X(net816));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout818 (.A(_11907_),
    .X(net817));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout819 (.A(net820),
    .X(net818));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout820 (.A(net820),
    .X(net819));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout821 (.A(_01725_),
    .X(net820));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout822 (.A(_19641_),
    .X(net821));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout823 (.A(_19641_),
    .X(net822));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout824 (.A(_19630_),
    .X(net823));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout825 (.A(_19630_),
    .X(net824));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout826 (.A(net826),
    .X(net825));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout827 (.A(_19518_),
    .X(net826));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout828 (.A(_18741_),
    .X(net827));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout829 (.A(_18535_),
    .X(net828));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout830 (.A(_18048_),
    .X(net829));
 sky130_fd_sc_hd__buf_16 wire831 (.A(_14370_),
    .X(net830));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout832 (.A(net834),
    .X(net831));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout833 (.A(net834),
    .X(net832));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout834 (.A(net834),
    .X(net833));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout835 (.A(_11914_),
    .X(net834));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout836 (.A(_10307_),
    .X(net835));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout837 (.A(_10307_),
    .X(net836));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout838 (.A(net838),
    .X(net837));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout839 (.A(_20362_),
    .X(net838));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout840 (.A(net840),
    .X(net839));
 sky130_fd_sc_hd__buf_4 wire841 (.A(_18082_),
    .X(net840));
 sky130_fd_sc_hd__buf_4 wire842 (.A(_18073_),
    .X(net841));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout843 (.A(_17987_),
    .X(net842));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout844 (.A(_17987_),
    .X(net843));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout845 (.A(net845),
    .X(net844));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout846 (.A(_17933_),
    .X(net845));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout847 (.A(net848),
    .X(net846));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout848 (.A(net848),
    .X(net847));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout849 (.A(_11930_),
    .X(net848));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout850 (.A(net850),
    .X(net849));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout851 (.A(net851),
    .X(net850));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout852 (.A(_11930_),
    .X(net851));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout853 (.A(_10318_),
    .X(net852));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout854 (.A(_10318_),
    .X(net853));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout855 (.A(_09992_),
    .X(net854));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout856 (.A(_09992_),
    .X(net855));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout857 (.A(_09992_),
    .X(net856));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout858 (.A(_09992_),
    .X(net857));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout859 (.A(net859),
    .X(net858));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout860 (.A(net862),
    .X(net859));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout861 (.A(net862),
    .X(net860));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout862 (.A(net862),
    .X(net861));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout863 (.A(_09336_),
    .X(net862));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout864 (.A(_19670_),
    .X(net863));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout865 (.A(_19178_),
    .X(net864));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout866 (.A(_18483_),
    .X(net865));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout867 (.A(_18480_),
    .X(net866));
 sky130_fd_sc_hd__buf_12 load_slew868 (.A(_17967_),
    .X(net867));
 sky130_fd_sc_hd__buf_12 load_slew869 (.A(_17948_),
    .X(net868));
 sky130_fd_sc_hd__buf_16 wire870 (.A(_14252_),
    .X(net869));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout871 (.A(_11929_),
    .X(net870));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout872 (.A(_11929_),
    .X(net871));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout873 (.A(net875),
    .X(net872));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout874 (.A(net874),
    .X(net873));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout875 (.A(net875),
    .X(net874));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout876 (.A(net880),
    .X(net875));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout877 (.A(net880),
    .X(net876));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout878 (.A(net878),
    .X(net877));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout879 (.A(net879),
    .X(net878));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout880 (.A(net880),
    .X(net879));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout881 (.A(_20255_),
    .X(net880));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout882 (.A(_19170_),
    .X(net881));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout883 (.A(_18403_),
    .X(net882));
 sky130_fd_sc_hd__buf_4 wire884 (.A(_11912_),
    .X(net883));
 sky130_fd_sc_hd__buf_8 wire885 (.A(_06042_),
    .X(net884));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout886 (.A(net886),
    .X(net885));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout887 (.A(net889),
    .X(net886));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout888 (.A(net888),
    .X(net887));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout889 (.A(net889),
    .X(net888));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout890 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[15] ),
    .X(net889));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout891 (.A(net891),
    .X(net890));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout892 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[7] ),
    .X(net891));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout893 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout894 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[7] ),
    .X(net893));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout895 (.A(_19694_),
    .X(net894));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout896 (.A(_19694_),
    .X(net895));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout897 (.A(net897),
    .X(net896));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout898 (.A(_19674_),
    .X(net897));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout899 (.A(_19672_),
    .X(net898));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout900 (.A(_19672_),
    .X(net899));
 sky130_fd_sc_hd__buf_12 load_slew901 (.A(_17941_),
    .X(net900));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout902 (.A(net904),
    .X(net901));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout903 (.A(net903),
    .X(net902));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout904 (.A(net904),
    .X(net903));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout905 (.A(net905),
    .X(net904));
 sky130_fd_sc_hd__buf_2 fanout906 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[31] ),
    .X(net905));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout907 (.A(net909),
    .X(net906));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout908 (.A(net909),
    .X(net907));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout909 (.A(net909),
    .X(net908));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout910 (.A(net910),
    .X(net909));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout911 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[30] ),
    .X(net910));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout912 (.A(net914),
    .X(net911));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout913 (.A(net914),
    .X(net912));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout914 (.A(net914),
    .X(net913));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout915 (.A(net915),
    .X(net914));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout916 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[29] ),
    .X(net915));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout917 (.A(net919),
    .X(net916));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout918 (.A(net918),
    .X(net917));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout919 (.A(net919),
    .X(net918));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout920 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[28] ),
    .X(net919));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout921 (.A(net923),
    .X(net920));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout922 (.A(net922),
    .X(net921));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout923 (.A(net923),
    .X(net922));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout924 (.A(net924),
    .X(net923));
 sky130_fd_sc_hd__buf_2 fanout925 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[27] ),
    .X(net924));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout926 (.A(net928),
    .X(net925));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout927 (.A(net928),
    .X(net926));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout928 (.A(net928),
    .X(net927));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout929 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[26] ),
    .X(net928));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout930 (.A(net933),
    .X(net929));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout931 (.A(net932),
    .X(net930));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout932 (.A(net932),
    .X(net931));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout933 (.A(net933),
    .X(net932));
 sky130_fd_sc_hd__buf_2 fanout934 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[25] ),
    .X(net933));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout935 (.A(net935),
    .X(net934));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout936 (.A(net938),
    .X(net935));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout937 (.A(net937),
    .X(net936));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout938 (.A(net938),
    .X(net937));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout939 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[24] ),
    .X(net938));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout940 (.A(net941),
    .X(net939));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout941 (.A(net941),
    .X(net940));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout942 (.A(net942),
    .X(net941));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout943 (.A(net943),
    .X(net942));
 sky130_fd_sc_hd__buf_4 load_slew944 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[23] ),
    .X(net943));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout945 (.A(net947),
    .X(net944));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout946 (.A(net947),
    .X(net945));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout947 (.A(net947),
    .X(net946));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout948 (.A(net948),
    .X(net947));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout949 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[22] ),
    .X(net948));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout950 (.A(net951),
    .X(net949));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout951 (.A(net951),
    .X(net950));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout952 (.A(net952),
    .X(net951));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout953 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[21] ),
    .X(net952));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout954 (.A(net955),
    .X(net953));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout955 (.A(net955),
    .X(net954));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout956 (.A(net956),
    .X(net955));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout957 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__buf_4 load_slew958 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[20] ),
    .X(net957));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout959 (.A(net960),
    .X(net958));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout960 (.A(net960),
    .X(net959));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout961 (.A(net961),
    .X(net960));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout962 (.A(net962),
    .X(net961));
 sky130_fd_sc_hd__buf_8 load_slew963 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[19] ),
    .X(net962));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout964 (.A(net966),
    .X(net963));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout965 (.A(net966),
    .X(net964));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout966 (.A(net966),
    .X(net965));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout967 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[18] ),
    .X(net966));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout968 (.A(net969),
    .X(net967));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout969 (.A(net970),
    .X(net968));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout970 (.A(net970),
    .X(net969));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout971 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[17] ),
    .X(net970));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout972 (.A(net974),
    .X(net971));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout973 (.A(net973),
    .X(net972));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout974 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout975 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[16] ),
    .X(net974));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout976 (.A(net977),
    .X(net975));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout977 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout978 (.A(net978),
    .X(net977));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout979 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__buf_8 wire980 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[14] ),
    .X(net979));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout981 (.A(net982),
    .X(net980));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout982 (.A(net982),
    .X(net981));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout983 (.A(net983),
    .X(net982));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout984 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[13] ),
    .X(net983));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout985 (.A(net987),
    .X(net984));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout986 (.A(net986),
    .X(net985));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout987 (.A(net987),
    .X(net986));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout988 (.A(net988),
    .X(net987));
 sky130_fd_sc_hd__buf_8 wire989 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[12] ),
    .X(net988));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout990 (.A(net991),
    .X(net989));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout991 (.A(net991),
    .X(net990));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout992 (.A(net992),
    .X(net991));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout993 (.A(net993),
    .X(net992));
 sky130_fd_sc_hd__buf_4 wire994 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[11] ),
    .X(net993));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout995 (.A(net997),
    .X(net994));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout996 (.A(net996),
    .X(net995));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout997 (.A(net997),
    .X(net996));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout998 (.A(net998),
    .X(net997));
 sky130_fd_sc_hd__buf_6 wire999 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[10] ),
    .X(net998));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1000 (.A(net1002),
    .X(net999));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1001 (.A(net1002),
    .X(net1000));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1002 (.A(net1002),
    .X(net1001));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1003 (.A(net1003),
    .X(net1002));
 sky130_fd_sc_hd__buf_4 wire1004 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[9] ),
    .X(net1003));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1005 (.A(net1006),
    .X(net1004));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1006 (.A(net1006),
    .X(net1005));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1007 (.A(net1007),
    .X(net1006));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1008 (.A(net1008),
    .X(net1007));
 sky130_fd_sc_hd__buf_4 wire1009 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[8] ),
    .X(net1008));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1010 (.A(net1013),
    .X(net1009));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1011 (.A(net1012),
    .X(net1010));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1012 (.A(net1012),
    .X(net1011));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1013 (.A(net1013),
    .X(net1012));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1014 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[4] ),
    .X(net1013));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1015 (.A(net1017),
    .X(net1014));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1016 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1017 (.A(net1017),
    .X(net1016));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1018 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[1] ),
    .X(net1017));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1019 (.A(_20226_),
    .X(net1018));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1020 (.A(_20226_),
    .X(net1019));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1021 (.A(net1021),
    .X(net1020));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1022 (.A(_20226_),
    .X(net1021));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1023 (.A(_18460_),
    .X(net1022));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1024 (.A(_18460_),
    .X(net1023));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1025 (.A(_14881_),
    .X(net1024));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1026 (.A(_12721_),
    .X(net1025));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1027 (.A(_12721_),
    .X(net1026));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1028 (.A(net1030),
    .X(net1027));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1029 (.A(net1029),
    .X(net1028));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1030 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1031 (.A(_11722_),
    .X(net1030));
 sky130_fd_sc_hd__buf_6 wire1032 (.A(_11016_),
    .X(net1031));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1033 (.A(net1034),
    .X(net1032));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1034 (.A(net1034),
    .X(net1033));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1035 (.A(net1035),
    .X(net1034));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1036 (.A(_09993_),
    .X(net1035));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1037 (.A(net1040),
    .X(net1036));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1038 (.A(net1040),
    .X(net1037));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1039 (.A(net1040),
    .X(net1038));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1040 (.A(net1040),
    .X(net1039));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1041 (.A(_09993_),
    .X(net1040));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1042 (.A(net1042),
    .X(net1041));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1043 (.A(_09450_),
    .X(net1042));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1044 (.A(net1044),
    .X(net1043));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1045 (.A(_09450_),
    .X(net1044));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1046 (.A(net1047),
    .X(net1045));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1047 (.A(net1047),
    .X(net1046));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1048 (.A(_06014_),
    .X(net1047));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1049 (.A(net1050),
    .X(net1048));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1050 (.A(net1050),
    .X(net1049));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1051 (.A(net1051),
    .X(net1050));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1052 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[6] ),
    .X(net1051));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1053 (.A(net1053),
    .X(net1052));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1054 (.A(net1055),
    .X(net1053));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1055 (.A(net1055),
    .X(net1054));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1056 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[5] ),
    .X(net1055));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1057 (.A(net1058),
    .X(net1056));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1058 (.A(net1058),
    .X(net1057));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1059 (.A(net1059),
    .X(net1058));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1060 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[3] ),
    .X(net1059));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1061 (.A(net1061),
    .X(net1060));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1062 (.A(net1062),
    .X(net1061));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1063 (.A(net1063),
    .X(net1062));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1064 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[2] ),
    .X(net1063));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1065 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[0] ),
    .X(net1064));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1066 (.A(net1067),
    .X(net1065));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1067 (.A(net1067),
    .X(net1066));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1068 (.A(\inst$top.soc.cpu.gprf.bypass1.w_wp_data[0] ),
    .X(net1067));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1069 (.A(_20195_),
    .X(net1068));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1070 (.A(_20195_),
    .X(net1069));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1071 (.A(net1071),
    .X(net1070));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1072 (.A(_20195_),
    .X(net1071));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1073 (.A(net1074),
    .X(net1072));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1074 (.A(net1074),
    .X(net1073));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1075 (.A(net1075),
    .X(net1074));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1076 (.A(net1076),
    .X(net1075));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1077 (.A(net1077),
    .X(net1076));
 sky130_fd_sc_hd__buf_2 fanout1078 (.A(_20100_),
    .X(net1077));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1079 (.A(net1081),
    .X(net1078));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1080 (.A(net1081),
    .X(net1079));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1081 (.A(net1081),
    .X(net1080));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1082 (.A(_19103_),
    .X(net1081));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1083 (.A(_12707_),
    .X(net1082));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1084 (.A(_12707_),
    .X(net1083));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1085 (.A(net1087),
    .X(net1084));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1086 (.A(net1087),
    .X(net1085));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1087 (.A(net1087),
    .X(net1086));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1088 (.A(_12703_),
    .X(net1087));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1089 (.A(net1091),
    .X(net1088));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1090 (.A(net1090),
    .X(net1089));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1091 (.A(net1091),
    .X(net1090));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1092 (.A(_11399_),
    .X(net1091));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1093 (.A(net1095),
    .X(net1092));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1094 (.A(net1094),
    .X(net1093));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1095 (.A(net1095),
    .X(net1094));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1096 (.A(_11030_),
    .X(net1095));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1097 (.A(net1099),
    .X(net1096));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1098 (.A(net1098),
    .X(net1097));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1099 (.A(net1099),
    .X(net1098));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1100 (.A(_10915_),
    .X(net1099));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1101 (.A(net1103),
    .X(net1100));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1102 (.A(net1102),
    .X(net1101));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1103 (.A(net1103),
    .X(net1102));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1104 (.A(_09923_),
    .X(net1103));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1105 (.A(net1105),
    .X(net1104));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1106 (.A(_09909_),
    .X(net1105));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1107 (.A(net1107),
    .X(net1106));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1108 (.A(_06011_),
    .X(net1107));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1109 (.A(net1109),
    .X(net1108));
 sky130_fd_sc_hd__buf_16 wire1110 (.A(_06011_),
    .X(net1109));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1111 (.A(net1113),
    .X(net1110));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1112 (.A(net1113),
    .X(net1111));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1113 (.A(net1113),
    .X(net1112));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1114 (.A(_06002_),
    .X(net1113));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1115 (.A(net1116),
    .X(net1114));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1116 (.A(net1116),
    .X(net1115));
 sky130_fd_sc_hd__buf_2 fanout1117 (.A(_05997_),
    .X(net1116));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1118 (.A(net1119),
    .X(net1117));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1119 (.A(_05987_),
    .X(net1118));
 sky130_fd_sc_hd__buf_16 load_slew1120 (.A(net1118),
    .X(net1119));
 sky130_fd_sc_hd__buf_12 wire1121 (.A(_05987_),
    .X(net1120));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1122 (.A(net1122),
    .X(net1121));
 sky130_fd_sc_hd__buf_2 fanout1123 (.A(_05968_),
    .X(net1122));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1124 (.A(net1125),
    .X(net1123));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1125 (.A(_05962_),
    .X(net1124));
 sky130_fd_sc_hd__buf_16 max_cap1126 (.A(net1124),
    .X(net1125));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1127 (.A(net1128),
    .X(net1126));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1128 (.A(_05950_),
    .X(net1127));
 sky130_fd_sc_hd__buf_16 wire1129 (.A(net1127),
    .X(net1128));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1130 (.A(net1131),
    .X(net1129));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1131 (.A(_05948_),
    .X(net1130));
 sky130_fd_sc_hd__buf_16 wire1132 (.A(net1130),
    .X(net1131));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1133 (.A(net1133),
    .X(net1132));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1134 (.A(net1134),
    .X(net1133));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1135 (.A(net1135),
    .X(net1134));
 sky130_fd_sc_hd__buf_2 fanout1136 (.A(_05947_),
    .X(net1135));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1137 (.A(_05945_),
    .X(net1136));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1138 (.A(_05940_),
    .X(net1137));
 sky130_fd_sc_hd__buf_16 wire1139 (.A(net1137),
    .X(net1138));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1140 (.A(_05938_),
    .X(net1139));
 sky130_fd_sc_hd__buf_16 load_slew1141 (.A(net1139),
    .X(net1140));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1142 (.A(_05935_),
    .X(net1141));
 sky130_fd_sc_hd__buf_16 load_slew1143 (.A(net1141),
    .X(net1142));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1144 (.A(_05931_),
    .X(net1143));
 sky130_fd_sc_hd__buf_16 wire1145 (.A(net1143),
    .X(net1144));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1146 (.A(_05928_),
    .X(net1145));
 sky130_fd_sc_hd__buf_16 load_slew1147 (.A(net1145),
    .X(net1146));
 sky130_fd_sc_hd__buf_12 wire1148 (.A(_05928_),
    .X(net1147));
 sky130_fd_sc_hd__buf_2 fanout1149 (.A(_05920_),
    .X(net1148));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1150 (.A(_05920_),
    .X(net1149));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1151 (.A(_05916_),
    .X(net1150));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1152 (.A(_05916_),
    .X(net1151));
 sky130_fd_sc_hd__buf_2 fanout1153 (.A(_05912_),
    .X(net1152));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1154 (.A(net1155),
    .X(net1153));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1155 (.A(net1155),
    .X(net1154));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1156 (.A(_05910_),
    .X(net1155));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1157 (.A(_05908_),
    .X(net1156));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1158 (.A(_05903_),
    .X(net1157));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1159 (.A(_05901_),
    .X(net1158));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1160 (.A(_05897_),
    .X(net1159));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1161 (.A(net1162),
    .X(net1160));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1162 (.A(_20683_),
    .X(net1161));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1163 (.A(_20683_),
    .X(net1162));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1164 (.A(_20630_),
    .X(net1163));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1165 (.A(net1165),
    .X(net1164));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1166 (.A(_20630_),
    .X(net1165));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1167 (.A(net1169),
    .X(net1166));
 sky130_fd_sc_hd__buf_2 fanout1168 (.A(net1169),
    .X(net1167));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1169 (.A(net1169),
    .X(net1168));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1170 (.A(_20601_),
    .X(net1169));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1171 (.A(net1172),
    .X(net1170));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1172 (.A(_20572_),
    .X(net1171));
 sky130_fd_sc_hd__buf_12 wire1173 (.A(net1171),
    .X(net1172));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1174 (.A(net1174),
    .X(net1173));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1175 (.A(_20506_),
    .X(net1174));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1176 (.A(net1177),
    .X(net1175));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1177 (.A(net1177),
    .X(net1176));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1178 (.A(net1180),
    .X(net1177));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1179 (.A(net1179),
    .X(net1178));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1180 (.A(net1180),
    .X(net1179));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1181 (.A(_20506_),
    .X(net1180));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1182 (.A(net1182),
    .X(net1181));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1183 (.A(net1183),
    .X(net1182));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1184 (.A(_20465_),
    .X(net1183));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1185 (.A(net1185),
    .X(net1184));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1186 (.A(net1189),
    .X(net1185));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1187 (.A(net1187),
    .X(net1186));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1188 (.A(net1188),
    .X(net1187));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1189 (.A(net1189),
    .X(net1188));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1190 (.A(net1190),
    .X(net1189));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1191 (.A(_20465_),
    .X(net1190));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1192 (.A(_20349_),
    .X(net1191));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1193 (.A(net1195),
    .X(net1192));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1194 (.A(net1194),
    .X(net1193));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1195 (.A(net1195),
    .X(net1194));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1196 (.A(_20220_),
    .X(net1195));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1197 (.A(net1197),
    .X(net1196));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1198 (.A(net1202),
    .X(net1197));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1199 (.A(net1199),
    .X(net1198));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1200 (.A(net1201),
    .X(net1199));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1201 (.A(net1201),
    .X(net1200));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1202 (.A(net1202),
    .X(net1201));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1203 (.A(_20099_),
    .X(net1202));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1204 (.A(_20062_),
    .X(net1203));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1205 (.A(net1205),
    .X(net1204));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1206 (.A(net1206),
    .X(net1205));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1207 (.A(_20062_),
    .X(net1206));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1208 (.A(net1209),
    .X(net1207));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1209 (.A(net1209),
    .X(net1208));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1210 (.A(net1210),
    .X(net1209));
 sky130_fd_sc_hd__buf_2 fanout1211 (.A(_19998_),
    .X(net1210));
 sky130_fd_sc_hd__buf_2 fanout1212 (.A(_19992_),
    .X(net1211));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1213 (.A(_19984_),
    .X(net1212));
 sky130_fd_sc_hd__buf_16 max_cap1214 (.A(net1212),
    .X(net1213));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1215 (.A(net1216),
    .X(net1214));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1216 (.A(net1216),
    .X(net1215));
 sky130_fd_sc_hd__buf_2 fanout1217 (.A(_19974_),
    .X(net1216));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1218 (.A(_19946_),
    .X(net1217));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1219 (.A(_19932_),
    .X(net1218));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1220 (.A(_19919_),
    .X(net1219));
 sky130_fd_sc_hd__buf_12 wire1221 (.A(net1219),
    .X(net1220));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1222 (.A(net1223),
    .X(net1221));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1223 (.A(_19884_),
    .X(net1222));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1224 (.A(_19884_),
    .X(net1223));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1225 (.A(_18856_),
    .X(net1224));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1226 (.A(_18856_),
    .X(net1225));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1227 (.A(_18809_),
    .X(net1226));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1228 (.A(net1228),
    .X(net1227));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1229 (.A(_14887_),
    .X(net1228));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1230 (.A(net1230),
    .X(net1229));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1231 (.A(_12976_),
    .X(net1230));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1232 (.A(_12976_),
    .X(net1231));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1233 (.A(_12976_),
    .X(net1232));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1234 (.A(net1236),
    .X(net1233));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1235 (.A(net1235),
    .X(net1234));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1236 (.A(net1236),
    .X(net1235));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1237 (.A(_11402_),
    .X(net1236));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1238 (.A(net1240),
    .X(net1237));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1239 (.A(net1239),
    .X(net1238));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1240 (.A(net1240),
    .X(net1239));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1241 (.A(_11033_),
    .X(net1240));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1242 (.A(net1244),
    .X(net1241));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1243 (.A(net1243),
    .X(net1242));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1244 (.A(net1244),
    .X(net1243));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1245 (.A(_10918_),
    .X(net1244));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1246 (.A(_09907_),
    .X(net1245));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1247 (.A(net1247),
    .X(net1246));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1248 (.A(_09648_),
    .X(net1247));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1249 (.A(_09648_),
    .X(net1248));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1250 (.A(_09648_),
    .X(net1249));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1251 (.A(_09352_),
    .X(net1250));
 sky130_fd_sc_hd__buf_2 fanout1252 (.A(_09352_),
    .X(net1251));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1253 (.A(net1254),
    .X(net1252));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1254 (.A(_06023_),
    .X(net1253));
 sky130_fd_sc_hd__buf_12 wire1255 (.A(_06023_),
    .X(net1254));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1256 (.A(net1257),
    .X(net1255));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1257 (.A(_06018_),
    .X(net1256));
 sky130_fd_sc_hd__buf_16 wire1258 (.A(net1256),
    .X(net1257));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1259 (.A(net1261),
    .X(net1258));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1260 (.A(net1261),
    .X(net1259));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1261 (.A(_05972_),
    .X(net1260));
 sky130_fd_sc_hd__buf_12 wire1262 (.A(net1260),
    .X(net1261));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1263 (.A(_05893_),
    .X(net1262));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1264 (.A(_05893_),
    .X(net1263));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1265 (.A(_05826_),
    .X(net1264));
 sky130_fd_sc_hd__buf_2 fanout1266 (.A(_05813_),
    .X(net1265));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1267 (.A(_05813_),
    .X(net1266));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1268 (.A(net1269),
    .X(net1267));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1269 (.A(_05794_),
    .X(net1268));
 sky130_fd_sc_hd__buf_16 wire1270 (.A(net1268),
    .X(net1269));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1271 (.A(net1271),
    .X(net1270));
 sky130_fd_sc_hd__buf_2 fanout1272 (.A(_05773_),
    .X(net1271));
 sky130_fd_sc_hd__buf_2 fanout1273 (.A(_05773_),
    .X(net1272));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1274 (.A(net1277),
    .X(net1273));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1275 (.A(net1275),
    .X(net1274));
 sky130_fd_sc_hd__buf_2 fanout1276 (.A(net1277),
    .X(net1275));
 sky130_fd_sc_hd__buf_16 max_cap1277 (.A(net1275),
    .X(net1276));
 sky130_fd_sc_hd__buf_4 wire1278 (.A(_05754_),
    .X(net1277));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1279 (.A(_05715_),
    .X(net1278));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1280 (.A(net1282),
    .X(net1279));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1281 (.A(_05715_),
    .X(net1280));
 sky130_fd_sc_hd__buf_16 wire1282 (.A(net1280),
    .X(net1281));
 sky130_fd_sc_hd__buf_16 load_slew1283 (.A(net1280),
    .X(net1282));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1284 (.A(net1285),
    .X(net1283));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1285 (.A(net1285),
    .X(net1284));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1286 (.A(_05693_),
    .X(net1285));
 sky130_fd_sc_hd__buf_12 wire1287 (.A(net1285),
    .X(net1286));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1288 (.A(net1291),
    .X(net1287));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1289 (.A(net1290),
    .X(net1288));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1290 (.A(_05671_),
    .X(net1289));
 sky130_fd_sc_hd__buf_12 wire1291 (.A(net1289),
    .X(net1290));
 sky130_fd_sc_hd__buf_16 load_slew1292 (.A(_05671_),
    .X(net1291));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1293 (.A(net1294),
    .X(net1292));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1294 (.A(net1294),
    .X(net1293));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1295 (.A(net1295),
    .X(net1294));
 sky130_fd_sc_hd__buf_2 fanout1296 (.A(_05649_),
    .X(net1295));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1297 (.A(net1298),
    .X(net1296));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1298 (.A(net1298),
    .X(net1297));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1299 (.A(net1299),
    .X(net1298));
 sky130_fd_sc_hd__buf_2 fanout1300 (.A(_05627_),
    .X(net1299));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1301 (.A(net1304),
    .X(net1300));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1302 (.A(net1302),
    .X(net1301));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1303 (.A(net1304),
    .X(net1302));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1304 (.A(_05603_),
    .X(net1303));
 sky130_fd_sc_hd__buf_16 load_slew1305 (.A(net1303),
    .X(net1304));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1306 (.A(net1306),
    .X(net1305));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1307 (.A(net1307),
    .X(net1306));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1308 (.A(net1308),
    .X(net1307));
 sky130_fd_sc_hd__buf_2 fanout1309 (.A(_20812_),
    .X(net1308));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1310 (.A(net1310),
    .X(net1309));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1311 (.A(net1311),
    .X(net1310));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1312 (.A(net1312),
    .X(net1311));
 sky130_fd_sc_hd__buf_2 fanout1313 (.A(net1313),
    .X(net1312));
 sky130_fd_sc_hd__buf_2 wire1314 (.A(_20794_),
    .X(net1313));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1315 (.A(net1315),
    .X(net1314));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1316 (.A(net1316),
    .X(net1315));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1317 (.A(net1317),
    .X(net1316));
 sky130_fd_sc_hd__buf_2 fanout1318 (.A(_20776_),
    .X(net1317));
 sky130_fd_sc_hd__buf_12 wire1319 (.A(_20759_),
    .X(net1318));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1320 (.A(net1320),
    .X(net1319));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1321 (.A(net1321),
    .X(net1320));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1322 (.A(net1322),
    .X(net1321));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1323 (.A(_20756_),
    .X(net1322));
 sky130_fd_sc_hd__buf_12 load_slew1324 (.A(_20734_),
    .X(net1323));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1325 (.A(net1325),
    .X(net1324));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1326 (.A(net1326),
    .X(net1325));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1327 (.A(net1327),
    .X(net1326));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1328 (.A(_20731_),
    .X(net1327));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1329 (.A(net1329),
    .X(net1328));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1330 (.A(net1330),
    .X(net1329));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1331 (.A(net1331),
    .X(net1330));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1332 (.A(_20710_),
    .X(net1331));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1333 (.A(net1334),
    .X(net1332));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1334 (.A(net1334),
    .X(net1333));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1335 (.A(net1335),
    .X(net1334));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1336 (.A(net1337),
    .X(net1335));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1337 (.A(_20690_),
    .X(net1336));
 sky130_fd_sc_hd__buf_16 wire1338 (.A(net1336),
    .X(net1337));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1339 (.A(net1339),
    .X(net1338));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1340 (.A(net1340),
    .X(net1339));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1341 (.A(net1341),
    .X(net1340));
 sky130_fd_sc_hd__buf_2 fanout1342 (.A(_20670_),
    .X(net1341));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1343 (.A(net1343),
    .X(net1342));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1344 (.A(net1344),
    .X(net1343));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1345 (.A(net1346),
    .X(net1344));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1346 (.A(_20628_),
    .X(net1345));
 sky130_fd_sc_hd__buf_16 wire1347 (.A(net1345),
    .X(net1346));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1348 (.A(net1348),
    .X(net1347));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1349 (.A(net1349),
    .X(net1348));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1350 (.A(_20599_),
    .X(net1349));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1351 (.A(_20599_),
    .X(net1350));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1352 (.A(net1355),
    .X(net1351));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1353 (.A(net1354),
    .X(net1352));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1354 (.A(net1354),
    .X(net1353));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1355 (.A(net1355),
    .X(net1354));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1356 (.A(_20571_),
    .X(net1355));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1357 (.A(_20543_),
    .X(net1356));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1358 (.A(_20543_),
    .X(net1357));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1359 (.A(net1359),
    .X(net1358));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1360 (.A(net1360),
    .X(net1359));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1361 (.A(_20543_),
    .X(net1360));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1362 (.A(_20505_),
    .X(net1361));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1363 (.A(_20505_),
    .X(net1362));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1364 (.A(net1364),
    .X(net1363));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1365 (.A(net1365),
    .X(net1364));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1366 (.A(_20505_),
    .X(net1365));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1367 (.A(net1367),
    .X(net1366));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1368 (.A(_20464_),
    .X(net1367));
 sky130_fd_sc_hd__buf_16 wire1369 (.A(net1367),
    .X(net1368));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1370 (.A(_00136_),
    .X(net1369));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1371 (.A(_00136_),
    .X(net1370));
 sky130_fd_sc_hd__buf_2 fanout1372 (.A(_00136_),
    .X(net1371));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1373 (.A(_00136_),
    .X(net1372));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1374 (.A(net1374),
    .X(net1373));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1375 (.A(net1376),
    .X(net1374));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1376 (.A(_00156_),
    .X(net1375));
 sky130_fd_sc_hd__buf_16 wire1377 (.A(_00156_),
    .X(net1376));
 sky130_fd_sc_hd__buf_2 fanout1378 (.A(net1380),
    .X(net1377));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1379 (.A(net1379),
    .X(net1378));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1380 (.A(net1380),
    .X(net1379));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1381 (.A(_00129_),
    .X(net1380));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1382 (.A(_20167_),
    .X(net1381));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1383 (.A(net1384),
    .X(net1382));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1384 (.A(net1384),
    .X(net1383));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1385 (.A(net1385),
    .X(net1384));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1386 (.A(_20130_),
    .X(net1385));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1387 (.A(net1387),
    .X(net1386));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1388 (.A(net1388),
    .X(net1387));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1389 (.A(net1389),
    .X(net1388));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1390 (.A(_20115_),
    .X(net1389));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1391 (.A(net1392),
    .X(net1390));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1392 (.A(net1392),
    .X(net1391));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1393 (.A(net1393),
    .X(net1392));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1394 (.A(net1394),
    .X(net1393));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1395 (.A(_20107_),
    .X(net1394));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1396 (.A(net1396),
    .X(net1395));
 sky130_fd_sc_hd__buf_2 fanout1397 (.A(_20092_),
    .X(net1396));
 sky130_fd_sc_hd__buf_12 wire1398 (.A(_20086_),
    .X(net1397));
 sky130_fd_sc_hd__buf_12 wire1399 (.A(_20080_),
    .X(net1398));
 sky130_fd_sc_hd__buf_2 fanout1400 (.A(net1402),
    .X(net1399));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1401 (.A(net1401),
    .X(net1400));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1402 (.A(net1402),
    .X(net1401));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1403 (.A(_20074_),
    .X(net1402));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1404 (.A(net1406),
    .X(net1403));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1405 (.A(net1405),
    .X(net1404));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1406 (.A(net1406),
    .X(net1405));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1407 (.A(_20068_),
    .X(net1406));
 sky130_fd_sc_hd__buf_12 load_slew1408 (.A(_20061_),
    .X(net1407));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1409 (.A(net1409),
    .X(net1408));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1410 (.A(net1410),
    .X(net1409));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1411 (.A(net1411),
    .X(net1410));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1412 (.A(_20055_),
    .X(net1411));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1413 (.A(net1413),
    .X(net1412));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1414 (.A(net1414),
    .X(net1413));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1415 (.A(net1415),
    .X(net1414));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1416 (.A(net1416),
    .X(net1415));
 sky130_fd_sc_hd__buf_4 wire1417 (.A(_20048_),
    .X(net1416));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1418 (.A(net1418),
    .X(net1417));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1419 (.A(net1419),
    .X(net1418));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1420 (.A(net1420),
    .X(net1419));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1421 (.A(_20042_),
    .X(net1420));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1422 (.A(net1422),
    .X(net1421));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1423 (.A(net1423),
    .X(net1422));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1424 (.A(net1424),
    .X(net1423));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1425 (.A(_20036_),
    .X(net1424));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1426 (.A(net1426),
    .X(net1425));
 sky130_fd_sc_hd__buf_2 fanout1427 (.A(_20030_),
    .X(net1426));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1428 (.A(_20024_),
    .X(net1427));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1429 (.A(_20019_),
    .X(net1428));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1430 (.A(net1430),
    .X(net1429));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1431 (.A(net1431),
    .X(net1430));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1432 (.A(_20014_),
    .X(net1431));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1433 (.A(net1433),
    .X(net1432));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1434 (.A(net1434),
    .X(net1433));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1435 (.A(net1436),
    .X(net1434));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1436 (.A(_20009_),
    .X(net1435));
 sky130_fd_sc_hd__buf_12 wire1437 (.A(net1435),
    .X(net1436));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1438 (.A(_19997_),
    .X(net1437));
 sky130_fd_sc_hd__buf_16 wire1439 (.A(net1437),
    .X(net1438));
 sky130_fd_sc_hd__buf_16 load_slew1440 (.A(_19997_),
    .X(net1439));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1441 (.A(net1442),
    .X(net1440));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1442 (.A(net1442),
    .X(net1441));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1443 (.A(net1443),
    .X(net1442));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1444 (.A(_19990_),
    .X(net1443));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1445 (.A(net1446),
    .X(net1444));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1446 (.A(net1446),
    .X(net1445));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1447 (.A(net1447),
    .X(net1446));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1448 (.A(net1448),
    .X(net1447));
 sky130_fd_sc_hd__buf_6 wire1449 (.A(_19983_),
    .X(net1448));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1450 (.A(net1450),
    .X(net1449));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1451 (.A(net1451),
    .X(net1450));
 sky130_fd_sc_hd__buf_12 wire1452 (.A(_19973_),
    .X(net1451));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1453 (.A(_19952_),
    .X(net1452));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1454 (.A(_19952_),
    .X(net1453));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1455 (.A(net1455),
    .X(net1454));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1456 (.A(net1456),
    .X(net1455));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1457 (.A(net1457),
    .X(net1456));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1458 (.A(net1458),
    .X(net1457));
 sky130_fd_sc_hd__buf_4 wire1459 (.A(_19944_),
    .X(net1458));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1460 (.A(net1461),
    .X(net1459));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1461 (.A(_19938_),
    .X(net1460));
 sky130_fd_sc_hd__buf_16 wire1462 (.A(net1460),
    .X(net1461));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1463 (.A(net1463),
    .X(net1462));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1464 (.A(net1464),
    .X(net1463));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1465 (.A(net1465),
    .X(net1464));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1466 (.A(_19930_),
    .X(net1465));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1467 (.A(net1469),
    .X(net1466));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1468 (.A(_19924_),
    .X(net1467));
 sky130_fd_sc_hd__buf_8 load_slew1469 (.A(net1467),
    .X(net1468));
 sky130_fd_sc_hd__buf_8 load_slew1470 (.A(net1467),
    .X(net1469));
 sky130_fd_sc_hd__buf_16 wire1471 (.A(_19924_),
    .X(net1470));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1472 (.A(net1472),
    .X(net1471));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1473 (.A(net1473),
    .X(net1472));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1474 (.A(net1474),
    .X(net1473));
 sky130_fd_sc_hd__buf_12 wire1475 (.A(_19918_),
    .X(net1474));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1476 (.A(_19910_),
    .X(net1475));
 sky130_fd_sc_hd__buf_16 wire1477 (.A(net1475),
    .X(net1476));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1478 (.A(_19910_),
    .X(net1477));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1479 (.A(net1479),
    .X(net1478));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1480 (.A(net1480),
    .X(net1479));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1481 (.A(_19899_),
    .X(net1480));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1482 (.A(net1483),
    .X(net1481));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1483 (.A(_19883_),
    .X(net1482));
 sky130_fd_sc_hd__buf_16 load_slew1484 (.A(_19883_),
    .X(net1483));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1485 (.A(net1485),
    .X(net1484));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1486 (.A(net1487),
    .X(net1485));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1487 (.A(_00155_),
    .X(net1486));
 sky130_fd_sc_hd__buf_16 wire1488 (.A(_00155_),
    .X(net1487));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1489 (.A(_00137_),
    .X(net1488));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1490 (.A(_00137_),
    .X(net1489));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1491 (.A(_00137_),
    .X(net1490));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1492 (.A(_00137_),
    .X(net1491));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1493 (.A(_00138_),
    .X(net1492));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1494 (.A(_00138_),
    .X(net1493));
 sky130_fd_sc_hd__buf_2 fanout1495 (.A(_00138_),
    .X(net1494));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1496 (.A(_00138_),
    .X(net1495));
 sky130_fd_sc_hd__buf_2 fanout1497 (.A(_00139_),
    .X(net1496));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1498 (.A(_00139_),
    .X(net1497));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1499 (.A(_00139_),
    .X(net1498));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1500 (.A(_00139_),
    .X(net1499));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1501 (.A(_00141_),
    .X(net1500));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1502 (.A(_00141_),
    .X(net1501));
 sky130_fd_sc_hd__buf_2 fanout1503 (.A(_00141_),
    .X(net1502));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1504 (.A(_00141_),
    .X(net1503));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1505 (.A(_00142_),
    .X(net1504));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1506 (.A(_00142_),
    .X(net1505));
 sky130_fd_sc_hd__buf_2 fanout1507 (.A(_00142_),
    .X(net1506));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1508 (.A(_00142_),
    .X(net1507));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1509 (.A(_00143_),
    .X(net1508));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1510 (.A(_00143_),
    .X(net1509));
 sky130_fd_sc_hd__buf_2 fanout1511 (.A(_00143_),
    .X(net1510));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1512 (.A(_00143_),
    .X(net1511));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1513 (.A(_00144_),
    .X(net1512));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1514 (.A(_00144_),
    .X(net1513));
 sky130_fd_sc_hd__buf_2 fanout1515 (.A(_00144_),
    .X(net1514));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1516 (.A(_00144_),
    .X(net1515));
 sky130_fd_sc_hd__buf_2 fanout1517 (.A(net1519),
    .X(net1516));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1518 (.A(net1518),
    .X(net1517));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1519 (.A(net1519),
    .X(net1518));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1520 (.A(_00145_),
    .X(net1519));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1521 (.A(net1523),
    .X(net1520));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1522 (.A(net1522),
    .X(net1521));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1523 (.A(net1523),
    .X(net1522));
 sky130_fd_sc_hd__buf_2 fanout1524 (.A(_00146_),
    .X(net1523));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1525 (.A(net1527),
    .X(net1524));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1526 (.A(net1526),
    .X(net1525));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1527 (.A(net1527),
    .X(net1526));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1528 (.A(_00147_),
    .X(net1527));
 sky130_fd_sc_hd__buf_2 fanout1529 (.A(net1531),
    .X(net1528));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1530 (.A(net1530),
    .X(net1529));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1531 (.A(net1531),
    .X(net1530));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1532 (.A(_00148_),
    .X(net1531));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1533 (.A(net1535),
    .X(net1532));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1534 (.A(net1534),
    .X(net1533));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1535 (.A(net1535),
    .X(net1534));
 sky130_fd_sc_hd__buf_2 fanout1536 (.A(_00149_),
    .X(net1535));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1537 (.A(net1539),
    .X(net1536));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1538 (.A(net1538),
    .X(net1537));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1539 (.A(net1539),
    .X(net1538));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1540 (.A(_00150_),
    .X(net1539));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1541 (.A(net1543),
    .X(net1540));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1542 (.A(net1542),
    .X(net1541));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1543 (.A(net1543),
    .X(net1542));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1544 (.A(_00152_),
    .X(net1543));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1545 (.A(net1547),
    .X(net1544));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1546 (.A(net1546),
    .X(net1545));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1547 (.A(net1547),
    .X(net1546));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1548 (.A(_00153_),
    .X(net1547));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1549 (.A(net1551),
    .X(net1548));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1550 (.A(net1551),
    .X(net1549));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1551 (.A(_00157_),
    .X(net1550));
 sky130_fd_sc_hd__buf_16 wire1552 (.A(_00157_),
    .X(net1551));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1553 (.A(net1555),
    .X(net1552));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1554 (.A(net1555),
    .X(net1553));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1555 (.A(net1555),
    .X(net1554));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1556 (.A(_00135_),
    .X(net1555));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1557 (.A(net1559),
    .X(net1556));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1558 (.A(net1559),
    .X(net1557));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1559 (.A(_00154_),
    .X(net1558));
 sky130_fd_sc_hd__buf_8 load_slew1560 (.A(_00154_),
    .X(net1559));
 sky130_fd_sc_hd__buf_2 fanout1561 (.A(net1563),
    .X(net1560));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1562 (.A(net1562),
    .X(net1561));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1563 (.A(net1563),
    .X(net1562));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1564 (.A(_00131_),
    .X(net1563));
 sky130_fd_sc_hd__buf_2 fanout1565 (.A(net1567),
    .X(net1564));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1566 (.A(net1566),
    .X(net1565));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1567 (.A(net1567),
    .X(net1566));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1568 (.A(_00130_),
    .X(net1567));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1569 (.A(net1569),
    .X(net1568));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1570 (.A(net1571),
    .X(net1569));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1571 (.A(_00158_),
    .X(net1570));
 sky130_fd_sc_hd__buf_16 wire1572 (.A(_00158_),
    .X(net1571));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1573 (.A(net1575),
    .X(net1572));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1574 (.A(net1574),
    .X(net1573));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1575 (.A(net1575),
    .X(net1574));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1576 (.A(_00160_),
    .X(net1575));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1577 (.A(net1579),
    .X(net1576));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1578 (.A(net1579),
    .X(net1577));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1579 (.A(_00140_),
    .X(net1578));
 sky130_fd_sc_hd__buf_8 wire1580 (.A(_00140_),
    .X(net1579));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1581 (.A(net1583),
    .X(net1580));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1582 (.A(net1582),
    .X(net1581));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1583 (.A(net1583),
    .X(net1582));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1584 (.A(_00132_),
    .X(net1583));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1585 (.A(net1587),
    .X(net1584));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1586 (.A(net1586),
    .X(net1585));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1587 (.A(net1587),
    .X(net1586));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1588 (.A(_00159_),
    .X(net1587));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1589 (.A(net1592),
    .X(net1588));
 sky130_fd_sc_hd__buf_16 max_cap1590 (.A(net1588),
    .X(net1589));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1591 (.A(net1591),
    .X(net1590));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1592 (.A(net1592),
    .X(net1591));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1593 (.A(_00134_),
    .X(net1592));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1594 (.A(net1596),
    .X(net1593));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1595 (.A(net1595),
    .X(net1594));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1596 (.A(net1596),
    .X(net1595));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1597 (.A(_00151_),
    .X(net1596));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1598 (.A(net1600),
    .X(net1597));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1599 (.A(net1599),
    .X(net1598));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1600 (.A(net1600),
    .X(net1599));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1601 (.A(_00133_),
    .X(net1600));
 sky130_fd_sc_hd__buf_16 wire1602 (.A(net559),
    .X(net1601));
 sky130_fd_sc_hd__buf_16 wire1603 (.A(net1603),
    .X(net1602));
 sky130_fd_sc_hd__buf_16 wire1604 (.A(net1604),
    .X(net1603));
 sky130_fd_sc_hd__buf_16 wire1605 (.A(net1605),
    .X(net1604));
 sky130_fd_sc_hd__buf_12 wire1606 (.A(net555),
    .X(net1605));
 sky130_fd_sc_hd__buf_16 wire1607 (.A(net1607),
    .X(net1606));
 sky130_fd_sc_hd__buf_16 wire1608 (.A(net1608),
    .X(net1607));
 sky130_fd_sc_hd__buf_16 wire1609 (.A(net1609),
    .X(net1608));
 sky130_fd_sc_hd__buf_12 wire1610 (.A(net554),
    .X(net1609));
 sky130_fd_sc_hd__buf_16 wire1611 (.A(net558),
    .X(net1610));
 sky130_fd_sc_hd__buf_16 wire1612 (.A(net1612),
    .X(net1611));
 sky130_fd_sc_hd__buf_16 wire1613 (.A(net1613),
    .X(net1612));
 sky130_fd_sc_hd__buf_16 wire1614 (.A(net1614),
    .X(net1613));
 sky130_fd_sc_hd__buf_12 wire1615 (.A(net553),
    .X(net1614));
 sky130_fd_sc_hd__buf_16 wire1616 (.A(net1616),
    .X(net1615));
 sky130_fd_sc_hd__buf_16 wire1617 (.A(net1617),
    .X(net1616));
 sky130_fd_sc_hd__buf_16 wire1618 (.A(net1618),
    .X(net1617));
 sky130_fd_sc_hd__buf_12 wire1619 (.A(net552),
    .X(net1618));
 sky130_fd_sc_hd__buf_16 wire1620 (.A(net1620),
    .X(net1619));
 sky130_fd_sc_hd__buf_16 wire1621 (.A(net1621),
    .X(net1620));
 sky130_fd_sc_hd__buf_12 wire1622 (.A(net551),
    .X(net1621));
 sky130_fd_sc_hd__buf_16 wire1623 (.A(net1623),
    .X(net1622));
 sky130_fd_sc_hd__buf_16 wire1624 (.A(net1624),
    .X(net1623));
 sky130_fd_sc_hd__buf_12 wire1625 (.A(net550),
    .X(net1624));
 sky130_fd_sc_hd__buf_16 wire1626 (.A(net1626),
    .X(net1625));
 sky130_fd_sc_hd__buf_16 wire1627 (.A(net1627),
    .X(net1626));
 sky130_fd_sc_hd__buf_12 wire1628 (.A(net565),
    .X(net1627));
 sky130_fd_sc_hd__buf_16 wire1629 (.A(net1629),
    .X(net1628));
 sky130_fd_sc_hd__buf_16 wire1630 (.A(net1630),
    .X(net1629));
 sky130_fd_sc_hd__buf_12 wire1631 (.A(net564),
    .X(net1630));
 sky130_fd_sc_hd__buf_16 wire1632 (.A(net557),
    .X(net1631));
 sky130_fd_sc_hd__buf_16 wire1633 (.A(net1633),
    .X(net1632));
 sky130_fd_sc_hd__buf_12 wire1634 (.A(net556),
    .X(net1633));
 sky130_fd_sc_hd__buf_2 wire1635 (.A(_19737_),
    .X(net1634));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1636 (.A(net1636),
    .X(net1635));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1637 (.A(_18755_),
    .X(net1636));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1638 (.A(_18755_),
    .X(net1637));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1639 (.A(_18327_),
    .X(net1638));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1640 (.A(_14886_),
    .X(net1639));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1641 (.A(_14886_),
    .X(net1640));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1642 (.A(net1642),
    .X(net1641));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1643 (.A(net1648),
    .X(net1642));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1644 (.A(net1644),
    .X(net1643));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1645 (.A(net1648),
    .X(net1644));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1646 (.A(net1647),
    .X(net1645));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1647 (.A(net1647),
    .X(net1646));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1648 (.A(net1648),
    .X(net1647));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1649 (.A(_11516_),
    .X(net1648));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1650 (.A(_11295_),
    .X(net1649));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1651 (.A(_11295_),
    .X(net1650));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1652 (.A(_11295_),
    .X(net1651));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1653 (.A(_11295_),
    .X(net1652));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1654 (.A(net1654),
    .X(net1653));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1655 (.A(_11243_),
    .X(net1654));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1656 (.A(_11243_),
    .X(net1655));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1657 (.A(net1657),
    .X(net1656));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1658 (.A(net1659),
    .X(net1657));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1659 (.A(net1659),
    .X(net1658));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1660 (.A(_11243_),
    .X(net1659));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1661 (.A(net1662),
    .X(net1660));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1662 (.A(net1662),
    .X(net1661));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1663 (.A(net1663),
    .X(net1662));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1664 (.A(_11145_),
    .X(net1663));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1665 (.A(net1666),
    .X(net1664));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1666 (.A(_09906_),
    .X(net1665));
 sky130_fd_sc_hd__buf_4 wire1667 (.A(_09906_),
    .X(net1666));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1668 (.A(net1668),
    .X(net1667));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1669 (.A(_07483_),
    .X(net1668));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1670 (.A(net1670),
    .X(net1669));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1671 (.A(_05811_),
    .X(net1670));
 sky130_fd_sc_hd__buf_16 wire1672 (.A(_05811_),
    .X(net1671));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1673 (.A(net1676),
    .X(net1672));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1674 (.A(net1675),
    .X(net1673));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1675 (.A(net1676),
    .X(net1674));
 sky130_fd_sc_hd__buf_16 load_slew1676 (.A(net1674),
    .X(net1675));
 sky130_fd_sc_hd__buf_8 wire1677 (.A(_05792_),
    .X(net1676));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1678 (.A(net3044),
    .X(net1677));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1679 (.A(_05732_),
    .X(net1678));
 sky130_fd_sc_hd__buf_16 wire1680 (.A(_05732_),
    .X(net1679));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1681 (.A(net1681),
    .X(net1680));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1682 (.A(_05619_),
    .X(net1681));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1683 (.A(net1683),
    .X(net1682));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1684 (.A(net1684),
    .X(net1683));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1685 (.A(_20378_),
    .X(net1684));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1686 (.A(net1686),
    .X(net1685));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1687 (.A(net1689),
    .X(net1686));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1688 (.A(net1689),
    .X(net1687));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1689 (.A(net1689),
    .X(net1688));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1690 (.A(net1690),
    .X(net1689));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1691 (.A(_20378_),
    .X(net1690));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1692 (.A(net1692),
    .X(net1691));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1693 (.A(net1693),
    .X(net1692));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1694 (.A(net1696),
    .X(net1693));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1695 (.A(net1695),
    .X(net1694));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1696 (.A(net1696),
    .X(net1695));
 sky130_fd_sc_hd__buf_6 wire1697 (.A(_20137_),
    .X(net1696));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1698 (.A(net1698),
    .X(net1697));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1699 (.A(net1699),
    .X(net1698));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1700 (.A(_20129_),
    .X(net1699));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1701 (.A(net1701),
    .X(net1700));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1702 (.A(net1705),
    .X(net1701));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1703 (.A(net1703),
    .X(net1702));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1704 (.A(net1704),
    .X(net1703));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1705 (.A(net1705),
    .X(net1704));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1706 (.A(_20129_),
    .X(net1705));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1707 (.A(net1707),
    .X(net1706));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1708 (.A(_20124_),
    .X(net1707));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1709 (.A(_20124_),
    .X(net1708));
 sky130_fd_sc_hd__buf_12 wire1710 (.A(_20067_),
    .X(net1709));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1711 (.A(net1711),
    .X(net1710));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1712 (.A(net1712),
    .X(net1711));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1713 (.A(net1713),
    .X(net1712));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1714 (.A(_20029_),
    .X(net1713));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1715 (.A(net1715),
    .X(net1714));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1716 (.A(net1716),
    .X(net1715));
 sky130_fd_sc_hd__buf_2 fanout1717 (.A(_20023_),
    .X(net1716));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1718 (.A(net1718),
    .X(net1717));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1719 (.A(net1719),
    .X(net1718));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1720 (.A(_20018_),
    .X(net1719));
 sky130_fd_sc_hd__buf_16 load_slew1721 (.A(net1721),
    .X(net1720));
 sky130_fd_sc_hd__buf_8 load_slew1722 (.A(net1719),
    .X(net1721));
 sky130_fd_sc_hd__buf_12 wire1723 (.A(_20013_),
    .X(net1722));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1724 (.A(net1726),
    .X(net1723));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1725 (.A(net1726),
    .X(net1724));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1726 (.A(_19967_),
    .X(net1725));
 sky130_fd_sc_hd__buf_12 wire1727 (.A(net1725),
    .X(net1726));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1728 (.A(net1730),
    .X(net1727));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1729 (.A(net1730),
    .X(net1728));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1730 (.A(_19962_),
    .X(net1729));
 sky130_fd_sc_hd__buf_16 wire1731 (.A(net1729),
    .X(net1730));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1732 (.A(net1732),
    .X(net1731));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1733 (.A(net1733),
    .X(net1732));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1734 (.A(net1734),
    .X(net1733));
 sky130_fd_sc_hd__buf_12 wire1735 (.A(_19957_),
    .X(net1734));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1736 (.A(net1737),
    .X(net1735));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1737 (.A(net1738),
    .X(net1736));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1738 (.A(_19937_),
    .X(net1737));
 sky130_fd_sc_hd__buf_16 load_slew1739 (.A(net1737),
    .X(net1738));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1740 (.A(net1740),
    .X(net1739));
 sky130_fd_sc_hd__buf_2 fanout1741 (.A(_19898_),
    .X(net1740));
 sky130_fd_sc_hd__buf_16 wire1742 (.A(net593),
    .X(net1741));
 sky130_fd_sc_hd__buf_16 wire1743 (.A(net592),
    .X(net1742));
 sky130_fd_sc_hd__buf_16 wire1744 (.A(net591),
    .X(net1743));
 sky130_fd_sc_hd__buf_16 wire1745 (.A(net590),
    .X(net1744));
 sky130_fd_sc_hd__buf_16 wire1746 (.A(net588),
    .X(net1745));
 sky130_fd_sc_hd__buf_16 wire1747 (.A(net585),
    .X(net1746));
 sky130_fd_sc_hd__buf_16 wire1748 (.A(net1748),
    .X(net1747));
 sky130_fd_sc_hd__buf_16 wire1749 (.A(net1749),
    .X(net1748));
 sky130_fd_sc_hd__buf_16 wire1750 (.A(net584),
    .X(net1749));
 sky130_fd_sc_hd__buf_16 wire1751 (.A(net1751),
    .X(net1750));
 sky130_fd_sc_hd__buf_16 wire1752 (.A(net1752),
    .X(net1751));
 sky130_fd_sc_hd__buf_16 wire1753 (.A(net583),
    .X(net1752));
 sky130_fd_sc_hd__buf_16 wire1754 (.A(net1754),
    .X(net1753));
 sky130_fd_sc_hd__buf_16 wire1755 (.A(net1755),
    .X(net1754));
 sky130_fd_sc_hd__buf_16 wire1756 (.A(net600),
    .X(net1755));
 sky130_fd_sc_hd__buf_16 wire1757 (.A(net1757),
    .X(net1756));
 sky130_fd_sc_hd__buf_16 wire1758 (.A(net599),
    .X(net1757));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1759 (.A(_19111_),
    .X(net1758));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1760 (.A(_19111_),
    .X(net1759));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1761 (.A(_19049_),
    .X(net1760));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1762 (.A(_19049_),
    .X(net1761));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1763 (.A(net1765),
    .X(net1762));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1764 (.A(net1765),
    .X(net1763));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1765 (.A(net1765),
    .X(net1764));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1766 (.A(_18768_),
    .X(net1765));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1767 (.A(_18756_),
    .X(net1766));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1768 (.A(_15006_),
    .X(net1767));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1769 (.A(_15006_),
    .X(net1768));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1770 (.A(net1770),
    .X(net1769));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1771 (.A(net1774),
    .X(net1770));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1772 (.A(net1773),
    .X(net1771));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1773 (.A(net1773),
    .X(net1772));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1774 (.A(net1774),
    .X(net1773));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1775 (.A(_15006_),
    .X(net1774));
 sky130_fd_sc_hd__buf_8 wire1776 (.A(_14542_),
    .X(net1775));
 sky130_fd_sc_hd__buf_16 wire1777 (.A(_14514_),
    .X(net1776));
 sky130_fd_sc_hd__buf_6 wire1778 (.A(_14499_),
    .X(net1777));
 sky130_fd_sc_hd__buf_8 wire1779 (.A(_14456_),
    .X(net1778));
 sky130_fd_sc_hd__buf_6 wire1780 (.A(_14397_),
    .X(net1779));
 sky130_fd_sc_hd__buf_6 wire1781 (.A(_14383_),
    .X(net1780));
 sky130_fd_sc_hd__buf_4 wire1782 (.A(_14357_),
    .X(net1781));
 sky130_fd_sc_hd__buf_6 wire1783 (.A(_14247_),
    .X(net1782));
 sky130_fd_sc_hd__buf_6 wire1784 (.A(_14235_),
    .X(net1783));
 sky130_fd_sc_hd__buf_6 wire1785 (.A(_13957_),
    .X(net1784));
 sky130_fd_sc_hd__buf_6 wire1786 (.A(_13908_),
    .X(net1785));
 sky130_fd_sc_hd__buf_6 wire1787 (.A(_13754_),
    .X(net1786));
 sky130_fd_sc_hd__buf_6 wire1788 (.A(_13742_),
    .X(net1787));
 sky130_fd_sc_hd__buf_6 wire1789 (.A(_13674_),
    .X(net1788));
 sky130_fd_sc_hd__buf_6 wire1790 (.A(_13603_),
    .X(net1789));
 sky130_fd_sc_hd__buf_6 wire1791 (.A(_13583_),
    .X(net1790));
 sky130_fd_sc_hd__buf_8 wire1792 (.A(_13531_),
    .X(net1791));
 sky130_fd_sc_hd__buf_16 wire1793 (.A(_13347_),
    .X(net1792));
 sky130_fd_sc_hd__buf_8 wire1794 (.A(_13253_),
    .X(net1793));
 sky130_fd_sc_hd__buf_16 wire1795 (.A(_13237_),
    .X(net1794));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1796 (.A(net1796),
    .X(net1795));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1797 (.A(_12967_),
    .X(net1796));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1798 (.A(_12967_),
    .X(net1797));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1799 (.A(_12967_),
    .X(net1798));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1800 (.A(net1800),
    .X(net1799));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1801 (.A(net1803),
    .X(net1800));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1802 (.A(net1802),
    .X(net1801));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1803 (.A(net1803),
    .X(net1802));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1804 (.A(_12696_),
    .X(net1803));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1805 (.A(net1806),
    .X(net1804));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1806 (.A(net1806),
    .X(net1805));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1807 (.A(_12696_),
    .X(net1806));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1808 (.A(net1808),
    .X(net1807));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1809 (.A(net1810),
    .X(net1808));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1810 (.A(net1810),
    .X(net1809));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1811 (.A(_10911_),
    .X(net1810));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1812 (.A(net1814),
    .X(net1811));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1813 (.A(net1813),
    .X(net1812));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1814 (.A(net1814),
    .X(net1813));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1815 (.A(_10911_),
    .X(net1814));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1816 (.A(net1816),
    .X(net1815));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1817 (.A(net1821),
    .X(net1816));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1818 (.A(net1821),
    .X(net1817));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1819 (.A(net1820),
    .X(net1818));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1820 (.A(net1820),
    .X(net1819));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1821 (.A(net1821),
    .X(net1820));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1822 (.A(_20357_),
    .X(net1821));
 sky130_fd_sc_hd__buf_6 wire1823 (.A(_20001_),
    .X(net1822));
 sky130_fd_sc_hd__buf_6 wire1824 (.A(_19988_),
    .X(net1823));
 sky130_fd_sc_hd__buf_4 wire1825 (.A(_19981_),
    .X(net1824));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1826 (.A(net1826),
    .X(net1825));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1827 (.A(net1827),
    .X(net1826));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1828 (.A(_19976_),
    .X(net1827));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1829 (.A(_19881_),
    .X(net1828));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1830 (.A(net1830),
    .X(net1829));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1831 (.A(_19881_),
    .X(net1830));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1832 (.A(_19872_),
    .X(net1831));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1833 (.A(_19872_),
    .X(net1832));
 sky130_fd_sc_hd__buf_12 load_slew1834 (.A(\inst$top.soc.bus__adr[7] ),
    .X(net1833));
 sky130_fd_sc_hd__buf_12 load_slew1835 (.A(\inst$top.soc.bus__adr[5] ),
    .X(net1834));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1836 (.A(_02882_),
    .X(net1835));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1837 (.A(net1837),
    .X(net1836));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1838 (.A(_02881_),
    .X(net1837));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1839 (.A(_02865_),
    .X(net1838));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1840 (.A(net1840),
    .X(net1839));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1841 (.A(_02865_),
    .X(net1840));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1842 (.A(net1842),
    .X(net1841));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1843 (.A(_19542_),
    .X(net1842));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1844 (.A(net1844),
    .X(net1843));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1845 (.A(_19542_),
    .X(net1844));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1846 (.A(net1847),
    .X(net1845));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1847 (.A(net1847),
    .X(net1846));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1848 (.A(_19394_),
    .X(net1847));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1849 (.A(_19394_),
    .X(net1848));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1850 (.A(_19394_),
    .X(net1849));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1851 (.A(_19167_),
    .X(net1850));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1852 (.A(net1853),
    .X(net1851));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1853 (.A(net1853),
    .X(net1852));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1854 (.A(_19110_),
    .X(net1853));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1855 (.A(net1856),
    .X(net1854));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1856 (.A(net1856),
    .X(net1855));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1857 (.A(_18760_),
    .X(net1856));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1858 (.A(net1860),
    .X(net1857));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1859 (.A(net1860),
    .X(net1858));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1860 (.A(net1860),
    .X(net1859));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1861 (.A(_17148_),
    .X(net1860));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1862 (.A(_17034_),
    .X(net1861));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1863 (.A(net1863),
    .X(net1862));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1864 (.A(_17034_),
    .X(net1863));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1865 (.A(net1867),
    .X(net1864));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1866 (.A(net1867),
    .X(net1865));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1867 (.A(net1867),
    .X(net1866));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1868 (.A(_17034_),
    .X(net1867));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1869 (.A(net1869),
    .X(net1868));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1870 (.A(_12971_),
    .X(net1869));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1871 (.A(_12971_),
    .X(net1870));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1872 (.A(_12971_),
    .X(net1871));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1873 (.A(net1873),
    .X(net1872));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1874 (.A(_10921_),
    .X(net1873));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1875 (.A(net1875),
    .X(net1874));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1876 (.A(_10921_),
    .X(net1875));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1877 (.A(net1880),
    .X(net1876));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1878 (.A(net1878),
    .X(net1877));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1879 (.A(net1880),
    .X(net1878));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1880 (.A(net1880),
    .X(net1879));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1881 (.A(_10921_),
    .X(net1880));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1882 (.A(net1882),
    .X(net1881));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1883 (.A(net1886),
    .X(net1882));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1884 (.A(net1884),
    .X(net1883));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1885 (.A(net1885),
    .X(net1884));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1886 (.A(net1886),
    .X(net1885));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1887 (.A(net1893),
    .X(net1886));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1888 (.A(net1890),
    .X(net1887));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1889 (.A(net1890),
    .X(net1888));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1890 (.A(net1890),
    .X(net1889));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1891 (.A(net1893),
    .X(net1890));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1892 (.A(net1893),
    .X(net1891));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1893 (.A(net1893),
    .X(net1892));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1894 (.A(net1909),
    .X(net1893));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1895 (.A(net1895),
    .X(net1894));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1896 (.A(net1900),
    .X(net1895));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1897 (.A(net1900),
    .X(net1896));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1898 (.A(net1899),
    .X(net1897));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1899 (.A(net1899),
    .X(net1898));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1900 (.A(net1900),
    .X(net1899));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1901 (.A(net1909),
    .X(net1900));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1902 (.A(net1904),
    .X(net1901));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1903 (.A(net1904),
    .X(net1902));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1904 (.A(net1904),
    .X(net1903));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1905 (.A(net1909),
    .X(net1904));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1906 (.A(net1906),
    .X(net1905));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1907 (.A(net1909),
    .X(net1906));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1908 (.A(net1908),
    .X(net1907));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1909 (.A(net1909),
    .X(net1908));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1910 (.A(net1932),
    .X(net1909));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1911 (.A(net1912),
    .X(net1910));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1912 (.A(net1912),
    .X(net1911));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1913 (.A(net1913),
    .X(net1912));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1914 (.A(net1923),
    .X(net1913));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1915 (.A(net1915),
    .X(net1914));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1916 (.A(net1918),
    .X(net1915));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1917 (.A(net1917),
    .X(net1916));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1918 (.A(net1918),
    .X(net1917));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1919 (.A(net1923),
    .X(net1918));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1920 (.A(net1920),
    .X(net1919));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1921 (.A(net1921),
    .X(net1920));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1922 (.A(net1923),
    .X(net1921));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1923 (.A(net1923),
    .X(net1922));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1924 (.A(net1932),
    .X(net1923));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1925 (.A(net1925),
    .X(net1924));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1926 (.A(net1933),
    .X(net1925));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1927 (.A(net1927),
    .X(net1926));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1928 (.A(net1933),
    .X(net1927));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1929 (.A(net1929),
    .X(net1928));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1930 (.A(net1931),
    .X(net1929));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1931 (.A(net1931),
    .X(net1930));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1932 (.A(net1933),
    .X(net1931));
 sky130_fd_sc_hd__buf_2 fanout1933 (.A(_09405_),
    .X(net1932));
 sky130_fd_sc_hd__buf_16 wire1934 (.A(net1932),
    .X(net1933));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1935 (.A(net1936),
    .X(net1934));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1936 (.A(net1936),
    .X(net1935));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1937 (.A(net1943),
    .X(net1936));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1938 (.A(net1940),
    .X(net1937));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1939 (.A(net1940),
    .X(net1938));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1940 (.A(net1940),
    .X(net1939));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1941 (.A(net1941),
    .X(net1940));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1942 (.A(_06101_),
    .X(net1941));
 sky130_fd_sc_hd__buf_16 load_slew1943 (.A(net1943),
    .X(net1942));
 sky130_fd_sc_hd__buf_16 load_slew1944 (.A(net1941),
    .X(net1943));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1945 (.A(net1947),
    .X(net1944));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1946 (.A(net1947),
    .X(net1945));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1947 (.A(net1947),
    .X(net1946));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1948 (.A(net1948),
    .X(net1947));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1949 (.A(net1957),
    .X(net1948));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1950 (.A(net1950),
    .X(net1949));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1951 (.A(net1957),
    .X(net1950));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1952 (.A(net1957),
    .X(net1951));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1953 (.A(net1957),
    .X(net1952));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1954 (.A(net1956),
    .X(net1953));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1955 (.A(net1956),
    .X(net1954));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1956 (.A(net1956),
    .X(net1955));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1957 (.A(net1957),
    .X(net1956));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1958 (.A(_06064_),
    .X(net1957));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1959 (.A(net1959),
    .X(net1958));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1960 (.A(net1966),
    .X(net1959));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1961 (.A(net1966),
    .X(net1960));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1962 (.A(net1966),
    .X(net1961));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1963 (.A(net1963),
    .X(net1962));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1964 (.A(net1966),
    .X(net1963));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1965 (.A(net1966),
    .X(net1964));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1966 (.A(net1966),
    .X(net1965));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1967 (.A(_06064_),
    .X(net1966));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1968 (.A(net1976),
    .X(net1967));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1969 (.A(net1976),
    .X(net1968));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1970 (.A(net1970),
    .X(net1969));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1971 (.A(net1976),
    .X(net1970));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1972 (.A(net1972),
    .X(net1971));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1973 (.A(net1975),
    .X(net1972));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1974 (.A(net1975),
    .X(net1973));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1975 (.A(net1975),
    .X(net1974));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1976 (.A(net1976),
    .X(net1975));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1977 (.A(_06064_),
    .X(net1976));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1978 (.A(net1978),
    .X(net1977));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1979 (.A(net1979),
    .X(net1978));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1980 (.A(_20498_),
    .X(net1979));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1981 (.A(net1981),
    .X(net1980));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1982 (.A(_20481_),
    .X(net1981));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1983 (.A(net1985),
    .X(net1982));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1984 (.A(net1985),
    .X(net1983));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1985 (.A(net1985),
    .X(net1984));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1986 (.A(_20403_),
    .X(net1985));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1987 (.A(_19886_),
    .X(net1986));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1988 (.A(net1989),
    .X(net1987));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1989 (.A(net1989),
    .X(net1988));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1990 (.A(_19886_),
    .X(net1989));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1991 (.A(_19134_),
    .X(net1990));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1992 (.A(_19134_),
    .X(net1991));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1993 (.A(_19101_),
    .X(net1992));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1994 (.A(net1996),
    .X(net1993));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1995 (.A(net1995),
    .X(net1994));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1996 (.A(net1996),
    .X(net1995));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1997 (.A(_17147_),
    .X(net1996));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1998 (.A(net1998),
    .X(net1997));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout1999 (.A(net2000),
    .X(net1998));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2000 (.A(net2000),
    .X(net1999));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2001 (.A(_16055_),
    .X(net2000));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2002 (.A(_13129_),
    .X(net2001));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2003 (.A(net2004),
    .X(net2002));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2004 (.A(net2004),
    .X(net2003));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2005 (.A(_13102_),
    .X(net2004));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2006 (.A(net2007),
    .X(net2005));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2007 (.A(net2007),
    .X(net2006));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2008 (.A(net2008),
    .X(net2007));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2009 (.A(_13041_),
    .X(net2008));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2010 (.A(net2011),
    .X(net2009));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2011 (.A(net2011),
    .X(net2010));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2012 (.A(net2012),
    .X(net2011));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2013 (.A(_12994_),
    .X(net2012));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2014 (.A(net2016),
    .X(net2013));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2015 (.A(net2016),
    .X(net2014));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2016 (.A(net2016),
    .X(net2015));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2017 (.A(_12994_),
    .X(net2016));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2018 (.A(net2020),
    .X(net2017));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2019 (.A(net2019),
    .X(net2018));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2020 (.A(net2020),
    .X(net2019));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2021 (.A(_12961_),
    .X(net2020));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2022 (.A(_11194_),
    .X(net2021));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2023 (.A(_11194_),
    .X(net2022));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2024 (.A(net2025),
    .X(net2023));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2025 (.A(net2025),
    .X(net2024));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2026 (.A(net2026),
    .X(net2025));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2027 (.A(_09920_),
    .X(net2026));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2028 (.A(net2028),
    .X(net2027));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2029 (.A(net2082),
    .X(net2028));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2030 (.A(net2030),
    .X(net2029));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2031 (.A(net2036),
    .X(net2030));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2032 (.A(net2035),
    .X(net2031));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2033 (.A(net2035),
    .X(net2032));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2034 (.A(net2035),
    .X(net2033));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2035 (.A(net2035),
    .X(net2034));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2036 (.A(net2036),
    .X(net2035));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2037 (.A(net2082),
    .X(net2036));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2038 (.A(net2046),
    .X(net2037));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2039 (.A(net2046),
    .X(net2038));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2040 (.A(net2041),
    .X(net2039));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2041 (.A(net2041),
    .X(net2040));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2042 (.A(net2046),
    .X(net2041));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2043 (.A(net2046),
    .X(net2042));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2044 (.A(net2046),
    .X(net2043));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2045 (.A(net2046),
    .X(net2044));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2046 (.A(net2046),
    .X(net2045));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2047 (.A(net2082),
    .X(net2046));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2048 (.A(net2048),
    .X(net2047));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2049 (.A(net2050),
    .X(net2048));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2050 (.A(net2050),
    .X(net2049));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2051 (.A(net2064),
    .X(net2050));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2052 (.A(net2052),
    .X(net2051));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2053 (.A(net2053),
    .X(net2052));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2054 (.A(net2058),
    .X(net2053));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2055 (.A(net2058),
    .X(net2054));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2056 (.A(net2058),
    .X(net2055));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2057 (.A(net2058),
    .X(net2056));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2058 (.A(net2058),
    .X(net2057));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2059 (.A(net2064),
    .X(net2058));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2060 (.A(net2064),
    .X(net2059));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2061 (.A(net2064),
    .X(net2060));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2062 (.A(net2063),
    .X(net2061));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2063 (.A(net2063),
    .X(net2062));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2064 (.A(net2064),
    .X(net2063));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2065 (.A(net2082),
    .X(net2064));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2066 (.A(net2066),
    .X(net2065));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2067 (.A(net2072),
    .X(net2066));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2068 (.A(net2072),
    .X(net2067));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2069 (.A(net2072),
    .X(net2068));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2070 (.A(net2072),
    .X(net2069));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2071 (.A(net2071),
    .X(net2070));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2072 (.A(net2072),
    .X(net2071));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2073 (.A(net2082),
    .X(net2072));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2074 (.A(net2075),
    .X(net2073));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2075 (.A(net2075),
    .X(net2074));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2076 (.A(net2081),
    .X(net2075));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2077 (.A(net2077),
    .X(net2076));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2078 (.A(net2081),
    .X(net2077));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2079 (.A(net2079),
    .X(net2078));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2080 (.A(net2081),
    .X(net2079));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2081 (.A(net2081),
    .X(net2080));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2082 (.A(net2082),
    .X(net2081));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2083 (.A(net2188),
    .X(net2082));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2084 (.A(net2084),
    .X(net2083));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2085 (.A(net2089),
    .X(net2084));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2086 (.A(net2089),
    .X(net2085));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2087 (.A(net2089),
    .X(net2086));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2088 (.A(net2088),
    .X(net2087));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2089 (.A(net2089),
    .X(net2088));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2090 (.A(net2103),
    .X(net2089));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2091 (.A(net2091),
    .X(net2090));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2092 (.A(net2092),
    .X(net2091));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2093 (.A(net2103),
    .X(net2092));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2094 (.A(net2094),
    .X(net2093));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2095 (.A(net2102),
    .X(net2094));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2096 (.A(net2096),
    .X(net2095));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2097 (.A(net2102),
    .X(net2096));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2098 (.A(net2102),
    .X(net2097));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2099 (.A(net2101),
    .X(net2098));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2100 (.A(net2100),
    .X(net2099));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2101 (.A(net2101),
    .X(net2100));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2102 (.A(net2102),
    .X(net2101));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2103 (.A(net2103),
    .X(net2102));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2104 (.A(net2118),
    .X(net2103));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2105 (.A(net2108),
    .X(net2104));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2106 (.A(net2108),
    .X(net2105));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2107 (.A(net2108),
    .X(net2106));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2108 (.A(net2108),
    .X(net2107));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2109 (.A(net2114),
    .X(net2108));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2110 (.A(net2110),
    .X(net2109));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2111 (.A(net2114),
    .X(net2110));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2112 (.A(net2112),
    .X(net2111));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2113 (.A(net2114),
    .X(net2112));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2114 (.A(net2114),
    .X(net2113));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2115 (.A(net2118),
    .X(net2114));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2116 (.A(net2117),
    .X(net2115));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2117 (.A(net2117),
    .X(net2116));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2118 (.A(net2118),
    .X(net2117));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2119 (.A(net2188),
    .X(net2118));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2120 (.A(net2125),
    .X(net2119));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2121 (.A(net2125),
    .X(net2120));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2122 (.A(net2124),
    .X(net2121));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2123 (.A(net2124),
    .X(net2122));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2124 (.A(net2124),
    .X(net2123));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2125 (.A(net2125),
    .X(net2124));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2126 (.A(net2158),
    .X(net2125));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2127 (.A(net2128),
    .X(net2126));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2128 (.A(net2128),
    .X(net2127));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2129 (.A(net2158),
    .X(net2128));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2130 (.A(net2131),
    .X(net2129));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2131 (.A(net2131),
    .X(net2130));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2132 (.A(net2158),
    .X(net2131));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2133 (.A(net2140),
    .X(net2132));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2134 (.A(net2135),
    .X(net2133));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2135 (.A(net2135),
    .X(net2134));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2136 (.A(net2140),
    .X(net2135));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2137 (.A(net2137),
    .X(net2136));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2138 (.A(net2140),
    .X(net2137));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2139 (.A(net2139),
    .X(net2138));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2140 (.A(net2140),
    .X(net2139));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2141 (.A(net2158),
    .X(net2140));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2142 (.A(net2145),
    .X(net2141));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2143 (.A(net2145),
    .X(net2142));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2144 (.A(net2144),
    .X(net2143));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2145 (.A(net2145),
    .X(net2144));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2146 (.A(net2158),
    .X(net2145));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2147 (.A(net2149),
    .X(net2146));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2148 (.A(net2149),
    .X(net2147));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2149 (.A(net2149),
    .X(net2148));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2150 (.A(net2158),
    .X(net2149));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2151 (.A(net2153),
    .X(net2150));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2152 (.A(net2153),
    .X(net2151));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2153 (.A(net2153),
    .X(net2152));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2154 (.A(net2158),
    .X(net2153));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2155 (.A(net2155),
    .X(net2154));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2156 (.A(net2157),
    .X(net2155));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2157 (.A(net2157),
    .X(net2156));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2158 (.A(net2158),
    .X(net2157));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2159 (.A(net2189),
    .X(net2158));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2160 (.A(net2160),
    .X(net2159));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2161 (.A(net2163),
    .X(net2160));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2162 (.A(net2162),
    .X(net2161));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2163 (.A(net2163),
    .X(net2162));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2164 (.A(net2176),
    .X(net2163));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2165 (.A(net2165),
    .X(net2164));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2166 (.A(net2166),
    .X(net2165));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2167 (.A(net2170),
    .X(net2166));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2168 (.A(net2170),
    .X(net2167));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2169 (.A(net2170),
    .X(net2168));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2170 (.A(net2170),
    .X(net2169));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2171 (.A(net2176),
    .X(net2170));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2172 (.A(net2175),
    .X(net2171));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2173 (.A(net2174),
    .X(net2172));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2174 (.A(net2174),
    .X(net2173));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2175 (.A(net2175),
    .X(net2174));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2176 (.A(net2176),
    .X(net2175));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2177 (.A(net2189),
    .X(net2176));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2178 (.A(net2178),
    .X(net2177));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2179 (.A(net2187),
    .X(net2178));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2180 (.A(net2187),
    .X(net2179));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2181 (.A(net2187),
    .X(net2180));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2182 (.A(net2182),
    .X(net2181));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2183 (.A(net2183),
    .X(net2182));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2184 (.A(net2187),
    .X(net2183));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2185 (.A(net2185),
    .X(net2184));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2186 (.A(net2186),
    .X(net2185));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2187 (.A(net2187),
    .X(net2186));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2188 (.A(net2189),
    .X(net2187));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2189 (.A(_09401_),
    .X(net2188));
 sky130_fd_sc_hd__buf_12 wire2190 (.A(net2188),
    .X(net2189));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2191 (.A(_09184_),
    .X(net2190));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2192 (.A(_09184_),
    .X(net2191));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2193 (.A(_09184_),
    .X(net2192));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2194 (.A(_09184_),
    .X(net2193));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2195 (.A(net2195),
    .X(net2194));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2196 (.A(_05630_),
    .X(net2195));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2197 (.A(net2197),
    .X(net2196));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2198 (.A(_20422_),
    .X(net2197));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2199 (.A(net2200),
    .X(net2198));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2200 (.A(net2200),
    .X(net2199));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2201 (.A(_20422_),
    .X(net2200));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2202 (.A(net2204),
    .X(net2201));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2203 (.A(net2204),
    .X(net2202));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2204 (.A(net2204),
    .X(net2203));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2205 (.A(_20399_),
    .X(net2204));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2206 (.A(net2207),
    .X(net2205));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2207 (.A(net2207),
    .X(net2206));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2208 (.A(_20399_),
    .X(net2207));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2209 (.A(net2209),
    .X(net2208));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2210 (.A(_20386_),
    .X(net2209));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2211 (.A(_20386_),
    .X(net2210));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2212 (.A(net2213),
    .X(net2211));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2213 (.A(net2213),
    .X(net2212));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2214 (.A(_20383_),
    .X(net2213));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2215 (.A(net2215),
    .X(net2214));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2216 (.A(_20381_),
    .X(net2215));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2217 (.A(net2219),
    .X(net2216));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2218 (.A(net2219),
    .X(net2217));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2219 (.A(net2219),
    .X(net2218));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2220 (.A(net2236),
    .X(net2219));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2221 (.A(net2223),
    .X(net2220));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2222 (.A(net2222),
    .X(net2221));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2223 (.A(net2223),
    .X(net2222));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2224 (.A(net2236),
    .X(net2223));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2225 (.A(net2225),
    .X(net2224));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2226 (.A(net2236),
    .X(net2225));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2227 (.A(net2227),
    .X(net2226));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2228 (.A(net2235),
    .X(net2227));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2229 (.A(net2235),
    .X(net2228));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2230 (.A(net2235),
    .X(net2229));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2231 (.A(net2235),
    .X(net2230));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2232 (.A(net2235),
    .X(net2231));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2233 (.A(net2234),
    .X(net2232));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2234 (.A(net2234),
    .X(net2233));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2235 (.A(net2235),
    .X(net2234));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2236 (.A(net2236),
    .X(net2235));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2237 (.A(net2237),
    .X(net2236));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2238 (.A(net2250),
    .X(net2237));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2239 (.A(net2250),
    .X(net2238));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2240 (.A(net2249),
    .X(net2239));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2241 (.A(net2241),
    .X(net2240));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2242 (.A(net2249),
    .X(net2241));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2243 (.A(net2246),
    .X(net2242));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2244 (.A(net2245),
    .X(net2243));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2245 (.A(net2245),
    .X(net2244));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2246 (.A(net2246),
    .X(net2245));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2247 (.A(net2249),
    .X(net2246));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2248 (.A(net2249),
    .X(net2247));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2249 (.A(net2249),
    .X(net2248));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2250 (.A(net2250),
    .X(net2249));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2251 (.A(_20367_),
    .X(net2250));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2252 (.A(net2252),
    .X(net2251));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2253 (.A(net2259),
    .X(net2252));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2254 (.A(net2254),
    .X(net2253));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2255 (.A(net2259),
    .X(net2254));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2256 (.A(net2259),
    .X(net2255));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2257 (.A(net2258),
    .X(net2256));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2258 (.A(net2258),
    .X(net2257));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2259 (.A(net2259),
    .X(net2258));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2260 (.A(net2313),
    .X(net2259));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2261 (.A(net2261),
    .X(net2260));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2262 (.A(net2262),
    .X(net2261));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2263 (.A(net2264),
    .X(net2262));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2264 (.A(net2264),
    .X(net2263));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2265 (.A(net2313),
    .X(net2264));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2266 (.A(net2266),
    .X(net2265));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2267 (.A(net2267),
    .X(net2266));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2268 (.A(net2285),
    .X(net2267));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2269 (.A(net2269),
    .X(net2268));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2270 (.A(net2270),
    .X(net2269));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2271 (.A(net2285),
    .X(net2270));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2272 (.A(net2273),
    .X(net2271));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2273 (.A(net2273),
    .X(net2272));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2274 (.A(net2285),
    .X(net2273));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2275 (.A(net2275),
    .X(net2274));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2276 (.A(net2285),
    .X(net2275));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2277 (.A(net2277),
    .X(net2276));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2278 (.A(net2284),
    .X(net2277));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2279 (.A(net2281),
    .X(net2278));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2280 (.A(net2281),
    .X(net2279));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2281 (.A(net2281),
    .X(net2280));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2282 (.A(net2284),
    .X(net2281));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2283 (.A(net2283),
    .X(net2282));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2284 (.A(net2284),
    .X(net2283));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2285 (.A(net2285),
    .X(net2284));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2286 (.A(net2298),
    .X(net2285));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2287 (.A(net2288),
    .X(net2286));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2288 (.A(net2288),
    .X(net2287));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2289 (.A(net2298),
    .X(net2288));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2290 (.A(net2291),
    .X(net2289));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2291 (.A(net2291),
    .X(net2290));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2292 (.A(net2292),
    .X(net2291));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2293 (.A(net2294),
    .X(net2292));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2294 (.A(net2294),
    .X(net2293));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2295 (.A(net2298),
    .X(net2294));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2296 (.A(net2296),
    .X(net2295));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2297 (.A(net2297),
    .X(net2296));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2298 (.A(net2298),
    .X(net2297));
 sky130_fd_sc_hd__buf_2 fanout2299 (.A(net2312),
    .X(net2298));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2300 (.A(net2302),
    .X(net2299));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2301 (.A(net2302),
    .X(net2300));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2302 (.A(net2302),
    .X(net2301));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2303 (.A(net2312),
    .X(net2302));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2304 (.A(net2312),
    .X(net2303));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2305 (.A(net2311),
    .X(net2304));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2306 (.A(net2306),
    .X(net2305));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2307 (.A(net2308),
    .X(net2306));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2308 (.A(net2308),
    .X(net2307));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2309 (.A(net2311),
    .X(net2308));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2310 (.A(net2311),
    .X(net2309));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2311 (.A(net2311),
    .X(net2310));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2312 (.A(net2312),
    .X(net2311));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2313 (.A(_20367_),
    .X(net2312));
 sky130_fd_sc_hd__buf_6 wire2314 (.A(_20367_),
    .X(net2313));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2315 (.A(net2315),
    .X(net2314));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2316 (.A(net2318),
    .X(net2315));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2317 (.A(net2317),
    .X(net2316));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2318 (.A(net2318),
    .X(net2317));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2319 (.A(net2321),
    .X(net2318));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2320 (.A(net2320),
    .X(net2319));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2321 (.A(net2321),
    .X(net2320));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2322 (.A(_20333_),
    .X(net2321));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2323 (.A(_20333_),
    .X(net2322));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2324 (.A(net2325),
    .X(net2323));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2325 (.A(net2325),
    .X(net2324));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2326 (.A(net2328),
    .X(net2325));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2327 (.A(net2328),
    .X(net2326));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2328 (.A(net2328),
    .X(net2327));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2329 (.A(net2346),
    .X(net2328));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2330 (.A(net2333),
    .X(net2329));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2331 (.A(net2333),
    .X(net2330));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2332 (.A(net2333),
    .X(net2331));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2333 (.A(net2333),
    .X(net2332));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2334 (.A(net2346),
    .X(net2333));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2335 (.A(net2335),
    .X(net2334));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2336 (.A(net2339),
    .X(net2335));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2337 (.A(net2338),
    .X(net2336));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2338 (.A(net2338),
    .X(net2337));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2339 (.A(net2339),
    .X(net2338));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2340 (.A(net2346),
    .X(net2339));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2341 (.A(net2342),
    .X(net2340));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2342 (.A(net2342),
    .X(net2341));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2343 (.A(net2346),
    .X(net2342));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2344 (.A(net2345),
    .X(net2343));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2345 (.A(net2345),
    .X(net2344));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2346 (.A(net2346),
    .X(net2345));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2347 (.A(_20333_),
    .X(net2346));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2348 (.A(net2348),
    .X(net2347));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2349 (.A(net2349),
    .X(net2348));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2350 (.A(net2412),
    .X(net2349));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2351 (.A(net2351),
    .X(net2350));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2352 (.A(net2360),
    .X(net2351));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2353 (.A(net2360),
    .X(net2352));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2354 (.A(net2360),
    .X(net2353));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2355 (.A(net2360),
    .X(net2354));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2356 (.A(net2357),
    .X(net2355));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2357 (.A(net2357),
    .X(net2356));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2358 (.A(net2360),
    .X(net2357));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2359 (.A(net2360),
    .X(net2358));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2360 (.A(net2360),
    .X(net2359));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2361 (.A(net2412),
    .X(net2360));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2362 (.A(net2363),
    .X(net2361));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2363 (.A(net2363),
    .X(net2362));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2364 (.A(net2364),
    .X(net2363));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2365 (.A(net2412),
    .X(net2364));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2366 (.A(net2367),
    .X(net2365));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2367 (.A(net2367),
    .X(net2366));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2368 (.A(net2386),
    .X(net2367));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2369 (.A(net2370),
    .X(net2368));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2370 (.A(net2370),
    .X(net2369));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2371 (.A(net2386),
    .X(net2370));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2372 (.A(net2375),
    .X(net2371));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2373 (.A(net2375),
    .X(net2372));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2374 (.A(net2375),
    .X(net2373));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2375 (.A(net2375),
    .X(net2374));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2376 (.A(net2386),
    .X(net2375));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2377 (.A(net2380),
    .X(net2376));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2378 (.A(net2380),
    .X(net2377));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2379 (.A(net2380),
    .X(net2378));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2380 (.A(net2380),
    .X(net2379));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2381 (.A(net2386),
    .X(net2380));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2382 (.A(net2382),
    .X(net2381));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2383 (.A(net2386),
    .X(net2382));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2384 (.A(net2385),
    .X(net2383));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2385 (.A(net2385),
    .X(net2384));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2386 (.A(net2386),
    .X(net2385));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2387 (.A(net2412),
    .X(net2386));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2388 (.A(net2389),
    .X(net2387));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2389 (.A(net2389),
    .X(net2388));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2390 (.A(net2411),
    .X(net2389));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2391 (.A(net2391),
    .X(net2390));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2392 (.A(net2411),
    .X(net2391));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2393 (.A(net2394),
    .X(net2392));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2394 (.A(net2394),
    .X(net2393));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2395 (.A(net2411),
    .X(net2394));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2396 (.A(net2397),
    .X(net2395));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2397 (.A(net2397),
    .X(net2396));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2398 (.A(net2411),
    .X(net2397));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2399 (.A(net2399),
    .X(net2398));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2400 (.A(net2403),
    .X(net2399));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2401 (.A(net2402),
    .X(net2400));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2402 (.A(net2402),
    .X(net2401));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2403 (.A(net2403),
    .X(net2402));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2404 (.A(net2411),
    .X(net2403));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2405 (.A(net2407),
    .X(net2404));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2406 (.A(net2407),
    .X(net2405));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2407 (.A(net2407),
    .X(net2406));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2408 (.A(net2411),
    .X(net2407));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2409 (.A(net2410),
    .X(net2408));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2410 (.A(net2410),
    .X(net2409));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2411 (.A(net2411),
    .X(net2410));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2412 (.A(net2412),
    .X(net2411));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2413 (.A(_20327_),
    .X(net2412));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2414 (.A(net2414),
    .X(net2413));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2415 (.A(net2416),
    .X(net2414));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2416 (.A(net2416),
    .X(net2415));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2417 (.A(net2417),
    .X(net2416));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2418 (.A(_20324_),
    .X(net2417));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2419 (.A(net2420),
    .X(net2418));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2420 (.A(net2420),
    .X(net2419));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2421 (.A(net2429),
    .X(net2420));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2422 (.A(net2429),
    .X(net2421));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2423 (.A(net2429),
    .X(net2422));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2424 (.A(net2425),
    .X(net2423));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2425 (.A(net2425),
    .X(net2424));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2426 (.A(net2429),
    .X(net2425));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2427 (.A(net2428),
    .X(net2426));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2428 (.A(net2428),
    .X(net2427));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2429 (.A(net2429),
    .X(net2428));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2430 (.A(_20324_),
    .X(net2429));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2431 (.A(net2431),
    .X(net2430));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2432 (.A(net2432),
    .X(net2431));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2433 (.A(_20320_),
    .X(net2432));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2434 (.A(net2441),
    .X(net2433));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2435 (.A(net2441),
    .X(net2434));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2436 (.A(net2441),
    .X(net2435));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2437 (.A(net2441),
    .X(net2436));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2438 (.A(net2441),
    .X(net2437));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2439 (.A(net2441),
    .X(net2438));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2440 (.A(net2441),
    .X(net2439));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2441 (.A(net2441),
    .X(net2440));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2442 (.A(_20320_),
    .X(net2441));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2443 (.A(net2444),
    .X(net2442));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2444 (.A(net2444),
    .X(net2443));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2445 (.A(_20318_),
    .X(net2444));
 sky130_fd_sc_hd__buf_12 wire2446 (.A(net2444),
    .X(net2445));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2447 (.A(net2449),
    .X(net2446));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2448 (.A(net2449),
    .X(net2447));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2449 (.A(net2449),
    .X(net2448));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2450 (.A(net2450),
    .X(net2449));
 sky130_fd_sc_hd__buf_2 fanout2451 (.A(_20272_),
    .X(net2450));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2452 (.A(net2452),
    .X(net2451));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2453 (.A(net2460),
    .X(net2452));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2454 (.A(net2455),
    .X(net2453));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2455 (.A(net2455),
    .X(net2454));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2456 (.A(net2460),
    .X(net2455));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2457 (.A(net2459),
    .X(net2456));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2458 (.A(net2459),
    .X(net2457));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2459 (.A(net2459),
    .X(net2458));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2460 (.A(net2460),
    .X(net2459));
 sky130_fd_sc_hd__buf_2 fanout2461 (.A(_20264_),
    .X(net2460));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2462 (.A(net2462),
    .X(net2461));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2463 (.A(net2463),
    .X(net2462));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2464 (.A(net2464),
    .X(net2463));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2465 (.A(net2465),
    .X(net2464));
 sky130_fd_sc_hd__buf_2 fanout2466 (.A(_20263_),
    .X(net2465));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2467 (.A(net2469),
    .X(net2466));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2468 (.A(net2469),
    .X(net2467));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2469 (.A(net2469),
    .X(net2468));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2470 (.A(net2495),
    .X(net2469));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2471 (.A(net2472),
    .X(net2470));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2472 (.A(net2472),
    .X(net2471));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2473 (.A(net2495),
    .X(net2472));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2474 (.A(net2474),
    .X(net2473));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2475 (.A(net2478),
    .X(net2474));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2476 (.A(net2478),
    .X(net2475));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2477 (.A(net2478),
    .X(net2476));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2478 (.A(net2478),
    .X(net2477));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2479 (.A(net2495),
    .X(net2478));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2480 (.A(net2482),
    .X(net2479));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2481 (.A(net2482),
    .X(net2480));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2482 (.A(net2482),
    .X(net2481));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2483 (.A(net2495),
    .X(net2482));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2484 (.A(net2486),
    .X(net2483));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2485 (.A(net2486),
    .X(net2484));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2486 (.A(net2486),
    .X(net2485));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2487 (.A(net2495),
    .X(net2486));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2488 (.A(net2489),
    .X(net2487));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2489 (.A(net2489),
    .X(net2488));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2490 (.A(net2494),
    .X(net2489));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2491 (.A(net2494),
    .X(net2490));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2492 (.A(net2494),
    .X(net2491));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2493 (.A(net2494),
    .X(net2492));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2494 (.A(net2494),
    .X(net2493));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2495 (.A(net2495),
    .X(net2494));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2496 (.A(_20263_),
    .X(net2495));
 sky130_fd_sc_hd__buf_2 fanout2497 (.A(net2504),
    .X(net2496));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2498 (.A(net2504),
    .X(net2497));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2499 (.A(net2504),
    .X(net2498));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2500 (.A(net2504),
    .X(net2499));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2501 (.A(net2503),
    .X(net2500));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2502 (.A(net2503),
    .X(net2501));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2503 (.A(net2503),
    .X(net2502));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2504 (.A(net2504),
    .X(net2503));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2505 (.A(_20237_),
    .X(net2504));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2506 (.A(net2508),
    .X(net2505));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2507 (.A(net2508),
    .X(net2506));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2508 (.A(net2508),
    .X(net2507));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2509 (.A(net2509),
    .X(net2508));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2510 (.A(_20235_),
    .X(net2509));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2511 (.A(net2511),
    .X(net2510));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2512 (.A(net2517),
    .X(net2511));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2513 (.A(net2517),
    .X(net2512));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2514 (.A(net2517),
    .X(net2513));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2515 (.A(net2517),
    .X(net2514));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2516 (.A(net2517),
    .X(net2515));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2517 (.A(net2517),
    .X(net2516));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2518 (.A(_20235_),
    .X(net2517));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2519 (.A(net2519),
    .X(net2518));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2520 (.A(net2526),
    .X(net2519));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2521 (.A(net2526),
    .X(net2520));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2522 (.A(net2526),
    .X(net2521));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2523 (.A(net2523),
    .X(net2522));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2524 (.A(net2526),
    .X(net2523));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2525 (.A(net2526),
    .X(net2524));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2526 (.A(net2526),
    .X(net2525));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2527 (.A(_20235_),
    .X(net2526));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2528 (.A(net2536),
    .X(net2527));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2529 (.A(net2536),
    .X(net2528));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2530 (.A(net2530),
    .X(net2529));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2531 (.A(net2536),
    .X(net2530));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2532 (.A(net2532),
    .X(net2531));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2533 (.A(net2535),
    .X(net2532));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2534 (.A(net2535),
    .X(net2533));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2535 (.A(net2535),
    .X(net2534));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2536 (.A(net2536),
    .X(net2535));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2537 (.A(_20235_),
    .X(net2536));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2538 (.A(net2540),
    .X(net2537));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2539 (.A(net2539),
    .X(net2538));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2540 (.A(net2540),
    .X(net2539));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2541 (.A(net2545),
    .X(net2540));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2542 (.A(net2545),
    .X(net2541));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2543 (.A(net2543),
    .X(net2542));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2544 (.A(net2544),
    .X(net2543));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2545 (.A(net2545),
    .X(net2544));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2546 (.A(_20223_),
    .X(net2545));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2547 (.A(net2550),
    .X(net2546));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2548 (.A(net2550),
    .X(net2547));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2549 (.A(net2550),
    .X(net2548));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2550 (.A(net2550),
    .X(net2549));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2551 (.A(_19902_),
    .X(net2550));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2552 (.A(net2552),
    .X(net2551));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2553 (.A(net2554),
    .X(net2552));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2554 (.A(net2554),
    .X(net2553));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2555 (.A(_19889_),
    .X(net2554));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2556 (.A(net2556),
    .X(net2555));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2557 (.A(net2557),
    .X(net2556));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2558 (.A(_19847_),
    .X(net2557));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2559 (.A(net2560),
    .X(net2558));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2560 (.A(net2560),
    .X(net2559));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2561 (.A(\inst$top.soc.wb_arbiter.grant ),
    .X(net2560));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2562 (.A(net2566),
    .X(net2561));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2563 (.A(net2565),
    .X(net2562));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2564 (.A(net2565),
    .X(net2563));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2565 (.A(net2565),
    .X(net2564));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2566 (.A(net2566),
    .X(net2565));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2567 (.A(\inst$top.soc.wb_arbiter.grant ),
    .X(net2566));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2568 (.A(\inst$top.soc.uart_0._phy.tx.lower.fsm_state ),
    .X(net2567));
 sky130_fd_sc_hd__buf_16 wire2569 (.A(net582),
    .X(net2568));
 sky130_fd_sc_hd__buf_16 wire2570 (.A(net563),
    .X(net2569));
 sky130_fd_sc_hd__buf_16 wire2571 (.A(net597),
    .X(net2570));
 sky130_fd_sc_hd__buf_16 wire2572 (.A(net562),
    .X(net2571));
 sky130_fd_sc_hd__buf_16 wire2573 (.A(net596),
    .X(net2572));
 sky130_fd_sc_hd__buf_16 wire2574 (.A(net561),
    .X(net2573));
 sky130_fd_sc_hd__buf_16 wire2575 (.A(net595),
    .X(net2574));
 sky130_fd_sc_hd__buf_16 wire2576 (.A(net560),
    .X(net2575));
 sky130_fd_sc_hd__buf_16 wire2577 (.A(net594),
    .X(net2576));
 sky130_fd_sc_hd__buf_16 wire2578 (.A(\inst$top.soc.spiflash.phy.io_streamer.buffer_cs.o_ff ),
    .X(net2577));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2579 (.A(\inst$top.soc.spiflash.phy.enframer.cycle[1] ),
    .X(net2578));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2580 (.A(\inst$top.soc.spiflash.phy.enframer.cycle[0] ),
    .X(net2579));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2581 (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb$17 ),
    .X(net2580));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2582 (.A(\inst$top.soc.spiflash.ctrl.csr_bridge.mux.element__w_stb$17 ),
    .X(net2581));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2583 (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb ),
    .X(net2582));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2584 (.A(\inst$top.soc.gpio_open_drain._gpio.bridge.mux.element__w_stb ),
    .X(net2583));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2585 (.A(net2585),
    .X(net2584));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2586 (.A(net2586),
    .X(net2585));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2587 (.A(\inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb ),
    .X(net2586));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2588 (.A(\inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb$21 ),
    .X(net2587));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2589 (.A(\inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb$20 ),
    .X(net2588));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2590 (.A(\inst$top.soc.gpio_0._gpio.bridge.mux.element__w_stb$20 ),
    .X(net2589));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2591 (.A(net2595),
    .X(net2590));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2592 (.A(net2595),
    .X(net2591));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2593 (.A(net2596),
    .X(net2592));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2594 (.A(net2594),
    .X(net2593));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2595 (.A(net2596),
    .X(net2594));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2596 (.A(\inst$top.soc.cpu.sink__payload$6[56] ),
    .X(net2595));
 sky130_fd_sc_hd__buf_16 wire2597 (.A(net2595),
    .X(net2596));
 sky130_fd_sc_hd__buf_2 fanout2598 (.A(net2606),
    .X(net2597));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2599 (.A(net2600),
    .X(net2598));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2600 (.A(net2600),
    .X(net2599));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2601 (.A(net2606),
    .X(net2600));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2602 (.A(net2605),
    .X(net2601));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2603 (.A(net2605),
    .X(net2602));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2604 (.A(net2604),
    .X(net2603));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2605 (.A(net2605),
    .X(net2604));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2606 (.A(net2606),
    .X(net2605));
 sky130_fd_sc_hd__buf_2 fanout2607 (.A(\inst$top.soc.cpu.sink__payload$6[55] ),
    .X(net2606));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2608 (.A(net2608),
    .X(net2607));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2609 (.A(\inst$top.soc.cpu.sink__payload$6[54] ),
    .X(net2608));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2610 (.A(net2615),
    .X(net2609));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2611 (.A(net2615),
    .X(net2610));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2612 (.A(net2614),
    .X(net2611));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2613 (.A(net2614),
    .X(net2612));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2614 (.A(net2614),
    .X(net2613));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2615 (.A(net2615),
    .X(net2614));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2616 (.A(\inst$top.soc.cpu.sink__payload$6[54] ),
    .X(net2615));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2617 (.A(net2617),
    .X(net2616));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2618 (.A(net2618),
    .X(net2617));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2619 (.A(net2619),
    .X(net2618));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2620 (.A(net2620),
    .X(net2619));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2621 (.A(\inst$top.soc.cpu.sink__payload$6[53] ),
    .X(net2620));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2622 (.A(net2623),
    .X(net2621));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2623 (.A(net2623),
    .X(net2622));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2624 (.A(net2651),
    .X(net2623));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2625 (.A(net2626),
    .X(net2624));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2626 (.A(net2626),
    .X(net2625));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2627 (.A(net2651),
    .X(net2626));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2628 (.A(net2628),
    .X(net2627));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2629 (.A(net2632),
    .X(net2628));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2630 (.A(net2632),
    .X(net2629));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2631 (.A(net2632),
    .X(net2630));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2632 (.A(net2632),
    .X(net2631));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2633 (.A(net2651),
    .X(net2632));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2634 (.A(net2636),
    .X(net2633));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2635 (.A(net2636),
    .X(net2634));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2636 (.A(net2636),
    .X(net2635));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2637 (.A(net2641),
    .X(net2636));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2638 (.A(net2641),
    .X(net2637));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2639 (.A(net2641),
    .X(net2638));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2640 (.A(net2641),
    .X(net2639));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2641 (.A(net2641),
    .X(net2640));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2642 (.A(net2651),
    .X(net2641));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2643 (.A(net2645),
    .X(net2642));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2644 (.A(net2645),
    .X(net2643));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2645 (.A(net2645),
    .X(net2644));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2646 (.A(net2650),
    .X(net2645));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2647 (.A(net2650),
    .X(net2646));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2648 (.A(net2650),
    .X(net2647));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2649 (.A(net2650),
    .X(net2648));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2650 (.A(net2650),
    .X(net2649));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2651 (.A(net2651),
    .X(net2650));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2652 (.A(\inst$top.soc.cpu.sink__payload$6[53] ),
    .X(net2651));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2653 (.A(net2655),
    .X(net2652));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2654 (.A(net2655),
    .X(net2653));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2655 (.A(net2655),
    .X(net2654));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2656 (.A(net2656),
    .X(net2655));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2657 (.A(net2688),
    .X(net2656));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2658 (.A(net2665),
    .X(net2657));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2659 (.A(net2665),
    .X(net2658));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2660 (.A(net2665),
    .X(net2659));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2661 (.A(net2665),
    .X(net2660));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2662 (.A(net2664),
    .X(net2661));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2663 (.A(net2664),
    .X(net2662));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2664 (.A(net2664),
    .X(net2663));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2665 (.A(net2665),
    .X(net2664));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2666 (.A(net2688),
    .X(net2665));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2667 (.A(net2674),
    .X(net2666));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2668 (.A(net2674),
    .X(net2667));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2669 (.A(net2674),
    .X(net2668));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2670 (.A(net2674),
    .X(net2669));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2671 (.A(net2671),
    .X(net2670));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2672 (.A(net2674),
    .X(net2671));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2673 (.A(net2674),
    .X(net2672));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2674 (.A(net2674),
    .X(net2673));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2675 (.A(net2688),
    .X(net2674));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2676 (.A(net2685),
    .X(net2675));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2677 (.A(net2685),
    .X(net2676));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2678 (.A(net2678),
    .X(net2677));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2679 (.A(net2685),
    .X(net2678));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2680 (.A(net2685),
    .X(net2679));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2681 (.A(net2685),
    .X(net2680));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2682 (.A(net2685),
    .X(net2681));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2683 (.A(net2684),
    .X(net2682));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2684 (.A(net2684),
    .X(net2683));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2685 (.A(net2685),
    .X(net2684));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2686 (.A(net2688),
    .X(net2685));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2687 (.A(\inst$top.soc.cpu.sink__payload$6[52] ),
    .X(net2686));
 sky130_fd_sc_hd__buf_16 wire2688 (.A(net2686),
    .X(net2687));
 sky130_fd_sc_hd__buf_16 wire2689 (.A(\inst$top.soc.cpu.sink__payload$6[52] ),
    .X(net2688));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2690 (.A(net2690),
    .X(net2689));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2691 (.A(\inst$top.soc.cpu.sink__payload$6[51] ),
    .X(net2690));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2692 (.A(net2693),
    .X(net2691));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2693 (.A(net2693),
    .X(net2692));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2694 (.A(\inst$top.soc.cpu.sink__payload$6[51] ),
    .X(net2693));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2695 (.A(\inst$top.soc.cpu.sink__payload$6[51] ),
    .X(net2694));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2696 (.A(net2696),
    .X(net2695));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2697 (.A(\inst$top.soc.cpu.sink__payload$6[50] ),
    .X(net2696));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2698 (.A(net2699),
    .X(net2697));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2699 (.A(net2699),
    .X(net2698));
 sky130_fd_sc_hd__buf_2 fanout2700 (.A(\inst$top.soc.cpu.sink__payload$6[50] ),
    .X(net2699));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2701 (.A(net2701),
    .X(net2700));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2702 (.A(net2702),
    .X(net2701));
 sky130_fd_sc_hd__buf_2 fanout2703 (.A(net2703),
    .X(net2702));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2704 (.A(\inst$top.soc.cpu.sink__payload$6[49] ),
    .X(net2703));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2705 (.A(net2706),
    .X(net2704));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2706 (.A(net2706),
    .X(net2705));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2707 (.A(net2709),
    .X(net2706));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2708 (.A(net2709),
    .X(net2707));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2709 (.A(net2709),
    .X(net2708));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2710 (.A(\inst$top.soc.cpu.sink__payload$6[49] ),
    .X(net2709));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2711 (.A(net2712),
    .X(net2710));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2712 (.A(net2712),
    .X(net2711));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2713 (.A(net2716),
    .X(net2712));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2714 (.A(net2716),
    .X(net2713));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2715 (.A(net2716),
    .X(net2714));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2716 (.A(net2716),
    .X(net2715));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2717 (.A(\inst$top.soc.cpu.sink__payload$6[49] ),
    .X(net2716));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2718 (.A(net2718),
    .X(net2717));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2719 (.A(net2721),
    .X(net2718));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2720 (.A(net2721),
    .X(net2719));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2721 (.A(net2721),
    .X(net2720));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2722 (.A(\inst$top.soc.cpu.sink__payload$6[48] ),
    .X(net2721));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2723 (.A(net2723),
    .X(net2722));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2724 (.A(net2724),
    .X(net2723));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2725 (.A(\inst$top.soc.cpu.sink__payload$6[48] ),
    .X(net2724));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2726 (.A(net2727),
    .X(net2725));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2727 (.A(net2727),
    .X(net2726));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2728 (.A(net2750),
    .X(net2727));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2729 (.A(net2730),
    .X(net2728));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2730 (.A(net2730),
    .X(net2729));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2731 (.A(net2750),
    .X(net2730));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2732 (.A(net2733),
    .X(net2731));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2733 (.A(net2733),
    .X(net2732));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2734 (.A(net2736),
    .X(net2733));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2735 (.A(net2735),
    .X(net2734));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2736 (.A(net2736),
    .X(net2735));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2737 (.A(net2750),
    .X(net2736));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2738 (.A(net2739),
    .X(net2737));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2739 (.A(net2739),
    .X(net2738));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2740 (.A(net2750),
    .X(net2739));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2741 (.A(net2742),
    .X(net2740));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2742 (.A(net2742),
    .X(net2741));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2743 (.A(net2750),
    .X(net2742));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2744 (.A(net2745),
    .X(net2743));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2745 (.A(net2745),
    .X(net2744));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2746 (.A(net2750),
    .X(net2745));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2747 (.A(net2749),
    .X(net2746));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2748 (.A(net2749),
    .X(net2747));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2749 (.A(net2749),
    .X(net2748));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2750 (.A(net2750),
    .X(net2749));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2751 (.A(\inst$top.soc.cpu.sink__payload$6[48] ),
    .X(net2750));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2752 (.A(net2756),
    .X(net2751));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2753 (.A(net2756),
    .X(net2752));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2754 (.A(net2756),
    .X(net2753));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2755 (.A(net2756),
    .X(net2754));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2756 (.A(net2756),
    .X(net2755));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2757 (.A(net2762),
    .X(net2756));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2758 (.A(net2759),
    .X(net2757));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2759 (.A(net2759),
    .X(net2758));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2760 (.A(net2762),
    .X(net2759));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2761 (.A(net2761),
    .X(net2760));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2762 (.A(net2762),
    .X(net2761));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2763 (.A(net2819),
    .X(net2762));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2764 (.A(net2765),
    .X(net2763));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2765 (.A(net2765),
    .X(net2764));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2766 (.A(net2766),
    .X(net2765));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2767 (.A(net2819),
    .X(net2766));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2768 (.A(net2819),
    .X(net2767));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2769 (.A(net2770),
    .X(net2768));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2770 (.A(net2770),
    .X(net2769));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2771 (.A(net2791),
    .X(net2770));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2772 (.A(net2773),
    .X(net2771));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2773 (.A(net2773),
    .X(net2772));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2774 (.A(net2791),
    .X(net2773));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2775 (.A(net2776),
    .X(net2774));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2776 (.A(net2776),
    .X(net2775));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2777 (.A(net2791),
    .X(net2776));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2778 (.A(net2779),
    .X(net2777));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2779 (.A(net2779),
    .X(net2778));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2780 (.A(net2791),
    .X(net2779));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2781 (.A(net2781),
    .X(net2780));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2782 (.A(net2784),
    .X(net2781));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2783 (.A(net2784),
    .X(net2782));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2784 (.A(net2784),
    .X(net2783));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2785 (.A(net2791),
    .X(net2784));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2786 (.A(net2786),
    .X(net2785));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2787 (.A(net2790),
    .X(net2786));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2788 (.A(net2790),
    .X(net2787));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2789 (.A(net2790),
    .X(net2788));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2790 (.A(net2790),
    .X(net2789));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2791 (.A(net2791),
    .X(net2790));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2792 (.A(net2819),
    .X(net2791));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2793 (.A(net2794),
    .X(net2792));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2794 (.A(net2794),
    .X(net2793));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2795 (.A(net2804),
    .X(net2794));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2796 (.A(net2796),
    .X(net2795));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2797 (.A(net2804),
    .X(net2796));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2798 (.A(net2800),
    .X(net2797));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2799 (.A(net2800),
    .X(net2798));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2800 (.A(net2800),
    .X(net2799));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2801 (.A(net2804),
    .X(net2800));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2802 (.A(net2803),
    .X(net2801));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2803 (.A(net2803),
    .X(net2802));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2804 (.A(net2804),
    .X(net2803));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2805 (.A(net2818),
    .X(net2804));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2806 (.A(net2807),
    .X(net2805));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2807 (.A(net2807),
    .X(net2806));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2808 (.A(net2818),
    .X(net2807));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2809 (.A(net2810),
    .X(net2808));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2810 (.A(net2810),
    .X(net2809));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2811 (.A(net2818),
    .X(net2810));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2812 (.A(net2814),
    .X(net2811));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2813 (.A(net2814),
    .X(net2812));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2814 (.A(net2814),
    .X(net2813));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2815 (.A(net2818),
    .X(net2814));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2816 (.A(net2817),
    .X(net2815));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2817 (.A(net2817),
    .X(net2816));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2818 (.A(net2818),
    .X(net2817));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2819 (.A(net2819),
    .X(net2818));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2820 (.A(\inst$top.soc.cpu.sink__payload$6[47] ),
    .X(net2819));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2821 (.A(\inst$top.soc.cpu.csr_fmt_i ),
    .X(net2820));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2822 (.A(\inst$top.soc.cpu.sink__payload$6[38] ),
    .X(net2821));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2823 (.A(net2824),
    .X(net2822));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2824 (.A(net2824),
    .X(net2823));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2825 (.A(\inst$top.soc.cpu.sink__payload$24[42] ),
    .X(net2824));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2826 (.A(\inst$top.soc.cpu.d.sink__payload$16.multiply ),
    .X(net2825));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2827 (.A(\inst$top.soc.cpu.d.sink__payload$16.multiply ),
    .X(net2826));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2828 (.A(\inst$top.soc.cpu.d.sink__payload$16.multiply ),
    .X(net2827));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2829 (.A(\inst$top.soc.cpu.d.sink__payload$16.multiply ),
    .X(net2828));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2830 (.A(net2832),
    .X(net2829));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2831 (.A(net2832),
    .X(net2830));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2832 (.A(net2832),
    .X(net2831));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2833 (.A(\inst$top.soc.cpu.d.sink__payload$6.compare ),
    .X(net2832));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2834 (.A(net2834),
    .X(net2833));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2835 (.A(net2841),
    .X(net2834));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2836 (.A(net2836),
    .X(net2835));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2837 (.A(net2841),
    .X(net2836));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2838 (.A(net2838),
    .X(net2837));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2839 (.A(net2839),
    .X(net2838));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2840 (.A(net2840),
    .X(net2839));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2841 (.A(net2841),
    .X(net2840));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2842 (.A(\inst$top.soc.cpu.d.sink__payload$6.shift ),
    .X(net2841));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2843 (.A(\inst$top.soc.cpu.d.sink__payload.csr_fmt_i ),
    .X(net2842));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2844 (.A(net2844),
    .X(net2843));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2845 (.A(net2845),
    .X(net2844));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2846 (.A(net2846),
    .X(net2845));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2847 (.A(net2850),
    .X(net2846));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2848 (.A(net2850),
    .X(net2847));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2849 (.A(net2849),
    .X(net2848));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2850 (.A(net2850),
    .X(net2849));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2851 (.A(\inst$top.soc.cpu.d.sink__payload.csr_re ),
    .X(net2850));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2852 (.A(net2853),
    .X(net2851));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2853 (.A(net2853),
    .X(net2852));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2854 (.A(\inst$top.soc.cpu.d.sink__payload.jump ),
    .X(net2853));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2855 (.A(net2856),
    .X(net2854));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2856 (.A(net2856),
    .X(net2855));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2857 (.A(\inst$top.soc.cpu.d.sink__payload.jump ),
    .X(net2856));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2858 (.A(net2860),
    .X(net2857));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2859 (.A(net2860),
    .X(net2858));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2860 (.A(net2860),
    .X(net2859));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2861 (.A(\inst$top.soc.cpu.d.sink__payload.direction ),
    .X(net2860));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2862 (.A(net2864),
    .X(net2861));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2863 (.A(net2863),
    .X(net2862));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2864 (.A(net2864),
    .X(net2863));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2865 (.A(\inst$top.soc.cpu.d.sink__payload.logic ),
    .X(net2864));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2866 (.A(net2868),
    .X(net2865));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2867 (.A(net2868),
    .X(net2866));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2868 (.A(net2868),
    .X(net2867));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2869 (.A(\inst$top.soc.cpu.adder$307.x_sub ),
    .X(net2868));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2870 (.A(net2870),
    .X(net2869));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2871 (.A(net2873),
    .X(net2870));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2872 (.A(net2873),
    .X(net2871));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2873 (.A(net2873),
    .X(net2872));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2874 (.A(\inst$top.soc.cpu.shifter.m_direction ),
    .X(net2873));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2875 (.A(net2881),
    .X(net2874));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2876 (.A(net2876),
    .X(net2875));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2877 (.A(net2881),
    .X(net2876));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2878 (.A(net2880),
    .X(net2877));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2879 (.A(net2879),
    .X(net2878));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2880 (.A(net2880),
    .X(net2879));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2881 (.A(net2881),
    .X(net2880));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2882 (.A(\inst$top.soc.cpu.multiplier.m_low ),
    .X(net2881));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2883 (.A(net2883),
    .X(net2882));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2884 (.A(\inst$top.soc.cpu.gprf.x_bypass2_raw ),
    .X(net2883));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2885 (.A(net2885),
    .X(net2884));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2886 (.A(\inst$top.soc.cpu.gprf.x_bypass2_raw ),
    .X(net2885));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2887 (.A(net2889),
    .X(net2886));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2888 (.A(net2889),
    .X(net2887));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2889 (.A(net2889),
    .X(net2888));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2890 (.A(\inst$top.soc.cpu.gprf.x_bypass1_raw ),
    .X(net2889));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2891 (.A(\inst$top.soc.cpu.exception.m_mstatus.mie ),
    .X(net2890));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2892 (.A(\inst$top.soc.cpu.exception.m_mstatus.mie ),
    .X(net2891));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2893 (.A(\inst$top.soc.cpu.exception.csr_bank.mtvec_x_select ),
    .X(net2892));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2894 (.A(net2896),
    .X(net2893));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2895 (.A(net2895),
    .X(net2894));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2896 (.A(net2896),
    .X(net2895));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2897 (.A(\inst$top.soc.cpu.exception.csr_bank.mtval_x_select ),
    .X(net2896));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2898 (.A(net2900),
    .X(net2897));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2899 (.A(net2900),
    .X(net2898));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2900 (.A(net2900),
    .X(net2899));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2901 (.A(\inst$top.soc.cpu.exception.csr_bank.mscratch_x_select ),
    .X(net2900));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2902 (.A(net2904),
    .X(net2901));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2903 (.A(net2903),
    .X(net2902));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2904 (.A(net2904),
    .X(net2903));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2905 (.A(\inst$top.soc.cpu.exception.csr_bank.mscratch_w_select ),
    .X(net2904));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2906 (.A(\inst$top.soc.cpu.exception.csr_bank.mip_x_select ),
    .X(net2905));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2907 (.A(\inst$top.soc.cpu.exception.csr_bank.mip_w_select ),
    .X(net2906));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2908 (.A(\inst$top.soc.cpu.exception.csr_bank.mip_w_select ),
    .X(net2907));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2909 (.A(net2911),
    .X(net2908));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2910 (.A(net2910),
    .X(net2909));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2911 (.A(net2911),
    .X(net2910));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2912 (.A(\inst$top.soc.cpu.exception.csr_bank.mepc_x_select ),
    .X(net2911));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2913 (.A(net2915),
    .X(net2912));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2914 (.A(net2914),
    .X(net2913));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2915 (.A(net2915),
    .X(net2914));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2916 (.A(\inst$top.soc.cpu.exception.csr_bank.mcause_x_select ),
    .X(net2915));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2917 (.A(net2917),
    .X(net2916));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2918 (.A(net2918),
    .X(net2917));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2919 (.A(net2920),
    .X(net2918));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2920 (.A(net2920),
    .X(net2919));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2921 (.A(\inst$top.soc.cpu.divider.m_modulus ),
    .X(net2920));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2922 (.A(net2924),
    .X(net2921));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2923 (.A(net2924),
    .X(net2922));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2924 (.A(net2924),
    .X(net2923));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2925 (.A(\inst$top.soc.cpu.divider.m_modulus ),
    .X(net2924));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2926 (.A(net2927),
    .X(net2925));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2927 (.A(net2927),
    .X(net2926));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2928 (.A(net2931),
    .X(net2927));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2929 (.A(net2930),
    .X(net2928));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2930 (.A(net2930),
    .X(net2929));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2931 (.A(net2931),
    .X(net2930));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2932 (.A(\inst$top.soc.cpu.divider.fsm_state ),
    .X(net2931));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2933 (.A(net2934),
    .X(net2932));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2934 (.A(net2934),
    .X(net2933));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2935 (.A(net2935),
    .X(net2934));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2936 (.A(net2956),
    .X(net2935));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2937 (.A(net2937),
    .X(net2936));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2938 (.A(net2938),
    .X(net2937));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2939 (.A(net2956),
    .X(net2938));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2940 (.A(net2942),
    .X(net2939));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2941 (.A(net2942),
    .X(net2940));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2942 (.A(net2942),
    .X(net2941));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2943 (.A(net2943),
    .X(net2942));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2944 (.A(net2956),
    .X(net2943));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2945 (.A(net2945),
    .X(net2944));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2946 (.A(net2956),
    .X(net2945));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2947 (.A(net2947),
    .X(net2946));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2948 (.A(net2956),
    .X(net2947));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2949 (.A(net2951),
    .X(net2948));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2950 (.A(net2951),
    .X(net2949));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2951 (.A(net2951),
    .X(net2950));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2952 (.A(net2956),
    .X(net2951));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2953 (.A(net2953),
    .X(net2952));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2954 (.A(net2954),
    .X(net2953));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2955 (.A(net2955),
    .X(net2954));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2956 (.A(net2956),
    .X(net2955));
 sky130_fd_sc_hd__buf_2 fanout2957 (.A(\inst$top.rst_n_sync.rst ),
    .X(net2956));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2958 (.A(net2960),
    .X(net2957));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2959 (.A(net2960),
    .X(net2958));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2960 (.A(net2960),
    .X(net2959));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2961 (.A(net2966),
    .X(net2960));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2962 (.A(net2963),
    .X(net2961));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2963 (.A(net2963),
    .X(net2962));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2964 (.A(net2966),
    .X(net2963));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2965 (.A(net2965),
    .X(net2964));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2966 (.A(net2966),
    .X(net2965));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2967 (.A(net2978),
    .X(net2966));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2968 (.A(net2978),
    .X(net2967));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2969 (.A(net2970),
    .X(net2968));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2970 (.A(net2970),
    .X(net2969));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2971 (.A(net2973),
    .X(net2970));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2972 (.A(net2972),
    .X(net2971));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2973 (.A(net2973),
    .X(net2972));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2974 (.A(net2978),
    .X(net2973));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2975 (.A(net2975),
    .X(net2974));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2976 (.A(net2976),
    .X(net2975));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2977 (.A(net2977),
    .X(net2976));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2978 (.A(net2978),
    .X(net2977));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2979 (.A(\inst$top.rst_n_sync.rst ),
    .X(net2978));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2980 (.A(net2983),
    .X(net2979));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2981 (.A(net2981),
    .X(net2980));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2982 (.A(net2982),
    .X(net2981));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2983 (.A(net2983),
    .X(net2982));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2984 (.A(net2994),
    .X(net2983));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2985 (.A(net2985),
    .X(net2984));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2986 (.A(net2992),
    .X(net2985));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2987 (.A(net2987),
    .X(net2986));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2988 (.A(net2992),
    .X(net2987));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2989 (.A(net2991),
    .X(net2988));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2990 (.A(net2991),
    .X(net2989));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2991 (.A(net2991),
    .X(net2990));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2992 (.A(net2992),
    .X(net2991));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2993 (.A(net2994),
    .X(net2992));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2994 (.A(net2994),
    .X(net2993));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2995 (.A(net3004),
    .X(net2994));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2996 (.A(net2998),
    .X(net2995));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2997 (.A(net2998),
    .X(net2996));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2998 (.A(net2998),
    .X(net2997));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout2999 (.A(net3003),
    .X(net2998));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3000 (.A(net3000),
    .X(net2999));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3001 (.A(net3003),
    .X(net3000));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3002 (.A(net3002),
    .X(net3001));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3003 (.A(net3003),
    .X(net3002));
 sky130_fd_sc_hd__buf_2 fanout3004 (.A(net3004),
    .X(net3003));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3005 (.A(net3015),
    .X(net3004));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3006 (.A(net3014),
    .X(net3005));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3007 (.A(net3014),
    .X(net3006));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3008 (.A(net3008),
    .X(net3007));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3009 (.A(net3009),
    .X(net3008));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3010 (.A(net3014),
    .X(net3009));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3011 (.A(net3011),
    .X(net3010));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3012 (.A(net3014),
    .X(net3011));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3013 (.A(net3014),
    .X(net3012));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3014 (.A(net3014),
    .X(net3013));
 sky130_fd_sc_hd__buf_2 fanout3015 (.A(net3015),
    .X(net3014));
 sky130_fd_sc_hd__buf_12 load_slew3016 (.A(\inst$top.rst_n_sync.rst ),
    .X(net3015));
 sky130_fd_sc_hd__buf_16 wire3017 (.A(net549),
    .X(net3016));
 sky130_fd_sc_hd__buf_16 wire3018 (.A(net548),
    .X(net3017));
 sky130_fd_sc_hd__buf_16 wire3019 (.A(net546),
    .X(net3018));
 sky130_fd_sc_hd__buf_16 wire3020 (.A(net545),
    .X(net3019));
 sky130_fd_sc_hd__buf_16 wire3021 (.A(net541),
    .X(net3020));
 sky130_fd_sc_hd__buf_16 wire3022 (.A(net540),
    .X(net3021));
 sky130_fd_sc_hd__buf_16 wire3023 (.A(net539),
    .X(net3022));
 sky130_fd_sc_hd__buf_16 wire3024 (.A(net538),
    .X(net3023));
 sky130_fd_sc_hd__buf_16 wire3025 (.A(net537),
    .X(net3024));
 sky130_fd_sc_hd__buf_16 wire3026 (.A(net536),
    .X(net3025));
 sky130_fd_sc_hd__buf_16 wire3027 (.A(net535),
    .X(net3026));
 sky130_fd_sc_hd__buf_16 wire3028 (.A(net534),
    .X(net3027));
 sky130_fd_sc_hd__buf_16 wire3029 (.A(net533),
    .X(net3028));
 sky130_fd_sc_hd__buf_16 wire3030 (.A(net532),
    .X(net3029));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3031 (.A(_00128_),
    .X(net3030));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3032 (.A(_00128_),
    .X(net3031));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3033 (.A(net3033),
    .X(net3032));
 sky130_fd_sc_hd__clkdlybuf4s50_1 fanout3034 (.A(_00128_),
    .X(net3033));
 sky130_fd_sc_hd__buf_16 wire3035 (.A(gpio_in[7]),
    .X(net3034));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_regs_0_sys_clk_in (.A(clk_in),
    .X(clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_in (.A(delaynet_7_sys_clk_in),
    .X(clknet_0_clk_in));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk_in (.A(clknet_0_clk_in),
    .X(clknet_1_0__leaf_clk_in));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk_in_regs (.A(clknet_6_25__leaf_clk_in_regs),
    .X(clknet_leaf_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_1_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk_in_regs (.A(clknet_6_25__leaf_clk_in_regs),
    .X(clknet_leaf_2_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk_in_regs (.A(clknet_6_25__leaf_clk_in_regs),
    .X(clknet_leaf_4_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk_in_regs (.A(clknet_6_25__leaf_clk_in_regs),
    .X(clknet_leaf_5_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk_in_regs (.A(clknet_6_10__leaf_clk_in_regs),
    .X(clknet_leaf_6_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk_in_regs (.A(clknet_6_10__leaf_clk_in_regs),
    .X(clknet_leaf_8_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk_in_regs (.A(clknet_6_10__leaf_clk_in_regs),
    .X(clknet_leaf_9_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk_in_regs (.A(clknet_6_10__leaf_clk_in_regs),
    .X(clknet_leaf_10_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk_in_regs (.A(clknet_6_11__leaf_clk_in_regs),
    .X(clknet_leaf_11_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk_in_regs (.A(clknet_6_11__leaf_clk_in_regs),
    .X(clknet_leaf_12_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk_in_regs (.A(clknet_6_11__leaf_clk_in_regs),
    .X(clknet_leaf_13_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk_in_regs (.A(clknet_6_11__leaf_clk_in_regs),
    .X(clknet_leaf_14_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk_in_regs (.A(clknet_6_11__leaf_clk_in_regs),
    .X(clknet_leaf_15_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk_in_regs (.A(clknet_6_11__leaf_clk_in_regs),
    .X(clknet_leaf_16_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk_in_regs (.A(clknet_6_11__leaf_clk_in_regs),
    .X(clknet_leaf_17_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk_in_regs (.A(clknet_6_14__leaf_clk_in_regs),
    .X(clknet_leaf_18_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk_in_regs (.A(clknet_6_14__leaf_clk_in_regs),
    .X(clknet_leaf_19_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk_in_regs (.A(clknet_6_25__leaf_clk_in_regs),
    .X(clknet_leaf_21_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk_in_regs (.A(clknet_6_25__leaf_clk_in_regs),
    .X(clknet_leaf_22_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk_in_regs (.A(clknet_6_14__leaf_clk_in_regs),
    .X(clknet_leaf_23_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk_in_regs (.A(clknet_6_25__leaf_clk_in_regs),
    .X(clknet_leaf_24_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_25_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk_in_regs (.A(clknet_6_14__leaf_clk_in_regs),
    .X(clknet_leaf_26_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk_in_regs (.A(clknet_6_25__leaf_clk_in_regs),
    .X(clknet_leaf_27_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_28_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk_in_regs (.A(clknet_6_14__leaf_clk_in_regs),
    .X(clknet_leaf_29_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_30_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_31_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_32_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk_in_regs (.A(clknet_6_11__leaf_clk_in_regs),
    .X(clknet_leaf_33_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk_in_regs (.A(clknet_6_25__leaf_clk_in_regs),
    .X(clknet_leaf_34_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk_in_regs (.A(clknet_6_25__leaf_clk_in_regs),
    .X(clknet_leaf_35_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_36_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_37_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk_in_regs (.A(clknet_6_36__leaf_clk_in_regs),
    .X(clknet_leaf_38_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_39_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_40_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_41_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_42_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_43_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_44_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_45_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_46_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_47_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_48_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_49_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_50_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_51_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk_in_regs (.A(clknet_6_36__leaf_clk_in_regs),
    .X(clknet_leaf_52_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk_in_regs (.A(clknet_6_36__leaf_clk_in_regs),
    .X(clknet_leaf_53_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk_in_regs (.A(clknet_6_36__leaf_clk_in_regs),
    .X(clknet_leaf_54_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk_in_regs (.A(clknet_6_36__leaf_clk_in_regs),
    .X(clknet_leaf_55_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_56_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_57_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_58_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_59_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk_in_regs (.A(clknet_6_36__leaf_clk_in_regs),
    .X(clknet_leaf_60_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk_in_regs (.A(clknet_6_36__leaf_clk_in_regs),
    .X(clknet_leaf_61_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk_in_regs (.A(clknet_6_36__leaf_clk_in_regs),
    .X(clknet_leaf_62_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_63_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_64_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_65_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_66_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk_in_regs (.A(clknet_6_32__leaf_clk_in_regs),
    .X(clknet_leaf_67_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk_in_regs (.A(clknet_6_32__leaf_clk_in_regs),
    .X(clknet_leaf_68_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk_in_regs (.A(clknet_6_32__leaf_clk_in_regs),
    .X(clknet_leaf_69_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk_in_regs (.A(clknet_6_36__leaf_clk_in_regs),
    .X(clknet_leaf_70_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk_in_regs (.A(clknet_6_32__leaf_clk_in_regs),
    .X(clknet_leaf_71_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk_in_regs (.A(clknet_6_32__leaf_clk_in_regs),
    .X(clknet_leaf_72_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk_in_regs (.A(clknet_6_32__leaf_clk_in_regs),
    .X(clknet_leaf_73_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk_in_regs (.A(clknet_6_32__leaf_clk_in_regs),
    .X(clknet_leaf_74_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_75_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_76_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_77_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_78_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_79_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk_in_regs (.A(clknet_6_36__leaf_clk_in_regs),
    .X(clknet_leaf_80_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk_in_regs (.A(clknet_6_36__leaf_clk_in_regs),
    .X(clknet_leaf_81_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk_in_regs (.A(clknet_6_36__leaf_clk_in_regs),
    .X(clknet_leaf_82_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_83_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_84_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_85_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_86_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_87_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_89_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_90_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_91_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_92_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_93_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_94_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_95_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_96_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_97_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_98_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_99_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_100_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_102_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_103_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_104_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_105_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_106_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_107_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_108_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_109_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_110_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_111_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_113_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_114_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_115_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_116_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_117_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_118_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_119_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_121_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk_in_regs (.A(clknet_6_33__leaf_clk_in_regs),
    .X(clknet_leaf_123_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk_in_regs (.A(clknet_6_32__leaf_clk_in_regs),
    .X(clknet_leaf_124_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk_in_regs (.A(clknet_6_32__leaf_clk_in_regs),
    .X(clknet_leaf_127_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_128_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_129_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_130_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk_in_regs (.A(clknet_6_32__leaf_clk_in_regs),
    .X(clknet_leaf_131_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk_in_regs (.A(clknet_6_32__leaf_clk_in_regs),
    .X(clknet_leaf_132_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_134_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_135_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_138_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_140_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_143_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_144_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_145_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_146_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_147_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_148_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_149_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_150_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_151_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_152_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_153_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_154_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_155_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_156_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_157_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_158_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_159_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_160_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_161_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_162_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_163_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk_in_regs (.A(clknet_6_58__leaf_clk_in_regs),
    .X(clknet_leaf_164_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_165_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_166_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_167_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_168_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_169_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_170_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_171_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_172_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_173_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_174_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_175_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_176_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_177_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_178_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_179_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_180_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_181_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_182_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_183_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_184_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_185_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_186_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_187_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_188_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_189_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_190_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_191_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_192_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_193_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk_in_regs (.A(clknet_6_48__leaf_clk_in_regs),
    .X(clknet_leaf_194_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_195_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_196_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_197_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_198_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_199_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_200_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_201_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk_in_regs (.A(clknet_6_48__leaf_clk_in_regs),
    .X(clknet_leaf_202_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk_in_regs (.A(clknet_6_48__leaf_clk_in_regs),
    .X(clknet_leaf_203_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk_in_regs (.A(clknet_6_48__leaf_clk_in_regs),
    .X(clknet_leaf_204_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_205_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_206_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_207_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_208_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_209_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_210_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_211_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_212_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_213_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_214_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_215_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk_in_regs (.A(clknet_6_48__leaf_clk_in_regs),
    .X(clknet_leaf_216_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_217_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_218_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_219_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_220_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_221_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_222_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_223_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk_in_regs (.A(clknet_6_48__leaf_clk_in_regs),
    .X(clknet_leaf_224_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_225_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk_in_regs (.A(clknet_6_48__leaf_clk_in_regs),
    .X(clknet_leaf_226_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk_in_regs (.A(clknet_6_48__leaf_clk_in_regs),
    .X(clknet_leaf_227_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk_in_regs (.A(clknet_6_48__leaf_clk_in_regs),
    .X(clknet_leaf_228_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_229_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_231_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_232_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk_in_regs (.A(clknet_6_56__leaf_clk_in_regs),
    .X(clknet_leaf_233_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk_in_regs (.A(clknet_6_48__leaf_clk_in_regs),
    .X(clknet_leaf_236_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk_in_regs (.A(clknet_6_48__leaf_clk_in_regs),
    .X(clknet_leaf_237_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_238_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_239_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_240_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_241_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_242_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_243_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_244_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_245_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_246_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_247_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_248_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk_in_regs (.A(clknet_6_50__leaf_clk_in_regs),
    .X(clknet_leaf_249_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_250_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_251_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_252_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_253_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_254_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_255_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_256_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_clk_in_regs (.A(clknet_6_34__leaf_clk_in_regs),
    .X(clknet_leaf_257_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_258_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_259_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_260_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_261_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_262_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_263_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_264_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_265_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_266_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_clk_in_regs (.A(clknet_6_42__leaf_clk_in_regs),
    .X(clknet_leaf_267_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_268_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_269_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_270_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_271_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_272_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_273_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_274_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_274_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_275_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_275_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_276_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_276_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_277_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_277_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_278_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_278_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_279_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_279_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_280_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_280_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_281_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_281_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_282_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_282_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_283_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_283_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_284_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_284_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_285_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_285_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_286_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_286_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_287_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_287_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_288_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_288_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_289_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_289_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_290_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_290_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_291_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_291_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_292_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_292_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_293_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_293_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_294_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_294_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_295_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_295_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_296_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_296_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_297_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_297_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_298_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_298_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_299_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_299_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_300_clk_in_regs (.A(clknet_6_40__leaf_clk_in_regs),
    .X(clknet_leaf_300_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_302_clk_in_regs (.A(clknet_6_41__leaf_clk_in_regs),
    .X(clknet_leaf_302_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_303_clk_in_regs (.A(clknet_6_41__leaf_clk_in_regs),
    .X(clknet_leaf_303_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_304_clk_in_regs (.A(clknet_6_38__leaf_clk_in_regs),
    .X(clknet_leaf_304_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_305_clk_in_regs (.A(clknet_6_38__leaf_clk_in_regs),
    .X(clknet_leaf_305_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_308_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_308_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_309_clk_in_regs (.A(clknet_6_38__leaf_clk_in_regs),
    .X(clknet_leaf_309_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_310_clk_in_regs (.A(clknet_6_35__leaf_clk_in_regs),
    .X(clknet_leaf_310_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_311_clk_in_regs (.A(clknet_6_38__leaf_clk_in_regs),
    .X(clknet_leaf_311_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_312_clk_in_regs (.A(clknet_6_38__leaf_clk_in_regs),
    .X(clknet_leaf_312_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_313_clk_in_regs (.A(clknet_6_38__leaf_clk_in_regs),
    .X(clknet_leaf_313_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_314_clk_in_regs (.A(clknet_6_38__leaf_clk_in_regs),
    .X(clknet_leaf_314_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_315_clk_in_regs (.A(clknet_6_38__leaf_clk_in_regs),
    .X(clknet_leaf_315_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_316_clk_in_regs (.A(clknet_6_38__leaf_clk_in_regs),
    .X(clknet_leaf_316_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_317_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_317_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_318_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_318_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_319_clk_in_regs (.A(clknet_6_39__leaf_clk_in_regs),
    .X(clknet_leaf_319_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_320_clk_in_regs (.A(clknet_6_38__leaf_clk_in_regs),
    .X(clknet_leaf_320_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_321_clk_in_regs (.A(clknet_6_38__leaf_clk_in_regs),
    .X(clknet_leaf_321_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_322_clk_in_regs (.A(clknet_6_39__leaf_clk_in_regs),
    .X(clknet_leaf_322_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_323_clk_in_regs (.A(clknet_6_38__leaf_clk_in_regs),
    .X(clknet_leaf_323_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_324_clk_in_regs (.A(clknet_6_39__leaf_clk_in_regs),
    .X(clknet_leaf_324_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_325_clk_in_regs (.A(clknet_6_39__leaf_clk_in_regs),
    .X(clknet_leaf_325_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_327_clk_in_regs (.A(clknet_6_39__leaf_clk_in_regs),
    .X(clknet_leaf_327_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_328_clk_in_regs (.A(clknet_6_39__leaf_clk_in_regs),
    .X(clknet_leaf_328_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_329_clk_in_regs (.A(clknet_6_37__leaf_clk_in_regs),
    .X(clknet_leaf_329_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_330_clk_in_regs (.A(clknet_6_14__leaf_clk_in_regs),
    .X(clknet_leaf_330_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_331_clk_in_regs (.A(clknet_6_14__leaf_clk_in_regs),
    .X(clknet_leaf_331_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_332_clk_in_regs (.A(clknet_6_14__leaf_clk_in_regs),
    .X(clknet_leaf_332_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_333_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_333_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_334_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_334_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_335_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_335_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_337_clk_in_regs (.A(clknet_6_27__leaf_clk_in_regs),
    .X(clknet_leaf_337_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_338_clk_in_regs (.A(clknet_6_39__leaf_clk_in_regs),
    .X(clknet_leaf_338_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_339_clk_in_regs (.A(clknet_6_39__leaf_clk_in_regs),
    .X(clknet_leaf_339_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_340_clk_in_regs (.A(clknet_6_39__leaf_clk_in_regs),
    .X(clknet_leaf_340_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_341_clk_in_regs (.A(clknet_6_45__leaf_clk_in_regs),
    .X(clknet_leaf_341_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_342_clk_in_regs (.A(clknet_6_39__leaf_clk_in_regs),
    .X(clknet_leaf_342_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_343_clk_in_regs (.A(clknet_6_27__leaf_clk_in_regs),
    .X(clknet_leaf_343_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_344_clk_in_regs (.A(clknet_6_27__leaf_clk_in_regs),
    .X(clknet_leaf_344_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_345_clk_in_regs (.A(clknet_6_27__leaf_clk_in_regs),
    .X(clknet_leaf_345_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_346_clk_in_regs (.A(clknet_6_45__leaf_clk_in_regs),
    .X(clknet_leaf_346_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_347_clk_in_regs (.A(clknet_6_45__leaf_clk_in_regs),
    .X(clknet_leaf_347_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_348_clk_in_regs (.A(clknet_6_45__leaf_clk_in_regs),
    .X(clknet_leaf_348_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_349_clk_in_regs (.A(clknet_6_45__leaf_clk_in_regs),
    .X(clknet_leaf_349_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_350_clk_in_regs (.A(clknet_6_45__leaf_clk_in_regs),
    .X(clknet_leaf_350_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_351_clk_in_regs (.A(clknet_6_44__leaf_clk_in_regs),
    .X(clknet_leaf_351_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_352_clk_in_regs (.A(clknet_6_44__leaf_clk_in_regs),
    .X(clknet_leaf_352_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_353_clk_in_regs (.A(clknet_6_45__leaf_clk_in_regs),
    .X(clknet_leaf_353_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_354_clk_in_regs (.A(clknet_6_45__leaf_clk_in_regs),
    .X(clknet_leaf_354_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_355_clk_in_regs (.A(clknet_6_45__leaf_clk_in_regs),
    .X(clknet_leaf_355_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_356_clk_in_regs (.A(clknet_6_41__leaf_clk_in_regs),
    .X(clknet_leaf_356_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_357_clk_in_regs (.A(clknet_6_41__leaf_clk_in_regs),
    .X(clknet_leaf_357_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_358_clk_in_regs (.A(clknet_6_41__leaf_clk_in_regs),
    .X(clknet_leaf_358_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_359_clk_in_regs (.A(clknet_6_44__leaf_clk_in_regs),
    .X(clknet_leaf_359_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_360_clk_in_regs (.A(clknet_6_44__leaf_clk_in_regs),
    .X(clknet_leaf_360_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_361_clk_in_regs (.A(clknet_6_41__leaf_clk_in_regs),
    .X(clknet_leaf_361_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_362_clk_in_regs (.A(clknet_6_41__leaf_clk_in_regs),
    .X(clknet_leaf_362_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_363_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_363_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_364_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_364_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_365_clk_in_regs (.A(clknet_6_52__leaf_clk_in_regs),
    .X(clknet_leaf_365_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_366_clk_in_regs (.A(clknet_6_52__leaf_clk_in_regs),
    .X(clknet_leaf_366_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_367_clk_in_regs (.A(clknet_6_43__leaf_clk_in_regs),
    .X(clknet_leaf_367_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_368_clk_in_regs (.A(clknet_6_41__leaf_clk_in_regs),
    .X(clknet_leaf_368_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_369_clk_in_regs (.A(clknet_6_44__leaf_clk_in_regs),
    .X(clknet_leaf_369_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_370_clk_in_regs (.A(clknet_6_44__leaf_clk_in_regs),
    .X(clknet_leaf_370_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_371_clk_in_regs (.A(clknet_6_52__leaf_clk_in_regs),
    .X(clknet_leaf_371_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_372_clk_in_regs (.A(clknet_6_52__leaf_clk_in_regs),
    .X(clknet_leaf_372_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_373_clk_in_regs (.A(clknet_6_52__leaf_clk_in_regs),
    .X(clknet_leaf_373_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_374_clk_in_regs (.A(clknet_6_52__leaf_clk_in_regs),
    .X(clknet_leaf_374_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_375_clk_in_regs (.A(clknet_6_46__leaf_clk_in_regs),
    .X(clknet_leaf_375_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_376_clk_in_regs (.A(clknet_6_44__leaf_clk_in_regs),
    .X(clknet_leaf_376_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_377_clk_in_regs (.A(clknet_6_44__leaf_clk_in_regs),
    .X(clknet_leaf_377_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_378_clk_in_regs (.A(clknet_6_44__leaf_clk_in_regs),
    .X(clknet_leaf_378_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_379_clk_in_regs (.A(clknet_6_44__leaf_clk_in_regs),
    .X(clknet_leaf_379_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_381_clk_in_regs (.A(clknet_6_45__leaf_clk_in_regs),
    .X(clknet_leaf_381_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_383_clk_in_regs (.A(clknet_6_45__leaf_clk_in_regs),
    .X(clknet_leaf_383_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_384_clk_in_regs (.A(clknet_6_44__leaf_clk_in_regs),
    .X(clknet_leaf_384_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_385_clk_in_regs (.A(clknet_6_44__leaf_clk_in_regs),
    .X(clknet_leaf_385_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_387_clk_in_regs (.A(clknet_6_46__leaf_clk_in_regs),
    .X(clknet_leaf_387_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_388_clk_in_regs (.A(clknet_6_46__leaf_clk_in_regs),
    .X(clknet_leaf_388_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_389_clk_in_regs (.A(clknet_6_46__leaf_clk_in_regs),
    .X(clknet_leaf_389_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_390_clk_in_regs (.A(clknet_6_52__leaf_clk_in_regs),
    .X(clknet_leaf_390_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_391_clk_in_regs (.A(clknet_6_46__leaf_clk_in_regs),
    .X(clknet_leaf_391_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_392_clk_in_regs (.A(clknet_6_53__leaf_clk_in_regs),
    .X(clknet_leaf_392_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_393_clk_in_regs (.A(clknet_6_52__leaf_clk_in_regs),
    .X(clknet_leaf_393_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_394_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_394_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_395_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_395_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_396_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_396_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_397_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_397_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_398_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_398_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_399_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_399_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_400_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_400_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_401_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_401_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_402_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_402_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_403_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_403_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_404_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_404_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_405_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_405_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_406_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_406_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_407_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_407_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_408_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_408_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_409_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_409_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_410_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_410_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_411_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_411_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_412_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_412_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_413_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_413_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_414_clk_in_regs (.A(clknet_6_52__leaf_clk_in_regs),
    .X(clknet_leaf_414_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_415_clk_in_regs (.A(clknet_6_55__leaf_clk_in_regs),
    .X(clknet_leaf_415_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_416_clk_in_regs (.A(clknet_6_54__leaf_clk_in_regs),
    .X(clknet_leaf_416_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_417_clk_in_regs (.A(clknet_6_54__leaf_clk_in_regs),
    .X(clknet_leaf_417_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_418_clk_in_regs (.A(clknet_6_54__leaf_clk_in_regs),
    .X(clknet_leaf_418_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_419_clk_in_regs (.A(clknet_6_54__leaf_clk_in_regs),
    .X(clknet_leaf_419_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_421_clk_in_regs (.A(clknet_6_54__leaf_clk_in_regs),
    .X(clknet_leaf_421_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_423_clk_in_regs (.A(clknet_6_54__leaf_clk_in_regs),
    .X(clknet_leaf_423_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_424_clk_in_regs (.A(clknet_6_51__leaf_clk_in_regs),
    .X(clknet_leaf_424_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_425_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_425_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_426_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_426_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_427_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_427_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_428_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_428_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_429_clk_in_regs (.A(clknet_6_54__leaf_clk_in_regs),
    .X(clknet_leaf_429_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_430_clk_in_regs (.A(clknet_6_54__leaf_clk_in_regs),
    .X(clknet_leaf_430_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_431_clk_in_regs (.A(clknet_6_54__leaf_clk_in_regs),
    .X(clknet_leaf_431_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_432_clk_in_regs (.A(clknet_6_54__leaf_clk_in_regs),
    .X(clknet_leaf_432_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_433_clk_in_regs (.A(clknet_6_49__leaf_clk_in_regs),
    .X(clknet_leaf_433_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_434_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_434_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_435_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_435_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_436_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_436_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_437_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_437_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_438_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_438_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_439_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_439_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_440_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_440_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_441_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_441_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_442_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_442_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_443_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_443_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_444_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_444_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_445_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_445_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_446_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_446_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_447_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_447_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_448_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_448_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_449_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_449_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_450_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_450_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_451_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_451_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_452_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_452_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_453_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_453_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_454_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_454_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_455_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_455_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_456_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_456_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_457_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_457_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_458_clk_in_regs (.A(clknet_6_57__leaf_clk_in_regs),
    .X(clknet_leaf_458_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_459_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_459_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_460_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_460_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_461_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_461_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_462_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_462_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_463_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_463_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_464_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_464_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_465_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_465_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_466_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_466_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_467_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_467_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_468_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_468_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_469_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_469_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_470_clk_in_regs (.A(clknet_6_59__leaf_clk_in_regs),
    .X(clknet_leaf_470_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_471_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_471_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_472_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_472_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_473_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_473_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_474_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_474_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_475_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_475_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_476_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_476_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_477_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_477_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_478_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_478_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_479_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_479_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_480_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_480_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_481_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_481_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_482_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_482_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_483_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_483_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_484_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_484_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_485_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_485_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_486_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_486_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_487_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_487_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_488_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_488_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_489_clk_in_regs (.A(clknet_6_62__leaf_clk_in_regs),
    .X(clknet_leaf_489_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_490_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_490_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_491_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_491_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_492_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_492_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_493_clk_in_regs (.A(clknet_6_60__leaf_clk_in_regs),
    .X(clknet_leaf_493_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_494_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_494_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_495_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_495_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_496_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_496_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_497_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_497_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_498_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_498_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_499_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_499_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_500_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_500_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_501_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_501_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_502_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_502_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_503_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_503_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_504_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_504_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_505_clk_in_regs (.A(clknet_6_63__leaf_clk_in_regs),
    .X(clknet_leaf_505_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_506_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_506_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_507_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_507_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_508_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_508_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_509_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_509_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_510_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_510_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_511_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_511_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_512_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_512_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_513_clk_in_regs (.A(clknet_6_61__leaf_clk_in_regs),
    .X(clknet_leaf_513_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_515_clk_in_regs (.A(clknet_6_53__leaf_clk_in_regs),
    .X(clknet_leaf_515_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_519_clk_in_regs (.A(clknet_6_47__leaf_clk_in_regs),
    .X(clknet_leaf_519_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_520_clk_in_regs (.A(clknet_6_22__leaf_clk_in_regs),
    .X(clknet_leaf_520_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_525_clk_in_regs (.A(clknet_6_53__leaf_clk_in_regs),
    .X(clknet_leaf_525_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_527_clk_in_regs (.A(clknet_6_47__leaf_clk_in_regs),
    .X(clknet_leaf_527_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_528_clk_in_regs (.A(clknet_6_47__leaf_clk_in_regs),
    .X(clknet_leaf_528_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_529_clk_in_regs (.A(clknet_6_53__leaf_clk_in_regs),
    .X(clknet_leaf_529_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_530_clk_in_regs (.A(clknet_6_47__leaf_clk_in_regs),
    .X(clknet_leaf_530_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_531_clk_in_regs (.A(clknet_6_47__leaf_clk_in_regs),
    .X(clknet_leaf_531_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_532_clk_in_regs (.A(clknet_6_47__leaf_clk_in_regs),
    .X(clknet_leaf_532_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_533_clk_in_regs (.A(clknet_6_47__leaf_clk_in_regs),
    .X(clknet_leaf_533_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_534_clk_in_regs (.A(clknet_6_47__leaf_clk_in_regs),
    .X(clknet_leaf_534_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_535_clk_in_regs (.A(clknet_6_47__leaf_clk_in_regs),
    .X(clknet_leaf_535_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_536_clk_in_regs (.A(clknet_6_23__leaf_clk_in_regs),
    .X(clknet_leaf_536_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_537_clk_in_regs (.A(clknet_6_23__leaf_clk_in_regs),
    .X(clknet_leaf_537_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_538_clk_in_regs (.A(clknet_6_23__leaf_clk_in_regs),
    .X(clknet_leaf_538_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_542_clk_in_regs (.A(clknet_6_23__leaf_clk_in_regs),
    .X(clknet_leaf_542_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_543_clk_in_regs (.A(clknet_6_23__leaf_clk_in_regs),
    .X(clknet_leaf_543_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_544_clk_in_regs (.A(clknet_6_23__leaf_clk_in_regs),
    .X(clknet_leaf_544_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_545_clk_in_regs (.A(clknet_6_23__leaf_clk_in_regs),
    .X(clknet_leaf_545_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_546_clk_in_regs (.A(clknet_6_21__leaf_clk_in_regs),
    .X(clknet_leaf_546_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_547_clk_in_regs (.A(clknet_6_21__leaf_clk_in_regs),
    .X(clknet_leaf_547_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_549_clk_in_regs (.A(clknet_6_21__leaf_clk_in_regs),
    .X(clknet_leaf_549_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_550_clk_in_regs (.A(clknet_6_21__leaf_clk_in_regs),
    .X(clknet_leaf_550_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_551_clk_in_regs (.A(clknet_6_20__leaf_clk_in_regs),
    .X(clknet_leaf_551_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_554_clk_in_regs (.A(clknet_6_22__leaf_clk_in_regs),
    .X(clknet_leaf_554_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_555_clk_in_regs (.A(clknet_6_20__leaf_clk_in_regs),
    .X(clknet_leaf_555_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_557_clk_in_regs (.A(clknet_6_22__leaf_clk_in_regs),
    .X(clknet_leaf_557_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_559_clk_in_regs (.A(clknet_6_22__leaf_clk_in_regs),
    .X(clknet_leaf_559_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_560_clk_in_regs (.A(clknet_6_46__leaf_clk_in_regs),
    .X(clknet_leaf_560_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_561_clk_in_regs (.A(clknet_6_45__leaf_clk_in_regs),
    .X(clknet_leaf_561_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_562_clk_in_regs (.A(clknet_6_31__leaf_clk_in_regs),
    .X(clknet_leaf_562_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_564_clk_in_regs (.A(clknet_6_20__leaf_clk_in_regs),
    .X(clknet_leaf_564_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_565_clk_in_regs (.A(clknet_6_20__leaf_clk_in_regs),
    .X(clknet_leaf_565_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_566_clk_in_regs (.A(clknet_6_19__leaf_clk_in_regs),
    .X(clknet_leaf_566_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_567_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_567_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_568_clk_in_regs (.A(clknet_6_20__leaf_clk_in_regs),
    .X(clknet_leaf_568_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_570_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_570_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_572_clk_in_regs (.A(clknet_6_31__leaf_clk_in_regs),
    .X(clknet_leaf_572_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_573_clk_in_regs (.A(clknet_6_31__leaf_clk_in_regs),
    .X(clknet_leaf_573_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_574_clk_in_regs (.A(clknet_6_31__leaf_clk_in_regs),
    .X(clknet_leaf_574_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_575_clk_in_regs (.A(clknet_6_31__leaf_clk_in_regs),
    .X(clknet_leaf_575_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_576_clk_in_regs (.A(clknet_6_31__leaf_clk_in_regs),
    .X(clknet_leaf_576_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_577_clk_in_regs (.A(clknet_6_31__leaf_clk_in_regs),
    .X(clknet_leaf_577_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_578_clk_in_regs (.A(clknet_6_31__leaf_clk_in_regs),
    .X(clknet_leaf_578_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_579_clk_in_regs (.A(clknet_6_31__leaf_clk_in_regs),
    .X(clknet_leaf_579_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_580_clk_in_regs (.A(clknet_6_27__leaf_clk_in_regs),
    .X(clknet_leaf_580_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_584_clk_in_regs (.A(clknet_6_27__leaf_clk_in_regs),
    .X(clknet_leaf_584_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_585_clk_in_regs (.A(clknet_6_15__leaf_clk_in_regs),
    .X(clknet_leaf_585_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_586_clk_in_regs (.A(clknet_6_27__leaf_clk_in_regs),
    .X(clknet_leaf_586_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_587_clk_in_regs (.A(clknet_6_15__leaf_clk_in_regs),
    .X(clknet_leaf_587_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_588_clk_in_regs (.A(clknet_6_27__leaf_clk_in_regs),
    .X(clknet_leaf_588_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_589_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_589_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_590_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_590_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_591_clk_in_regs (.A(clknet_6_15__leaf_clk_in_regs),
    .X(clknet_leaf_591_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_592_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_592_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_593_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_593_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_594_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_594_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_595_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_595_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_596_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_596_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_597_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_597_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_598_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_598_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_599_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_599_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_600_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_600_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_601_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_601_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_602_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_602_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_603_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_603_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_604_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_604_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_605_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_605_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_606_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_606_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_607_clk_in_regs (.A(clknet_6_15__leaf_clk_in_regs),
    .X(clknet_leaf_607_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_608_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_608_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_609_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_609_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_610_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_610_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_611_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_611_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_612_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_612_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_613_clk_in_regs (.A(clknet_6_3__leaf_clk_in_regs),
    .X(clknet_leaf_613_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_614_clk_in_regs (.A(clknet_6_3__leaf_clk_in_regs),
    .X(clknet_leaf_614_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_615_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_615_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_616_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_616_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_617_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_617_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_618_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_618_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_619_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_619_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_620_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_620_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_621_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_621_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_622_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_622_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_623_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_623_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_624_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_624_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_625_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_625_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_626_clk_in_regs (.A(clknet_6_30__leaf_clk_in_regs),
    .X(clknet_leaf_626_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_627_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_627_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_628_clk_in_regs (.A(clknet_6_28__leaf_clk_in_regs),
    .X(clknet_leaf_628_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_629_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_629_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_630_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_630_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_632_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_632_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_633_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_633_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_634_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_634_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_635_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_635_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_636_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_636_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_637_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_637_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_638_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_638_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_640_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_640_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_641_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_641_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_642_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_642_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_643_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_643_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_644_clk_in_regs (.A(clknet_6_7__leaf_clk_in_regs),
    .X(clknet_leaf_644_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_645_clk_in_regs (.A(clknet_6_7__leaf_clk_in_regs),
    .X(clknet_leaf_645_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_646_clk_in_regs (.A(clknet_6_7__leaf_clk_in_regs),
    .X(clknet_leaf_646_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_647_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_647_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_648_clk_in_regs (.A(clknet_6_29__leaf_clk_in_regs),
    .X(clknet_leaf_648_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_649_clk_in_regs (.A(clknet_6_6__leaf_clk_in_regs),
    .X(clknet_leaf_649_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_650_clk_in_regs (.A(clknet_6_6__leaf_clk_in_regs),
    .X(clknet_leaf_650_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_651_clk_in_regs (.A(clknet_6_3__leaf_clk_in_regs),
    .X(clknet_leaf_651_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_652_clk_in_regs (.A(clknet_6_3__leaf_clk_in_regs),
    .X(clknet_leaf_652_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_653_clk_in_regs (.A(clknet_6_3__leaf_clk_in_regs),
    .X(clknet_leaf_653_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_654_clk_in_regs (.A(clknet_6_3__leaf_clk_in_regs),
    .X(clknet_leaf_654_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_655_clk_in_regs (.A(clknet_6_3__leaf_clk_in_regs),
    .X(clknet_leaf_655_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_656_clk_in_regs (.A(clknet_6_6__leaf_clk_in_regs),
    .X(clknet_leaf_656_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_657_clk_in_regs (.A(clknet_6_6__leaf_clk_in_regs),
    .X(clknet_leaf_657_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_658_clk_in_regs (.A(clknet_6_6__leaf_clk_in_regs),
    .X(clknet_leaf_658_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_659_clk_in_regs (.A(clknet_6_4__leaf_clk_in_regs),
    .X(clknet_leaf_659_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_660_clk_in_regs (.A(clknet_6_4__leaf_clk_in_regs),
    .X(clknet_leaf_660_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_661_clk_in_regs (.A(clknet_6_4__leaf_clk_in_regs),
    .X(clknet_leaf_661_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_662_clk_in_regs (.A(clknet_6_6__leaf_clk_in_regs),
    .X(clknet_leaf_662_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_663_clk_in_regs (.A(clknet_6_7__leaf_clk_in_regs),
    .X(clknet_leaf_663_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_664_clk_in_regs (.A(clknet_6_7__leaf_clk_in_regs),
    .X(clknet_leaf_664_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_665_clk_in_regs (.A(clknet_6_7__leaf_clk_in_regs),
    .X(clknet_leaf_665_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_666_clk_in_regs (.A(clknet_6_5__leaf_clk_in_regs),
    .X(clknet_leaf_666_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_667_clk_in_regs (.A(clknet_6_5__leaf_clk_in_regs),
    .X(clknet_leaf_667_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_669_clk_in_regs (.A(clknet_6_16__leaf_clk_in_regs),
    .X(clknet_leaf_669_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_671_clk_in_regs (.A(clknet_6_16__leaf_clk_in_regs),
    .X(clknet_leaf_671_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_672_clk_in_regs (.A(clknet_6_16__leaf_clk_in_regs),
    .X(clknet_leaf_672_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_673_clk_in_regs (.A(clknet_6_16__leaf_clk_in_regs),
    .X(clknet_leaf_673_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_675_clk_in_regs (.A(clknet_6_16__leaf_clk_in_regs),
    .X(clknet_leaf_675_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_678_clk_in_regs (.A(clknet_6_16__leaf_clk_in_regs),
    .X(clknet_leaf_678_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_679_clk_in_regs (.A(clknet_6_16__leaf_clk_in_regs),
    .X(clknet_leaf_679_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_680_clk_in_regs (.A(clknet_6_16__leaf_clk_in_regs),
    .X(clknet_leaf_680_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_681_clk_in_regs (.A(clknet_6_16__leaf_clk_in_regs),
    .X(clknet_leaf_681_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_682_clk_in_regs (.A(clknet_6_16__leaf_clk_in_regs),
    .X(clknet_leaf_682_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_683_clk_in_regs (.A(clknet_6_19__leaf_clk_in_regs),
    .X(clknet_leaf_683_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_684_clk_in_regs (.A(clknet_6_19__leaf_clk_in_regs),
    .X(clknet_leaf_684_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_685_clk_in_regs (.A(clknet_6_19__leaf_clk_in_regs),
    .X(clknet_leaf_685_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_686_clk_in_regs (.A(clknet_6_19__leaf_clk_in_regs),
    .X(clknet_leaf_686_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_687_clk_in_regs (.A(clknet_6_19__leaf_clk_in_regs),
    .X(clknet_leaf_687_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_688_clk_in_regs (.A(clknet_6_18__leaf_clk_in_regs),
    .X(clknet_leaf_688_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_689_clk_in_regs (.A(clknet_6_18__leaf_clk_in_regs),
    .X(clknet_leaf_689_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_690_clk_in_regs (.A(clknet_6_19__leaf_clk_in_regs),
    .X(clknet_leaf_690_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_691_clk_in_regs (.A(clknet_6_19__leaf_clk_in_regs),
    .X(clknet_leaf_691_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_692_clk_in_regs (.A(clknet_6_18__leaf_clk_in_regs),
    .X(clknet_leaf_692_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_694_clk_in_regs (.A(clknet_6_18__leaf_clk_in_regs),
    .X(clknet_leaf_694_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_695_clk_in_regs (.A(clknet_6_21__leaf_clk_in_regs),
    .X(clknet_leaf_695_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_696_clk_in_regs (.A(clknet_6_17__leaf_clk_in_regs),
    .X(clknet_leaf_696_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_697_clk_in_regs (.A(clknet_6_17__leaf_clk_in_regs),
    .X(clknet_leaf_697_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_698_clk_in_regs (.A(clknet_6_16__leaf_clk_in_regs),
    .X(clknet_leaf_698_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_700_clk_in_regs (.A(clknet_6_17__leaf_clk_in_regs),
    .X(clknet_leaf_700_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_701_clk_in_regs (.A(clknet_6_16__leaf_clk_in_regs),
    .X(clknet_leaf_701_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_702_clk_in_regs (.A(clknet_6_17__leaf_clk_in_regs),
    .X(clknet_leaf_702_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_703_clk_in_regs (.A(clknet_6_17__leaf_clk_in_regs),
    .X(clknet_leaf_703_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_704_clk_in_regs (.A(clknet_6_17__leaf_clk_in_regs),
    .X(clknet_leaf_704_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_705_clk_in_regs (.A(clknet_6_17__leaf_clk_in_regs),
    .X(clknet_leaf_705_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_706_clk_in_regs (.A(clknet_6_18__leaf_clk_in_regs),
    .X(clknet_leaf_706_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_707_clk_in_regs (.A(clknet_6_21__leaf_clk_in_regs),
    .X(clknet_leaf_707_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_708_clk_in_regs (.A(clknet_6_17__leaf_clk_in_regs),
    .X(clknet_leaf_708_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_709_clk_in_regs (.A(clknet_6_18__leaf_clk_in_regs),
    .X(clknet_leaf_709_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_711_clk_in_regs (.A(clknet_6_17__leaf_clk_in_regs),
    .X(clknet_leaf_711_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_712_clk_in_regs (.A(clknet_6_17__leaf_clk_in_regs),
    .X(clknet_leaf_712_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_715_clk_in_regs (.A(clknet_6_4__leaf_clk_in_regs),
    .X(clknet_leaf_715_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_716_clk_in_regs (.A(clknet_6_1__leaf_clk_in_regs),
    .X(clknet_leaf_716_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_717_clk_in_regs (.A(clknet_6_1__leaf_clk_in_regs),
    .X(clknet_leaf_717_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_718_clk_in_regs (.A(clknet_6_2__leaf_clk_in_regs),
    .X(clknet_leaf_718_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_719_clk_in_regs (.A(clknet_6_2__leaf_clk_in_regs),
    .X(clknet_leaf_719_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_720_clk_in_regs (.A(clknet_6_2__leaf_clk_in_regs),
    .X(clknet_leaf_720_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_721_clk_in_regs (.A(clknet_6_2__leaf_clk_in_regs),
    .X(clknet_leaf_721_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_722_clk_in_regs (.A(clknet_6_1__leaf_clk_in_regs),
    .X(clknet_leaf_722_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_723_clk_in_regs (.A(clknet_6_1__leaf_clk_in_regs),
    .X(clknet_leaf_723_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_724_clk_in_regs (.A(clknet_6_1__leaf_clk_in_regs),
    .X(clknet_leaf_724_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_725_clk_in_regs (.A(clknet_6_0__leaf_clk_in_regs),
    .X(clknet_leaf_725_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_726_clk_in_regs (.A(clknet_6_0__leaf_clk_in_regs),
    .X(clknet_leaf_726_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_727_clk_in_regs (.A(clknet_6_0__leaf_clk_in_regs),
    .X(clknet_leaf_727_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_728_clk_in_regs (.A(clknet_6_12__leaf_clk_in_regs),
    .X(clknet_leaf_728_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_729_clk_in_regs (.A(clknet_6_0__leaf_clk_in_regs),
    .X(clknet_leaf_729_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_730_clk_in_regs (.A(clknet_6_2__leaf_clk_in_regs),
    .X(clknet_leaf_730_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_731_clk_in_regs (.A(clknet_6_1__leaf_clk_in_regs),
    .X(clknet_leaf_731_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_732_clk_in_regs (.A(clknet_6_0__leaf_clk_in_regs),
    .X(clknet_leaf_732_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_733_clk_in_regs (.A(clknet_6_1__leaf_clk_in_regs),
    .X(clknet_leaf_733_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_734_clk_in_regs (.A(clknet_6_2__leaf_clk_in_regs),
    .X(clknet_leaf_734_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_735_clk_in_regs (.A(clknet_6_2__leaf_clk_in_regs),
    .X(clknet_leaf_735_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_736_clk_in_regs (.A(clknet_6_2__leaf_clk_in_regs),
    .X(clknet_leaf_736_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_737_clk_in_regs (.A(clknet_6_2__leaf_clk_in_regs),
    .X(clknet_leaf_737_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_738_clk_in_regs (.A(clknet_6_3__leaf_clk_in_regs),
    .X(clknet_leaf_738_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_739_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_739_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_740_clk_in_regs (.A(clknet_6_2__leaf_clk_in_regs),
    .X(clknet_leaf_740_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_741_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_741_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_742_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_742_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_743_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_743_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_744_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_744_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_745_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_745_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_746_clk_in_regs (.A(clknet_6_12__leaf_clk_in_regs),
    .X(clknet_leaf_746_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_748_clk_in_regs (.A(clknet_6_12__leaf_clk_in_regs),
    .X(clknet_leaf_748_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_749_clk_in_regs (.A(clknet_6_12__leaf_clk_in_regs),
    .X(clknet_leaf_749_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_750_clk_in_regs (.A(clknet_6_12__leaf_clk_in_regs),
    .X(clknet_leaf_750_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_751_clk_in_regs (.A(clknet_6_12__leaf_clk_in_regs),
    .X(clknet_leaf_751_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_752_clk_in_regs (.A(clknet_6_15__leaf_clk_in_regs),
    .X(clknet_leaf_752_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_753_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_753_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_754_clk_in_regs (.A(clknet_6_13__leaf_clk_in_regs),
    .X(clknet_leaf_754_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_755_clk_in_regs (.A(clknet_6_15__leaf_clk_in_regs),
    .X(clknet_leaf_755_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_756_clk_in_regs (.A(clknet_6_15__leaf_clk_in_regs),
    .X(clknet_leaf_756_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_757_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_757_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_758_clk_in_regs (.A(clknet_6_26__leaf_clk_in_regs),
    .X(clknet_leaf_758_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_759_clk_in_regs (.A(clknet_6_14__leaf_clk_in_regs),
    .X(clknet_leaf_759_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_760_clk_in_regs (.A(clknet_6_12__leaf_clk_in_regs),
    .X(clknet_leaf_760_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_761_clk_in_regs (.A(clknet_6_12__leaf_clk_in_regs),
    .X(clknet_leaf_761_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_762_clk_in_regs (.A(clknet_6_9__leaf_clk_in_regs),
    .X(clknet_leaf_762_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_763_clk_in_regs (.A(clknet_6_9__leaf_clk_in_regs),
    .X(clknet_leaf_763_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_764_clk_in_regs (.A(clknet_6_9__leaf_clk_in_regs),
    .X(clknet_leaf_764_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_765_clk_in_regs (.A(clknet_6_8__leaf_clk_in_regs),
    .X(clknet_leaf_765_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_766_clk_in_regs (.A(clknet_6_9__leaf_clk_in_regs),
    .X(clknet_leaf_766_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_767_clk_in_regs (.A(clknet_6_9__leaf_clk_in_regs),
    .X(clknet_leaf_767_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_768_clk_in_regs (.A(clknet_6_11__leaf_clk_in_regs),
    .X(clknet_leaf_768_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_769_clk_in_regs (.A(clknet_6_11__leaf_clk_in_regs),
    .X(clknet_leaf_769_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_770_clk_in_regs (.A(clknet_6_8__leaf_clk_in_regs),
    .X(clknet_leaf_770_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_771_clk_in_regs (.A(clknet_6_8__leaf_clk_in_regs),
    .X(clknet_leaf_771_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_772_clk_in_regs (.A(clknet_6_8__leaf_clk_in_regs),
    .X(clknet_leaf_772_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_773_clk_in_regs (.A(clknet_6_8__leaf_clk_in_regs),
    .X(clknet_leaf_773_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_774_clk_in_regs (.A(clknet_6_8__leaf_clk_in_regs),
    .X(clknet_leaf_774_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_776_clk_in_regs (.A(clknet_6_8__leaf_clk_in_regs),
    .X(clknet_leaf_776_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_777_clk_in_regs (.A(clknet_6_8__leaf_clk_in_regs),
    .X(clknet_leaf_777_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_778_clk_in_regs (.A(clknet_6_9__leaf_clk_in_regs),
    .X(clknet_leaf_778_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_779_clk_in_regs (.A(clknet_6_9__leaf_clk_in_regs),
    .X(clknet_leaf_779_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_781_clk_in_regs (.A(clknet_6_10__leaf_clk_in_regs),
    .X(clknet_leaf_781_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_783_clk_in_regs (.A(clknet_6_10__leaf_clk_in_regs),
    .X(clknet_leaf_783_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_784_clk_in_regs (.A(clknet_6_10__leaf_clk_in_regs),
    .X(clknet_leaf_784_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_785_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_785_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_786_clk_in_regs (.A(clknet_6_10__leaf_clk_in_regs),
    .X(clknet_leaf_786_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_787_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_787_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_788_clk_in_regs (.A(clknet_6_24__leaf_clk_in_regs),
    .X(clknet_leaf_788_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_789_clk_in_regs (.A(clknet_6_10__leaf_clk_in_regs),
    .X(clknet_leaf_789_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_790_clk_in_regs (.A(clknet_6_10__leaf_clk_in_regs),
    .X(clknet_leaf_790_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_in_regs (.A(clk_in_regs),
    .X(clknet_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0_0_clk_in_regs (.A(clknet_0_clk_in_regs),
    .X(clknet_1_0_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1_0_clk_in_regs (.A(clknet_0_clk_in_regs),
    .X(clknet_1_1_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0_0_clk_in_regs (.A(clknet_1_0_0_clk_in_regs),
    .X(clknet_3_0_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1_0_clk_in_regs (.A(clknet_1_0_0_clk_in_regs),
    .X(clknet_3_1_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2_0_clk_in_regs (.A(clknet_1_0_0_clk_in_regs),
    .X(clknet_3_2_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3_0_clk_in_regs (.A(clknet_1_0_0_clk_in_regs),
    .X(clknet_3_3_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4_0_clk_in_regs (.A(clknet_1_1_0_clk_in_regs),
    .X(clknet_3_4_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5_0_clk_in_regs (.A(clknet_1_1_0_clk_in_regs),
    .X(clknet_3_5_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6_0_clk_in_regs (.A(clknet_1_1_0_clk_in_regs),
    .X(clknet_3_6_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7_0_clk_in_regs (.A(clknet_1_1_0_clk_in_regs),
    .X(clknet_3_7_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_0_0_clk_in_regs (.A(clknet_3_0_0_clk_in_regs),
    .X(clknet_5_0_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_1_0_clk_in_regs (.A(clknet_3_0_0_clk_in_regs),
    .X(clknet_5_1_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_2_0_clk_in_regs (.A(clknet_3_0_0_clk_in_regs),
    .X(clknet_5_2_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_3_0_clk_in_regs (.A(clknet_3_0_0_clk_in_regs),
    .X(clknet_5_3_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_4_0_clk_in_regs (.A(clknet_3_1_0_clk_in_regs),
    .X(clknet_5_4_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_5_0_clk_in_regs (.A(clknet_3_1_0_clk_in_regs),
    .X(clknet_5_5_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_6_0_clk_in_regs (.A(clknet_3_1_0_clk_in_regs),
    .X(clknet_5_6_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_7_0_clk_in_regs (.A(clknet_3_1_0_clk_in_regs),
    .X(clknet_5_7_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_8_0_clk_in_regs (.A(clknet_3_2_0_clk_in_regs),
    .X(clknet_5_8_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_9_0_clk_in_regs (.A(clknet_3_2_0_clk_in_regs),
    .X(clknet_5_9_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_10_0_clk_in_regs (.A(clknet_3_2_0_clk_in_regs),
    .X(clknet_5_10_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_11_0_clk_in_regs (.A(clknet_3_2_0_clk_in_regs),
    .X(clknet_5_11_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_12_0_clk_in_regs (.A(clknet_3_3_0_clk_in_regs),
    .X(clknet_5_12_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_13_0_clk_in_regs (.A(clknet_3_3_0_clk_in_regs),
    .X(clknet_5_13_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_14_0_clk_in_regs (.A(clknet_3_3_0_clk_in_regs),
    .X(clknet_5_14_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_15_0_clk_in_regs (.A(clknet_3_3_0_clk_in_regs),
    .X(clknet_5_15_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_16_0_clk_in_regs (.A(clknet_3_4_0_clk_in_regs),
    .X(clknet_5_16_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_17_0_clk_in_regs (.A(clknet_3_4_0_clk_in_regs),
    .X(clknet_5_17_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_18_0_clk_in_regs (.A(clknet_3_4_0_clk_in_regs),
    .X(clknet_5_18_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_19_0_clk_in_regs (.A(clknet_3_4_0_clk_in_regs),
    .X(clknet_5_19_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_20_0_clk_in_regs (.A(clknet_3_5_0_clk_in_regs),
    .X(clknet_5_20_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_21_0_clk_in_regs (.A(clknet_3_5_0_clk_in_regs),
    .X(clknet_5_21_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_22_0_clk_in_regs (.A(clknet_3_5_0_clk_in_regs),
    .X(clknet_5_22_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_23_0_clk_in_regs (.A(clknet_3_5_0_clk_in_regs),
    .X(clknet_5_23_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_24_0_clk_in_regs (.A(clknet_3_6_0_clk_in_regs),
    .X(clknet_5_24_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_25_0_clk_in_regs (.A(clknet_3_6_0_clk_in_regs),
    .X(clknet_5_25_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_26_0_clk_in_regs (.A(clknet_3_6_0_clk_in_regs),
    .X(clknet_5_26_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_27_0_clk_in_regs (.A(clknet_3_6_0_clk_in_regs),
    .X(clknet_5_27_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_28_0_clk_in_regs (.A(clknet_3_7_0_clk_in_regs),
    .X(clknet_5_28_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_29_0_clk_in_regs (.A(clknet_3_7_0_clk_in_regs),
    .X(clknet_5_29_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_30_0_clk_in_regs (.A(clknet_3_7_0_clk_in_regs),
    .X(clknet_5_30_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_31_0_clk_in_regs (.A(clknet_3_7_0_clk_in_regs),
    .X(clknet_5_31_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_0__f_clk_in_regs (.A(clknet_5_0_0_clk_in_regs),
    .X(clknet_6_0__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_1__f_clk_in_regs (.A(clknet_5_0_0_clk_in_regs),
    .X(clknet_6_1__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_2__f_clk_in_regs (.A(clknet_5_1_0_clk_in_regs),
    .X(clknet_6_2__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_3__f_clk_in_regs (.A(clknet_5_1_0_clk_in_regs),
    .X(clknet_6_3__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_4__f_clk_in_regs (.A(clknet_5_2_0_clk_in_regs),
    .X(clknet_6_4__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_5__f_clk_in_regs (.A(clknet_5_2_0_clk_in_regs),
    .X(clknet_6_5__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_6__f_clk_in_regs (.A(clknet_5_3_0_clk_in_regs),
    .X(clknet_6_6__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_7__f_clk_in_regs (.A(clknet_5_3_0_clk_in_regs),
    .X(clknet_6_7__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_8__f_clk_in_regs (.A(clknet_5_4_0_clk_in_regs),
    .X(clknet_6_8__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_9__f_clk_in_regs (.A(clknet_5_4_0_clk_in_regs),
    .X(clknet_6_9__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_10__f_clk_in_regs (.A(clknet_5_5_0_clk_in_regs),
    .X(clknet_6_10__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_11__f_clk_in_regs (.A(clknet_5_5_0_clk_in_regs),
    .X(clknet_6_11__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_12__f_clk_in_regs (.A(clknet_5_6_0_clk_in_regs),
    .X(clknet_6_12__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_13__f_clk_in_regs (.A(clknet_5_6_0_clk_in_regs),
    .X(clknet_6_13__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_14__f_clk_in_regs (.A(clknet_5_7_0_clk_in_regs),
    .X(clknet_6_14__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_15__f_clk_in_regs (.A(clknet_5_7_0_clk_in_regs),
    .X(clknet_6_15__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_16__f_clk_in_regs (.A(clknet_5_8_0_clk_in_regs),
    .X(clknet_6_16__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_17__f_clk_in_regs (.A(clknet_5_8_0_clk_in_regs),
    .X(clknet_6_17__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_18__f_clk_in_regs (.A(clknet_5_9_0_clk_in_regs),
    .X(clknet_6_18__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_19__f_clk_in_regs (.A(clknet_5_9_0_clk_in_regs),
    .X(clknet_6_19__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_20__f_clk_in_regs (.A(clknet_5_10_0_clk_in_regs),
    .X(clknet_6_20__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_21__f_clk_in_regs (.A(clknet_5_10_0_clk_in_regs),
    .X(clknet_6_21__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_22__f_clk_in_regs (.A(clknet_5_11_0_clk_in_regs),
    .X(clknet_6_22__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_23__f_clk_in_regs (.A(clknet_5_11_0_clk_in_regs),
    .X(clknet_6_23__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_24__f_clk_in_regs (.A(clknet_5_12_0_clk_in_regs),
    .X(clknet_6_24__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_25__f_clk_in_regs (.A(clknet_5_12_0_clk_in_regs),
    .X(clknet_6_25__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_26__f_clk_in_regs (.A(clknet_5_13_0_clk_in_regs),
    .X(clknet_6_26__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_27__f_clk_in_regs (.A(clknet_5_13_0_clk_in_regs),
    .X(clknet_6_27__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_28__f_clk_in_regs (.A(clknet_5_14_0_clk_in_regs),
    .X(clknet_6_28__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_29__f_clk_in_regs (.A(clknet_5_14_0_clk_in_regs),
    .X(clknet_6_29__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_30__f_clk_in_regs (.A(clknet_5_15_0_clk_in_regs),
    .X(clknet_6_30__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_31__f_clk_in_regs (.A(clknet_5_15_0_clk_in_regs),
    .X(clknet_6_31__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_32__f_clk_in_regs (.A(clknet_5_16_0_clk_in_regs),
    .X(clknet_6_32__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_33__f_clk_in_regs (.A(clknet_5_16_0_clk_in_regs),
    .X(clknet_6_33__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_34__f_clk_in_regs (.A(clknet_5_17_0_clk_in_regs),
    .X(clknet_6_34__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_35__f_clk_in_regs (.A(clknet_5_17_0_clk_in_regs),
    .X(clknet_6_35__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_36__f_clk_in_regs (.A(clknet_5_18_0_clk_in_regs),
    .X(clknet_6_36__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_37__f_clk_in_regs (.A(clknet_5_18_0_clk_in_regs),
    .X(clknet_6_37__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_38__f_clk_in_regs (.A(clknet_5_19_0_clk_in_regs),
    .X(clknet_6_38__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_39__f_clk_in_regs (.A(clknet_5_19_0_clk_in_regs),
    .X(clknet_6_39__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_40__f_clk_in_regs (.A(clknet_5_20_0_clk_in_regs),
    .X(clknet_6_40__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_41__f_clk_in_regs (.A(clknet_5_20_0_clk_in_regs),
    .X(clknet_6_41__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_42__f_clk_in_regs (.A(clknet_5_21_0_clk_in_regs),
    .X(clknet_6_42__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_43__f_clk_in_regs (.A(clknet_5_21_0_clk_in_regs),
    .X(clknet_6_43__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_44__f_clk_in_regs (.A(clknet_5_22_0_clk_in_regs),
    .X(clknet_6_44__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_45__f_clk_in_regs (.A(clknet_5_22_0_clk_in_regs),
    .X(clknet_6_45__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_46__f_clk_in_regs (.A(clknet_5_23_0_clk_in_regs),
    .X(clknet_6_46__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_47__f_clk_in_regs (.A(clknet_5_23_0_clk_in_regs),
    .X(clknet_6_47__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_48__f_clk_in_regs (.A(clknet_5_24_0_clk_in_regs),
    .X(clknet_6_48__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_49__f_clk_in_regs (.A(clknet_5_24_0_clk_in_regs),
    .X(clknet_6_49__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_50__f_clk_in_regs (.A(clknet_5_25_0_clk_in_regs),
    .X(clknet_6_50__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_51__f_clk_in_regs (.A(clknet_5_25_0_clk_in_regs),
    .X(clknet_6_51__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_52__f_clk_in_regs (.A(clknet_5_26_0_clk_in_regs),
    .X(clknet_6_52__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_53__f_clk_in_regs (.A(clknet_5_26_0_clk_in_regs),
    .X(clknet_6_53__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_54__f_clk_in_regs (.A(clknet_5_27_0_clk_in_regs),
    .X(clknet_6_54__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_55__f_clk_in_regs (.A(clknet_5_27_0_clk_in_regs),
    .X(clknet_6_55__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_56__f_clk_in_regs (.A(clknet_5_28_0_clk_in_regs),
    .X(clknet_6_56__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_57__f_clk_in_regs (.A(clknet_5_28_0_clk_in_regs),
    .X(clknet_6_57__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_58__f_clk_in_regs (.A(clknet_5_29_0_clk_in_regs),
    .X(clknet_6_58__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_59__f_clk_in_regs (.A(clknet_5_29_0_clk_in_regs),
    .X(clknet_6_59__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_60__f_clk_in_regs (.A(clknet_5_30_0_clk_in_regs),
    .X(clknet_6_60__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_61__f_clk_in_regs (.A(clknet_5_30_0_clk_in_regs),
    .X(clknet_6_61__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_62__f_clk_in_regs (.A(clknet_5_31_0_clk_in_regs),
    .X(clknet_6_62__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_6_63__f_clk_in_regs (.A(clknet_5_31_0_clk_in_regs),
    .X(clknet_6_63__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_6_0__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_6_3__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload2 (.A(clknet_6_5__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload3 (.A(clknet_6_9__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload4 (.A(clknet_6_11__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_16 clkload5 (.A(clknet_6_12__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload6 (.A(clknet_6_15__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_8 clkload7 (.A(clknet_6_17__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload8 (.A(clknet_6_18__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkload9 (.A(clknet_6_20__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkinv_8 clkload10 (.A(clknet_6_22__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_16 clkload11 (.A(clknet_6_25__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkinv_16 clkload12 (.A(clknet_6_27__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_12 clkload13 (.A(clknet_6_29__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_12 clkload14 (.A(clknet_6_31__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkinv_16 clkload15 (.A(clknet_6_32__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkinv_8 clkload16 (.A(clknet_6_35__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkinv_16 clkload17 (.A(clknet_6_36__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload18 (.A(clknet_6_39__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkinv_16 clkload19 (.A(clknet_6_41__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_12 clkload20 (.A(clknet_6_43__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkinv_8 clkload21 (.A(clknet_6_46__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload22 (.A(clknet_6_48__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_8 clkload23 (.A(clknet_6_51__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_16 clkload24 (.A(clknet_6_53__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_16 clkload25 (.A(clknet_6_54__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkinv_16 clkload26 (.A(clknet_6_56__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkload27 (.A(clknet_6_58__leaf_clk_in_regs));
 sky130_fd_sc_hd__clkinv_16 clkload28 (.A(clknet_6_61__leaf_clk_in_regs));
 sky130_fd_sc_hd__inv_16 clkload29 (.A(clknet_6_63__leaf_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload30 (.A(clknet_leaf_725_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload31 (.A(clknet_leaf_727_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload32 (.A(clknet_leaf_729_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload33 (.A(clknet_leaf_732_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload34 (.A(clknet_leaf_716_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload35 (.A(clknet_leaf_717_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload36 (.A(clknet_leaf_723_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload37 (.A(clknet_leaf_724_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload38 (.A(clknet_leaf_733_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload39 (.A(clknet_leaf_718_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload40 (.A(clknet_leaf_719_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload41 (.A(clknet_leaf_720_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload42 (.A(clknet_leaf_721_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload43 (.A(clknet_leaf_734_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload44 (.A(clknet_leaf_735_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload45 (.A(clknet_leaf_736_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload46 (.A(clknet_leaf_737_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload47 (.A(clknet_leaf_740_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload48 (.A(clknet_leaf_613_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload49 (.A(clknet_leaf_651_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload50 (.A(clknet_leaf_652_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload51 (.A(clknet_leaf_653_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload52 (.A(clknet_leaf_654_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload53 (.A(clknet_leaf_655_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload54 (.A(clknet_leaf_738_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload55 (.A(clknet_leaf_660_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload56 (.A(clknet_leaf_661_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload57 (.A(clknet_leaf_715_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload58 (.A(clknet_leaf_667_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload59 (.A(clknet_leaf_650_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload60 (.A(clknet_leaf_656_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload61 (.A(clknet_leaf_657_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload62 (.A(clknet_leaf_658_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload63 (.A(clknet_leaf_662_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload64 (.A(clknet_leaf_644_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload65 (.A(clknet_leaf_645_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload66 (.A(clknet_leaf_646_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload67 (.A(clknet_leaf_663_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload68 (.A(clknet_leaf_665_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload69 (.A(clknet_leaf_765_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload70 (.A(clknet_leaf_771_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload71 (.A(clknet_leaf_772_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload72 (.A(clknet_leaf_773_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload73 (.A(clknet_leaf_774_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload74 (.A(clknet_leaf_776_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload75 (.A(clknet_leaf_777_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload76 (.A(clknet_leaf_762_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload77 (.A(clknet_leaf_763_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload78 (.A(clknet_leaf_766_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload79 (.A(clknet_leaf_767_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload80 (.A(clknet_leaf_778_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload81 (.A(clknet_leaf_779_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload82 (.A(clknet_leaf_6_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload83 (.A(clknet_leaf_9_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload84 (.A(clknet_leaf_10_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload85 (.A(clknet_leaf_781_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload86 (.A(clknet_leaf_783_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload87 (.A(clknet_leaf_784_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload88 (.A(clknet_leaf_786_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload89 (.A(clknet_leaf_789_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload90 (.A(clknet_leaf_790_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload91 (.A(clknet_leaf_11_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload92 (.A(clknet_leaf_12_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload93 (.A(clknet_leaf_13_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload94 (.A(clknet_leaf_14_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload95 (.A(clknet_leaf_15_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload96 (.A(clknet_leaf_16_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload97 (.A(clknet_leaf_17_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload98 (.A(clknet_leaf_768_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload99 (.A(clknet_leaf_769_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload100 (.A(clknet_leaf_728_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload101 (.A(clknet_leaf_746_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload102 (.A(clknet_leaf_748_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload103 (.A(clknet_leaf_750_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload104 (.A(clknet_leaf_751_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload105 (.A(clknet_leaf_760_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload106 (.A(clknet_leaf_761_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload107 (.A(clknet_leaf_608_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload108 (.A(clknet_leaf_609_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload109 (.A(clknet_leaf_610_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload110 (.A(clknet_leaf_611_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload111 (.A(clknet_leaf_739_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload112 (.A(clknet_leaf_741_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload113 (.A(clknet_leaf_744_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload114 (.A(clknet_leaf_745_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload115 (.A(clknet_leaf_753_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload116 (.A(clknet_leaf_754_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload117 (.A(clknet_leaf_18_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload118 (.A(clknet_leaf_19_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload119 (.A(clknet_leaf_23_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload120 (.A(clknet_leaf_26_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload121 (.A(clknet_leaf_330_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload122 (.A(clknet_leaf_331_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload123 (.A(clknet_leaf_332_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload124 (.A(clknet_leaf_759_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload125 (.A(clknet_leaf_585_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload126 (.A(clknet_leaf_587_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload127 (.A(clknet_leaf_591_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload128 (.A(clknet_leaf_752_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload129 (.A(clknet_leaf_755_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload130 (.A(clknet_leaf_756_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload131 (.A(clknet_leaf_669_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload132 (.A(clknet_leaf_671_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload133 (.A(clknet_leaf_672_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload134 (.A(clknet_leaf_673_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload135 (.A(clknet_leaf_675_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload136 (.A(clknet_leaf_678_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload137 (.A(clknet_leaf_680_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload138 (.A(clknet_leaf_681_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload139 (.A(clknet_leaf_682_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload140 (.A(clknet_leaf_698_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload141 (.A(clknet_leaf_701_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload142 (.A(clknet_leaf_696_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload143 (.A(clknet_leaf_700_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload144 (.A(clknet_leaf_702_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload145 (.A(clknet_leaf_703_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload146 (.A(clknet_leaf_704_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload147 (.A(clknet_leaf_705_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload148 (.A(clknet_leaf_708_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload149 (.A(clknet_leaf_711_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload150 (.A(clknet_leaf_712_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload151 (.A(clknet_leaf_688_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload152 (.A(clknet_leaf_689_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload153 (.A(clknet_leaf_692_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload154 (.A(clknet_leaf_709_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload155 (.A(clknet_leaf_566_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload156 (.A(clknet_leaf_683_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload157 (.A(clknet_leaf_684_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload158 (.A(clknet_leaf_686_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload159 (.A(clknet_leaf_687_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload160 (.A(clknet_leaf_690_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload161 (.A(clknet_leaf_691_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload162 (.A(clknet_leaf_551_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload163 (.A(clknet_leaf_564_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload164 (.A(clknet_leaf_568_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload165 (.A(clknet_leaf_546_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload166 (.A(clknet_leaf_547_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload167 (.A(clknet_leaf_695_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload168 (.A(clknet_leaf_707_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload169 (.A(clknet_leaf_554_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload170 (.A(clknet_leaf_557_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload171 (.A(clknet_leaf_559_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload172 (.A(clknet_leaf_536_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload173 (.A(clknet_leaf_537_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload174 (.A(clknet_leaf_538_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload175 (.A(clknet_leaf_542_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload176 (.A(clknet_leaf_543_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload177 (.A(clknet_leaf_545_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload178 (.A(clknet_leaf_1_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload179 (.A(clknet_leaf_56_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload180 (.A(clknet_leaf_57_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload181 (.A(clknet_leaf_58_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload182 (.A(clknet_leaf_59_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload183 (.A(clknet_leaf_63_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload184 (.A(clknet_leaf_64_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload185 (.A(clknet_leaf_65_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload186 (.A(clknet_leaf_66_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload187 (.A(clknet_leaf_128_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload188 (.A(clknet_leaf_130_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload189 (.A(clknet_leaf_785_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload190 (.A(clknet_leaf_787_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload191 (.A(clknet_leaf_788_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload192 (.A(clknet_leaf_0_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload193 (.A(clknet_leaf_2_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload194 (.A(clknet_leaf_4_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload195 (.A(clknet_leaf_5_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload196 (.A(clknet_leaf_21_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload197 (.A(clknet_leaf_22_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload198 (.A(clknet_leaf_24_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload199 (.A(clknet_leaf_27_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload200 (.A(clknet_leaf_35_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload201 (.A(clknet_leaf_25_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload202 (.A(clknet_leaf_28_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload203 (.A(clknet_leaf_30_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload204 (.A(clknet_leaf_31_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload205 (.A(clknet_leaf_32_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload206 (.A(clknet_leaf_36_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload207 (.A(clknet_leaf_37_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload208 (.A(clknet_leaf_39_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload209 (.A(clknet_leaf_333_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload210 (.A(clknet_leaf_335_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload211 (.A(clknet_leaf_589_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload212 (.A(clknet_leaf_757_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload213 (.A(clknet_leaf_758_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload214 (.A(clknet_leaf_337_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload215 (.A(clknet_leaf_343_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload216 (.A(clknet_leaf_344_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload217 (.A(clknet_leaf_345_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload218 (.A(clknet_leaf_580_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload219 (.A(clknet_leaf_584_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload220 (.A(clknet_leaf_588_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload221 (.A(clknet_leaf_594_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload222 (.A(clknet_leaf_595_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload223 (.A(clknet_leaf_596_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload224 (.A(clknet_leaf_597_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload225 (.A(clknet_leaf_604_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload226 (.A(clknet_leaf_605_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload227 (.A(clknet_leaf_606_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload228 (.A(clknet_leaf_615_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload229 (.A(clknet_leaf_618_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload230 (.A(clknet_leaf_619_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload231 (.A(clknet_leaf_620_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload232 (.A(clknet_leaf_621_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload233 (.A(clknet_leaf_622_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload234 (.A(clknet_leaf_625_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload235 (.A(clknet_leaf_628_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload236 (.A(clknet_leaf_629_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload237 (.A(clknet_leaf_630_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload238 (.A(clknet_leaf_632_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload239 (.A(clknet_leaf_633_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload240 (.A(clknet_leaf_634_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload241 (.A(clknet_leaf_635_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload242 (.A(clknet_leaf_636_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload243 (.A(clknet_leaf_637_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload244 (.A(clknet_leaf_640_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload245 (.A(clknet_leaf_641_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload246 (.A(clknet_leaf_642_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload247 (.A(clknet_leaf_643_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload248 (.A(clknet_leaf_647_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload249 (.A(clknet_leaf_648_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload250 (.A(clknet_leaf_567_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload251 (.A(clknet_leaf_570_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload252 (.A(clknet_leaf_590_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload253 (.A(clknet_leaf_592_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload254 (.A(clknet_leaf_598_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload255 (.A(clknet_leaf_599_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload256 (.A(clknet_leaf_600_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload257 (.A(clknet_leaf_601_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload258 (.A(clknet_leaf_602_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload259 (.A(clknet_leaf_623_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload260 (.A(clknet_leaf_624_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload261 (.A(clknet_leaf_626_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload262 (.A(clknet_leaf_562_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload263 (.A(clknet_leaf_572_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload264 (.A(clknet_leaf_573_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload265 (.A(clknet_leaf_574_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload266 (.A(clknet_leaf_575_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload267 (.A(clknet_leaf_576_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload268 (.A(clknet_leaf_577_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload269 (.A(clknet_leaf_579_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload270 (.A(clknet_leaf_67_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload271 (.A(clknet_leaf_68_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload272 (.A(clknet_leaf_69_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload273 (.A(clknet_leaf_72_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload274 (.A(clknet_leaf_74_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload275 (.A(clknet_leaf_124_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload276 (.A(clknet_leaf_127_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload277 (.A(clknet_leaf_131_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload278 (.A(clknet_leaf_132_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload279 (.A(clknet_leaf_75_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload280 (.A(clknet_leaf_76_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload281 (.A(clknet_leaf_79_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload282 (.A(clknet_leaf_84_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload283 (.A(clknet_leaf_85_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload284 (.A(clknet_leaf_87_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload285 (.A(clknet_leaf_97_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload286 (.A(clknet_leaf_98_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload287 (.A(clknet_leaf_99_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload288 (.A(clknet_leaf_117_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload289 (.A(clknet_leaf_118_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload290 (.A(clknet_leaf_119_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload291 (.A(clknet_leaf_123_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload292 (.A(clknet_leaf_94_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload293 (.A(clknet_leaf_100_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload294 (.A(clknet_leaf_102_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload295 (.A(clknet_leaf_103_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload296 (.A(clknet_leaf_104_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload297 (.A(clknet_leaf_105_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload298 (.A(clknet_leaf_106_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload299 (.A(clknet_leaf_107_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload300 (.A(clknet_leaf_108_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload301 (.A(clknet_leaf_109_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload302 (.A(clknet_leaf_113_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload303 (.A(clknet_leaf_114_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload304 (.A(clknet_leaf_115_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload305 (.A(clknet_leaf_116_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload306 (.A(clknet_leaf_257_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload307 (.A(clknet_leaf_89_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload308 (.A(clknet_leaf_90_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload309 (.A(clknet_leaf_91_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload310 (.A(clknet_leaf_92_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload311 (.A(clknet_leaf_95_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload312 (.A(clknet_leaf_269_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload313 (.A(clknet_leaf_270_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload314 (.A(clknet_leaf_271_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload315 (.A(clknet_leaf_272_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload316 (.A(clknet_leaf_273_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload317 (.A(clknet_leaf_274_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload318 (.A(clknet_leaf_276_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload319 (.A(clknet_leaf_308_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload320 (.A(clknet_leaf_310_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload321 (.A(clknet_leaf_53_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload322 (.A(clknet_leaf_54_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload323 (.A(clknet_leaf_55_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload324 (.A(clknet_leaf_60_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload325 (.A(clknet_leaf_61_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload326 (.A(clknet_leaf_62_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload327 (.A(clknet_leaf_70_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload328 (.A(clknet_leaf_80_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload329 (.A(clknet_leaf_81_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload330 (.A(clknet_leaf_82_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload331 (.A(clknet_leaf_40_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload332 (.A(clknet_leaf_41_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload333 (.A(clknet_leaf_42_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload334 (.A(clknet_leaf_43_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload335 (.A(clknet_leaf_44_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload336 (.A(clknet_leaf_45_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload337 (.A(clknet_leaf_46_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload338 (.A(clknet_leaf_48_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload339 (.A(clknet_leaf_49_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload340 (.A(clknet_leaf_50_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload341 (.A(clknet_leaf_51_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload342 (.A(clknet_leaf_83_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload343 (.A(clknet_leaf_86_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload344 (.A(clknet_leaf_317_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload345 (.A(clknet_leaf_318_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload346 (.A(clknet_leaf_329_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload347 (.A(clknet_leaf_304_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload348 (.A(clknet_leaf_305_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload349 (.A(clknet_leaf_311_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload350 (.A(clknet_leaf_312_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload351 (.A(clknet_leaf_313_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload352 (.A(clknet_leaf_314_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload353 (.A(clknet_leaf_315_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload354 (.A(clknet_leaf_316_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload355 (.A(clknet_leaf_320_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload356 (.A(clknet_leaf_321_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload357 (.A(clknet_leaf_323_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload358 (.A(clknet_leaf_322_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload359 (.A(clknet_leaf_324_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload360 (.A(clknet_leaf_325_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload361 (.A(clknet_leaf_327_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload362 (.A(clknet_leaf_328_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload363 (.A(clknet_leaf_338_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload364 (.A(clknet_leaf_339_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload365 (.A(clknet_leaf_342_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload366 (.A(clknet_leaf_275_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload367 (.A(clknet_leaf_277_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload368 (.A(clknet_leaf_278_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload369 (.A(clknet_leaf_279_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload370 (.A(clknet_leaf_288_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload371 (.A(clknet_leaf_289_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload372 (.A(clknet_leaf_290_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload373 (.A(clknet_leaf_295_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload374 (.A(clknet_leaf_296_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload375 (.A(clknet_leaf_297_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload376 (.A(clknet_leaf_298_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload377 (.A(clknet_leaf_299_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload378 (.A(clknet_leaf_300_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload379 (.A(clknet_leaf_302_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload380 (.A(clknet_leaf_356_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload381 (.A(clknet_leaf_357_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload382 (.A(clknet_leaf_358_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload383 (.A(clknet_leaf_361_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload384 (.A(clknet_leaf_362_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload385 (.A(clknet_leaf_368_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload386 (.A(clknet_leaf_111_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload387 (.A(clknet_leaf_134_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload388 (.A(clknet_leaf_138_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload389 (.A(clknet_leaf_242_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload390 (.A(clknet_leaf_248_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload391 (.A(clknet_leaf_250_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload392 (.A(clknet_leaf_251_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload393 (.A(clknet_leaf_252_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload394 (.A(clknet_leaf_253_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload395 (.A(clknet_leaf_254_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload396 (.A(clknet_leaf_258_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload397 (.A(clknet_leaf_259_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload398 (.A(clknet_leaf_260_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload399 (.A(clknet_leaf_261_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload400 (.A(clknet_leaf_262_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload401 (.A(clknet_leaf_263_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload402 (.A(clknet_leaf_218_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload403 (.A(clknet_leaf_221_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload404 (.A(clknet_leaf_264_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload405 (.A(clknet_leaf_265_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload406 (.A(clknet_leaf_266_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload407 (.A(clknet_leaf_281_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload408 (.A(clknet_leaf_283_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload409 (.A(clknet_leaf_284_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload410 (.A(clknet_leaf_285_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload411 (.A(clknet_leaf_286_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload412 (.A(clknet_leaf_287_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload413 (.A(clknet_leaf_291_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload414 (.A(clknet_leaf_292_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload415 (.A(clknet_leaf_293_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload416 (.A(clknet_leaf_367_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload417 (.A(clknet_leaf_352_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload418 (.A(clknet_leaf_359_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload419 (.A(clknet_leaf_360_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload420 (.A(clknet_leaf_369_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload421 (.A(clknet_leaf_370_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload422 (.A(clknet_leaf_376_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload423 (.A(clknet_leaf_377_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload424 (.A(clknet_leaf_378_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload425 (.A(clknet_leaf_384_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload426 (.A(clknet_leaf_385_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload427 (.A(clknet_leaf_341_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload428 (.A(clknet_leaf_346_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload429 (.A(clknet_leaf_347_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload430 (.A(clknet_leaf_348_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload431 (.A(clknet_leaf_349_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload432 (.A(clknet_leaf_350_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload433 (.A(clknet_leaf_353_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload434 (.A(clknet_leaf_354_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload435 (.A(clknet_leaf_355_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload436 (.A(clknet_leaf_381_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload437 (.A(clknet_leaf_383_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload438 (.A(clknet_leaf_375_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload439 (.A(clknet_leaf_387_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload440 (.A(clknet_leaf_389_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload441 (.A(clknet_leaf_560_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload442 (.A(clknet_leaf_519_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload443 (.A(clknet_leaf_527_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload444 (.A(clknet_leaf_528_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload445 (.A(clknet_leaf_530_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload446 (.A(clknet_leaf_531_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload447 (.A(clknet_leaf_532_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload448 (.A(clknet_leaf_533_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload449 (.A(clknet_leaf_534_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload450 (.A(clknet_leaf_202_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload451 (.A(clknet_leaf_204_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload452 (.A(clknet_leaf_216_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload453 (.A(clknet_leaf_224_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload454 (.A(clknet_leaf_226_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload455 (.A(clknet_leaf_227_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload456 (.A(clknet_leaf_228_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload457 (.A(clknet_leaf_236_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload458 (.A(clknet_leaf_237_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload459 (.A(clknet_leaf_205_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload460 (.A(clknet_leaf_206_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload461 (.A(clknet_leaf_207_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload462 (.A(clknet_leaf_208_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload463 (.A(clknet_leaf_214_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload464 (.A(clknet_leaf_215_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload465 (.A(clknet_leaf_363_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload466 (.A(clknet_leaf_425_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload467 (.A(clknet_leaf_427_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload468 (.A(clknet_leaf_428_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload469 (.A(clknet_leaf_433_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload470 (.A(clknet_leaf_135_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload471 (.A(clknet_leaf_140_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload472 (.A(clknet_leaf_223_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload473 (.A(clknet_leaf_225_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload474 (.A(clknet_leaf_238_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload475 (.A(clknet_leaf_240_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload476 (.A(clknet_leaf_241_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload477 (.A(clknet_leaf_243_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload478 (.A(clknet_leaf_244_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload479 (.A(clknet_leaf_245_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload480 (.A(clknet_leaf_246_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload481 (.A(clknet_leaf_247_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload482 (.A(clknet_leaf_249_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload483 (.A(clknet_leaf_209_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload484 (.A(clknet_leaf_210_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload485 (.A(clknet_leaf_211_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload486 (.A(clknet_leaf_212_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload487 (.A(clknet_leaf_217_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload488 (.A(clknet_leaf_219_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload489 (.A(clknet_leaf_220_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload490 (.A(clknet_leaf_222_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload491 (.A(clknet_leaf_239_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload492 (.A(clknet_leaf_294_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload493 (.A(clknet_leaf_364_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload494 (.A(clknet_leaf_424_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload495 (.A(clknet_leaf_365_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload496 (.A(clknet_leaf_366_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload497 (.A(clknet_leaf_371_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 clkload498 (.A(clknet_leaf_372_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload499 (.A(clknet_leaf_373_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload500 (.A(clknet_leaf_374_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload501 (.A(clknet_leaf_393_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload502 (.A(clknet_leaf_414_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload503 (.A(clknet_leaf_525_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload504 (.A(clknet_leaf_416_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload505 (.A(clknet_leaf_417_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload506 (.A(clknet_leaf_418_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload507 (.A(clknet_leaf_419_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload508 (.A(clknet_leaf_423_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload509 (.A(clknet_leaf_429_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload510 (.A(clknet_leaf_430_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload511 (.A(clknet_leaf_431_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload512 (.A(clknet_leaf_432_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload513 (.A(clknet_leaf_394_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload514 (.A(clknet_leaf_395_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload515 (.A(clknet_leaf_396_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload516 (.A(clknet_leaf_397_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload517 (.A(clknet_leaf_399_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload518 (.A(clknet_leaf_406_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload519 (.A(clknet_leaf_408_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload520 (.A(clknet_leaf_409_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload521 (.A(clknet_leaf_410_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload522 (.A(clknet_leaf_411_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload523 (.A(clknet_leaf_412_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload524 (.A(clknet_leaf_413_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload525 (.A(clknet_leaf_415_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload526 (.A(clknet_leaf_143_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload527 (.A(clknet_leaf_145_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload528 (.A(clknet_leaf_146_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload529 (.A(clknet_leaf_147_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload530 (.A(clknet_leaf_149_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload531 (.A(clknet_leaf_188_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload532 (.A(clknet_leaf_189_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload533 (.A(clknet_leaf_190_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload534 (.A(clknet_leaf_191_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload535 (.A(clknet_leaf_193_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload536 (.A(clknet_leaf_229_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload537 (.A(clknet_leaf_232_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload538 (.A(clknet_leaf_233_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload539 (.A(clknet_leaf_174_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload540 (.A(clknet_leaf_177_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload541 (.A(clknet_leaf_178_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload542 (.A(clknet_leaf_179_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload543 (.A(clknet_leaf_180_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload544 (.A(clknet_leaf_181_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload545 (.A(clknet_leaf_182_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload546 (.A(clknet_leaf_183_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload547 (.A(clknet_leaf_184_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload548 (.A(clknet_leaf_185_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload549 (.A(clknet_leaf_186_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload550 (.A(clknet_leaf_187_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload551 (.A(clknet_leaf_192_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload552 (.A(clknet_leaf_196_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload553 (.A(clknet_leaf_197_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload554 (.A(clknet_leaf_198_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload555 (.A(clknet_leaf_199_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload556 (.A(clknet_leaf_200_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload557 (.A(clknet_leaf_434_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload558 (.A(clknet_leaf_435_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload559 (.A(clknet_leaf_436_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload560 (.A(clknet_leaf_458_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload561 (.A(clknet_leaf_148_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload562 (.A(clknet_leaf_150_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload563 (.A(clknet_leaf_151_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload564 (.A(clknet_leaf_152_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload565 (.A(clknet_leaf_153_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload566 (.A(clknet_leaf_154_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload567 (.A(clknet_leaf_155_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload568 (.A(clknet_leaf_156_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload569 (.A(clknet_leaf_158_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload570 (.A(clknet_leaf_159_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload571 (.A(clknet_leaf_160_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload572 (.A(clknet_leaf_161_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload573 (.A(clknet_leaf_162_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload574 (.A(clknet_leaf_163_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload575 (.A(clknet_leaf_164_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload576 (.A(clknet_leaf_165_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload577 (.A(clknet_leaf_166_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload578 (.A(clknet_leaf_167_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload579 (.A(clknet_leaf_168_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload580 (.A(clknet_leaf_169_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload581 (.A(clknet_leaf_170_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload582 (.A(clknet_leaf_171_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload583 (.A(clknet_leaf_173_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload584 (.A(clknet_leaf_175_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload585 (.A(clknet_leaf_176_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload586 (.A(clknet_leaf_460_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload587 (.A(clknet_leaf_466_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload588 (.A(clknet_leaf_467_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload589 (.A(clknet_leaf_468_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload590 (.A(clknet_leaf_469_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload591 (.A(clknet_leaf_470_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload592 (.A(clknet_leaf_437_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload593 (.A(clknet_leaf_438_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload594 (.A(clknet_leaf_439_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload595 (.A(clknet_leaf_440_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload596 (.A(clknet_leaf_441_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload597 (.A(clknet_leaf_442_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload598 (.A(clknet_leaf_443_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload599 (.A(clknet_leaf_444_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload600 (.A(clknet_leaf_445_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload601 (.A(clknet_leaf_447_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload602 (.A(clknet_leaf_448_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload603 (.A(clknet_leaf_449_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload604 (.A(clknet_leaf_450_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload605 (.A(clknet_leaf_453_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload606 (.A(clknet_leaf_454_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload607 (.A(clknet_leaf_455_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload608 (.A(clknet_leaf_456_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload609 (.A(clknet_leaf_457_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload610 (.A(clknet_leaf_459_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload611 (.A(clknet_leaf_491_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload612 (.A(clknet_leaf_492_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload613 (.A(clknet_leaf_493_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload614 (.A(clknet_leaf_398_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload615 (.A(clknet_leaf_400_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload616 (.A(clknet_leaf_401_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload617 (.A(clknet_leaf_402_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload618 (.A(clknet_leaf_403_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload619 (.A(clknet_leaf_404_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload620 (.A(clknet_leaf_405_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload621 (.A(clknet_leaf_494_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload622 (.A(clknet_leaf_506_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload623 (.A(clknet_leaf_507_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload624 (.A(clknet_leaf_508_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload625 (.A(clknet_leaf_509_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload626 (.A(clknet_leaf_511_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload627 (.A(clknet_leaf_512_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload628 (.A(clknet_leaf_513_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload629 (.A(clknet_leaf_451_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload630 (.A(clknet_leaf_452_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload631 (.A(clknet_leaf_461_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload632 (.A(clknet_leaf_462_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload633 (.A(clknet_leaf_463_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload634 (.A(clknet_leaf_464_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload635 (.A(clknet_leaf_465_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload636 (.A(clknet_leaf_471_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload637 (.A(clknet_leaf_472_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload638 (.A(clknet_leaf_473_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload639 (.A(clknet_leaf_474_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload640 (.A(clknet_leaf_475_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload641 (.A(clknet_leaf_476_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload642 (.A(clknet_leaf_477_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload643 (.A(clknet_leaf_479_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload644 (.A(clknet_leaf_480_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload645 (.A(clknet_leaf_486_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload646 (.A(clknet_leaf_487_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload647 (.A(clknet_leaf_488_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload648 (.A(clknet_leaf_489_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload649 (.A(clknet_leaf_481_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload650 (.A(clknet_leaf_482_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload651 (.A(clknet_leaf_483_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload652 (.A(clknet_leaf_484_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload653 (.A(clknet_leaf_485_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload654 (.A(clknet_leaf_490_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload655 (.A(clknet_leaf_495_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload656 (.A(clknet_leaf_496_clk_in_regs));
 sky130_fd_sc_hd__clkinv_2 clkload657 (.A(clknet_leaf_498_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload658 (.A(clknet_leaf_499_clk_in_regs));
 sky130_fd_sc_hd__bufinv_16 clkload659 (.A(clknet_leaf_500_clk_in_regs));
 sky130_fd_sc_hd__inv_6 clkload660 (.A(clknet_leaf_501_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload661 (.A(clknet_leaf_502_clk_in_regs));
 sky130_fd_sc_hd__clkinv_1 clkload662 (.A(clknet_leaf_503_clk_in_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload663 (.A(clknet_leaf_504_clk_in_regs));
 sky130_fd_sc_hd__clkinv_4 clkload664 (.A(clknet_leaf_505_clk_in_regs));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_0_sys_clk_in (.A(clk_in),
    .X(delaynet_0_sys_clk_in));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_1_sys_clk_in (.A(delaynet_0_sys_clk_in),
    .X(delaynet_1_sys_clk_in));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_2_sys_clk_in (.A(delaynet_1_sys_clk_in),
    .X(delaynet_2_sys_clk_in));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_3_sys_clk_in (.A(delaynet_2_sys_clk_in),
    .X(delaynet_3_sys_clk_in));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_4_sys_clk_in (.A(delaynet_3_sys_clk_in),
    .X(delaynet_4_sys_clk_in));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_5_sys_clk_in (.A(delaynet_4_sys_clk_in),
    .X(delaynet_5_sys_clk_in));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_6_sys_clk_in (.A(delaynet_5_sys_clk_in),
    .X(delaynet_6_sys_clk_in));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_7_sys_clk_in (.A(delaynet_6_sys_clk_in),
    .X(delaynet_7_sys_clk_in));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3036 (.A(\inst$top.soc.cpu.loadstore.dbus__dat_w[9] ),
    .X(net3035));
 sky130_fd_sc_hd__buf_6 wire3037 (.A(_17158_),
    .X(net3036));
 sky130_fd_sc_hd__buf_4 wire3038 (.A(_12850_),
    .X(net3037));
 sky130_fd_sc_hd__buf_4 wire3039 (.A(_12836_),
    .X(net3038));
 sky130_fd_sc_hd__buf_4 wire3040 (.A(_12930_),
    .X(net3039));
 sky130_fd_sc_hd__clkbuf_8 wire3041 (.A(_12887_),
    .X(net3040));
 sky130_fd_sc_hd__buf_4 wire3042 (.A(_12873_),
    .X(net3041));
 sky130_fd_sc_hd__buf_16 load_slew3043 (.A(net1136),
    .X(net3042));
 sky130_fd_sc_hd__buf_8 load_slew3044 (.A(net1163),
    .X(net3043));
 sky130_fd_sc_hd__buf_16 wire3045 (.A(net1678),
    .X(net3044));
 sky130_fd_sc_hd__clkbuf_4 wire3046 (.A(_05616_),
    .X(net3045));
endmodule
